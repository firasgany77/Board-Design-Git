-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 5 2021 16:19:01

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "counter" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of counter
entity counter is
port (
    clk_2Hz : out std_logic;
    CLK_27mhz : in std_logic);
end counter;

-- Architecture of counter
-- View name is \INTERFACE\
architecture \INTERFACE\ of counter is

signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_1_0_\ : std_logic;
signal counter_1_1_cry_1 : std_logic;
signal counter_1_1_cry_2 : std_logic;
signal counter_1_1_cry_3 : std_logic;
signal counter_1_1_cry_4 : std_logic;
signal counter_1_1_cry_5 : std_logic;
signal counter_1_1_cry_6 : std_logic;
signal counter_1_1_cry_7 : std_logic;
signal counter_1_1_cry_8 : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal counter_1_1_cry_9 : std_logic;
signal counter_1_1_cry_10 : std_logic;
signal counter_1_1_cry_11 : std_logic;
signal counter_1_1_cry_12 : std_logic;
signal counter_1_1_cry_13 : std_logic;
signal counter_1_1_cry_14 : std_logic;
signal counter_1_1_cry_15 : std_logic;
signal counter_1_1_cry_16 : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal counter_1_1_cry_17 : std_logic;
signal counter_1_1_cry_18 : std_logic;
signal counter_1_1_cry_19 : std_logic;
signal counter_1_1_cry_20 : std_logic;
signal counter_1_1_cry_21 : std_logic;
signal counter_1_1_cry_22 : std_logic;
signal counter_1_1_cry_23 : std_logic;
signal counter_1_1_cry_24 : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal counter_1_1_cry_25 : std_logic;
signal counter_1_1_cry_26 : std_logic;
signal counter_1_1_cry_27 : std_logic;
signal counter_1_1_cry_28 : std_logic;
signal counter_1_1_cry_29 : std_logic;
signal counter_1_1_cry_30 : std_logic;
signal \counter_1Z0Z_29\ : std_logic;
signal \counter_1Z0Z_28\ : std_logic;
signal \counter_1Z0Z_30\ : std_logic;
signal \counter_1Z0Z_31\ : std_logic;
signal un4_counter_2_0_and : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal un4_counter_2_1_and : std_logic;
signal un4_counter_2_0 : std_logic;
signal un4_counter_2_1 : std_logic;
signal un4_counter_2_2 : std_logic;
signal un4_counter_2_3 : std_logic;
signal un4_counter_2_4 : std_logic;
signal un4_counter_2_5 : std_logic;
signal un4_counter_2_6 : std_logic;
signal un4_counter_2_7 : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal un4_counter_2_5_and : std_logic;
signal un4_counter_2_4_and : std_logic;
signal un4_counter_2_2_and : std_logic;
signal un4_counter_2_3_and : std_logic;
signal un4_counter_2_7_and : std_logic;
signal un4_counter_2_6_and : std_logic;
signal \counter_1Z0Z_5\ : std_logic;
signal \counter_1Z0Z_7\ : std_logic;
signal \counter_1Z0Z_6\ : std_logic;
signal \counter_1Z0Z_4\ : std_logic;
signal \counter_1Z0Z_8\ : std_logic;
signal \counter_1Z0Z_10\ : std_logic;
signal \counter_1Z0Z_9\ : std_logic;
signal \counter_1Z0Z_11\ : std_logic;
signal \counter_1Z0Z_13\ : std_logic;
signal \counter_1Z0Z_12\ : std_logic;
signal \counter_1Z0Z_15\ : std_logic;
signal \counter_1Z0Z_14\ : std_logic;
signal \counter_1Z0Z_18\ : std_logic;
signal \counter_1Z0Z_19\ : std_logic;
signal \counter_1Z0Z_17\ : std_logic;
signal \counter_1Z0Z_16\ : std_logic;
signal \counter_1Z0Z_20\ : std_logic;
signal \counter_1Z0Z_21\ : std_logic;
signal \counter_1Z0Z_23\ : std_logic;
signal \counter_1Z0Z_22\ : std_logic;
signal \counter_1Z0Z_27\ : std_logic;
signal \counter_1Z0Z_24\ : std_logic;
signal \counter_1Z0Z_25\ : std_logic;
signal \counter_1Z0Z_26\ : std_logic;
signal \counter_2Z0Z_0\ : std_logic;
signal \counter_2Z0Z_1\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \counter_2Z0Z_2\ : std_logic;
signal \counter_2_1_cry_1_THRU_CO\ : std_logic;
signal counter_2_1_cry_1 : std_logic;
signal \counter_2Z0Z_3\ : std_logic;
signal counter_2_1_cry_2 : std_logic;
signal \counter_2Z0Z_4\ : std_logic;
signal \counter_2_1_cry_3_THRU_CO\ : std_logic;
signal counter_2_1_cry_3 : std_logic;
signal \counter_2Z0Z_5\ : std_logic;
signal \counter_2_1_cry_4_THRU_CO\ : std_logic;
signal counter_2_1_cry_4 : std_logic;
signal \counter_2Z0Z_6\ : std_logic;
signal \counter_2_1_cry_5_THRU_CO\ : std_logic;
signal counter_2_1_cry_5 : std_logic;
signal \counter_2Z0Z_7\ : std_logic;
signal \counter_2_1_cry_6_THRU_CO\ : std_logic;
signal counter_2_1_cry_6 : std_logic;
signal \counter_2Z0Z_8\ : std_logic;
signal \counter_2_1_cry_7_THRU_CO\ : std_logic;
signal counter_2_1_cry_7 : std_logic;
signal counter_2_1_cry_8 : std_logic;
signal \counter_2Z0Z_9\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \counter_2Z0Z_10\ : std_logic;
signal counter_2_1_cry_9 : std_logic;
signal \counter_2Z0Z_11\ : std_logic;
signal counter_2_1_cry_10 : std_logic;
signal \counter_2Z0Z_12\ : std_logic;
signal counter_2_1_cry_11 : std_logic;
signal \counter_2Z0Z_13\ : std_logic;
signal counter_2_1_cry_12 : std_logic;
signal \counter_2Z0Z_14\ : std_logic;
signal counter_2_1_cry_13 : std_logic;
signal \counter_2Z0Z_15\ : std_logic;
signal counter_2_1_cry_14 : std_logic;
signal \counter_2Z0Z_16\ : std_logic;
signal counter_2_1_cry_15 : std_logic;
signal counter_2_1_cry_16 : std_logic;
signal \counter_2Z0Z_17\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \counter_2Z0Z_18\ : std_logic;
signal counter_2_1_cry_17 : std_logic;
signal \counter_2Z0Z_19\ : std_logic;
signal counter_2_1_cry_18 : std_logic;
signal \counter_2Z0Z_20\ : std_logic;
signal counter_2_1_cry_19 : std_logic;
signal \counter_2Z0Z_21\ : std_logic;
signal counter_2_1_cry_20 : std_logic;
signal \counter_2Z0Z_22\ : std_logic;
signal counter_2_1_cry_21 : std_logic;
signal \counter_2Z0Z_23\ : std_logic;
signal counter_2_1_cry_22 : std_logic;
signal \counter_2Z0Z_24\ : std_logic;
signal counter_2_1_cry_23 : std_logic;
signal counter_2_1_cry_24 : std_logic;
signal \counter_2Z0Z_25\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \counter_2Z0Z_26\ : std_logic;
signal counter_2_1_cry_25 : std_logic;
signal \counter_2Z0Z_27\ : std_logic;
signal counter_2_1_cry_26 : std_logic;
signal \counter_2Z0Z_28\ : std_logic;
signal counter_2_1_cry_27 : std_logic;
signal \counter_2Z0Z_29\ : std_logic;
signal counter_2_1_cry_28 : std_logic;
signal \counter_2Z0Z_30\ : std_logic;
signal counter_2_1_cry_29 : std_logic;
signal counter_2_1_cry_30 : std_logic;
signal \counter_2Z0Z_31\ : std_logic;
signal \clk_1Khz_cnv_0_g\ : std_logic;
signal \counter_1_1_cry_2_THRU_CO\ : std_logic;
signal \counter_1_1_cry_1_THRU_CO\ : std_logic;
signal \counter_1Z0Z_2\ : std_logic;
signal \counter_1Z0Z_3\ : std_logic;
signal \counter_1Z0Z_0\ : std_logic;
signal \counter_1Z0Z_1\ : std_logic;
signal un4_counter_1_0_and : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal un4_counter_1_1_and : std_logic;
signal un4_counter_1_0 : std_logic;
signal un4_counter_1_2_and : std_logic;
signal un4_counter_1_1 : std_logic;
signal un4_counter_1_3_and : std_logic;
signal un4_counter_1_2 : std_logic;
signal un4_counter_1_4_and : std_logic;
signal un4_counter_1_3 : std_logic;
signal un4_counter_1_5_and : std_logic;
signal un4_counter_1_4 : std_logic;
signal un4_counter_1_6_and : std_logic;
signal un4_counter_1_5 : std_logic;
signal un4_counter_1_7_and : std_logic;
signal un4_counter_1_6 : std_logic;
signal un4_counter_1_7 : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \un4_counter_1_7_THRU_CO_cascade_\ : std_logic;
signal \clk_1Khz_cnv_0\ : std_logic;
signal \clk_2Hz_cnv_m3_e_1\ : std_logic;
signal \clk_2Hz_c\ : std_logic;
signal \clk_1Khz_i\ : std_logic;
signal \clk_1MHz_i\ : std_logic;
signal \un4_counter_2_7_THRU_CO\ : std_logic;
signal \un4_counter_1_7_THRU_CO\ : std_logic;
signal \clk_1Khz_RNIDQNNZ0\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal un4_counter_3_1_and : std_logic;
signal un4_counter_3_0 : std_logic;
signal un4_counter_3_2_and : std_logic;
signal un4_counter_3_1 : std_logic;
signal un4_counter_3_3_and : std_logic;
signal un4_counter_3_2 : std_logic;
signal un4_counter_3_3 : std_logic;
signal un4_counter_3_4 : std_logic;
signal un4_counter_3_5 : std_logic;
signal un4_counter_3_6 : std_logic;
signal un4_counter_3_7 : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal un4_counter_3_7_and : std_logic;
signal un4_counter_3_5_and : std_logic;
signal un4_counter_3_4_and : std_logic;
signal un4_counter_3_0_and : std_logic;
signal un4_counter_3_6_and : std_logic;
signal \counter_3Z0Z_1\ : std_logic;
signal \counter_3Z0Z_0\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \counter_3Z0Z_2\ : std_logic;
signal counter_3_1_cry_1 : std_logic;
signal counter_3_1_cry_2 : std_logic;
signal \counter_3Z0Z_4\ : std_logic;
signal \counter_3_1_cry_3_THRU_CO\ : std_logic;
signal counter_3_1_cry_3 : std_logic;
signal \counter_3Z0Z_5\ : std_logic;
signal \counter_3_1_cry_4_THRU_CO\ : std_logic;
signal counter_3_1_cry_4 : std_logic;
signal \counter_3Z0Z_6\ : std_logic;
signal \counter_3_1_cry_5_THRU_CO\ : std_logic;
signal counter_3_1_cry_5 : std_logic;
signal \counter_3Z0Z_7\ : std_logic;
signal \counter_3_1_cry_6_THRU_CO\ : std_logic;
signal counter_3_1_cry_6 : std_logic;
signal \counter_3Z0Z_8\ : std_logic;
signal counter_3_1_cry_7 : std_logic;
signal counter_3_1_cry_8 : std_logic;
signal \counter_3Z0Z_9\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \counter_3Z0Z_10\ : std_logic;
signal counter_3_1_cry_9 : std_logic;
signal \counter_3Z0Z_11\ : std_logic;
signal counter_3_1_cry_10 : std_logic;
signal \counter_3Z0Z_12\ : std_logic;
signal counter_3_1_cry_11 : std_logic;
signal \counter_3Z0Z_13\ : std_logic;
signal counter_3_1_cry_12 : std_logic;
signal \counter_3Z0Z_14\ : std_logic;
signal counter_3_1_cry_13 : std_logic;
signal \counter_3Z0Z_15\ : std_logic;
signal counter_3_1_cry_14 : std_logic;
signal \counter_3Z0Z_16\ : std_logic;
signal counter_3_1_cry_15 : std_logic;
signal counter_3_1_cry_16 : std_logic;
signal \counter_3Z0Z_17\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \counter_3Z0Z_18\ : std_logic;
signal counter_3_1_cry_17 : std_logic;
signal \counter_3Z0Z_19\ : std_logic;
signal counter_3_1_cry_18 : std_logic;
signal \counter_3Z0Z_20\ : std_logic;
signal counter_3_1_cry_19 : std_logic;
signal \counter_3Z0Z_21\ : std_logic;
signal counter_3_1_cry_20 : std_logic;
signal \counter_3Z0Z_22\ : std_logic;
signal counter_3_1_cry_21 : std_logic;
signal \counter_3Z0Z_23\ : std_logic;
signal counter_3_1_cry_22 : std_logic;
signal \counter_3Z0Z_24\ : std_logic;
signal counter_3_1_cry_23 : std_logic;
signal counter_3_1_cry_24 : std_logic;
signal \counter_3Z0Z_25\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \counter_3Z0Z_26\ : std_logic;
signal counter_3_1_cry_25 : std_logic;
signal \counter_3Z0Z_27\ : std_logic;
signal counter_3_1_cry_26 : std_logic;
signal \counter_3Z0Z_28\ : std_logic;
signal counter_3_1_cry_27 : std_logic;
signal \counter_3Z0Z_29\ : std_logic;
signal counter_3_1_cry_28 : std_logic;
signal \counter_3Z0Z_30\ : std_logic;
signal counter_3_1_cry_29 : std_logic;
signal counter_3_1_cry_30 : std_logic;
signal \counter_3Z0Z_31\ : std_logic;
signal \counter_3_1_cry_2_THRU_CO\ : std_logic;
signal \un4_counter_3_7_THRU_CO\ : std_logic;
signal \counter_3Z0Z_3\ : std_logic;
signal \CLK_27mhz_0_0_c_g\ : std_logic;
signal \N_67_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_27mhz_wire\ : std_logic;
signal \clk_2Hz_wire\ : std_logic;

begin
    \CLK_27mhz_wire\ <= CLK_27mhz;
    clk_2Hz <= \clk_2Hz_wire\;

    \CLK_27mhz_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__4639\,
            GLOBALBUFFEROUTPUT => \CLK_27mhz_0_0_c_g\
        );

    \CLK_27mhz_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__4641\,
            DIN => \N__4640\,
            DOUT => \N__4639\,
            PACKAGEPIN => \CLK_27mhz_wire\
        );

    \CLK_27mhz_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4641\,
            PADOUT => \N__4640\,
            PADIN => \N__4639\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_2Hz_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__4630\,
            DIN => \N__4629\,
            DOUT => \N__4628\,
            PACKAGEPIN => \clk_2Hz_wire\
        );

    \clk_2Hz_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4630\,
            PADOUT => \N__4629\,
            PADIN => \N__4628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3774\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__995\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4607\
        );

    \I__994\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4604\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4607\,
            I => \counter_3Z0Z_25\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__4604\,
            I => \counter_3Z0Z_25\
        );

    \I__991\ : InMux
    port map (
            O => \N__4599\,
            I => \bfn_12_10_0_\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4596\,
            I => \N__4592\
        );

    \I__989\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4589\
        );

    \I__988\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4586\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4589\,
            I => \counter_3Z0Z_26\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4586\,
            I => \counter_3Z0Z_26\
        );

    \I__985\ : InMux
    port map (
            O => \N__4581\,
            I => counter_3_1_cry_25
        );

    \I__984\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4574\
        );

    \I__983\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4571\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4574\,
            I => \counter_3Z0Z_27\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4571\,
            I => \counter_3Z0Z_27\
        );

    \I__980\ : InMux
    port map (
            O => \N__4566\,
            I => counter_3_1_cry_26
        );

    \I__979\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4559\
        );

    \I__978\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4556\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4559\,
            I => \counter_3Z0Z_28\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4556\,
            I => \counter_3Z0Z_28\
        );

    \I__975\ : InMux
    port map (
            O => \N__4551\,
            I => counter_3_1_cry_27
        );

    \I__974\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4544\
        );

    \I__973\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4541\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4544\,
            I => \counter_3Z0Z_29\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4541\,
            I => \counter_3Z0Z_29\
        );

    \I__970\ : InMux
    port map (
            O => \N__4536\,
            I => counter_3_1_cry_28
        );

    \I__969\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4529\
        );

    \I__968\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4526\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4529\,
            I => \counter_3Z0Z_30\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4526\,
            I => \counter_3Z0Z_30\
        );

    \I__965\ : InMux
    port map (
            O => \N__4521\,
            I => counter_3_1_cry_29
        );

    \I__964\ : InMux
    port map (
            O => \N__4518\,
            I => counter_3_1_cry_30
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__4515\,
            I => \N__4511\
        );

    \I__962\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4508\
        );

    \I__961\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4505\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4508\,
            I => \counter_3Z0Z_31\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4505\,
            I => \counter_3Z0Z_31\
        );

    \I__958\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4497\,
            I => \N__4494\
        );

    \I__956\ : Odrv12
    port map (
            O => \N__4494\,
            I => \counter_3_1_cry_2_THRU_CO\
        );

    \I__955\ : InMux
    port map (
            O => \N__4491\,
            I => \N__4488\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4488\,
            I => \N__4481\
        );

    \I__953\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4478\
        );

    \I__952\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4471\
        );

    \I__951\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4471\
        );

    \I__950\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4471\
        );

    \I__949\ : Span4Mux_h
    port map (
            O => \N__4481\,
            I => \N__4466\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4463\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4471\,
            I => \N__4460\
        );

    \I__946\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4455\
        );

    \I__945\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4455\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__4466\,
            I => \un4_counter_3_7_THRU_CO\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__4463\,
            I => \un4_counter_3_7_THRU_CO\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__4460\,
            I => \un4_counter_3_7_THRU_CO\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4455\,
            I => \un4_counter_3_7_THRU_CO\
        );

    \I__940\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4442\
        );

    \I__939\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4438\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4442\,
            I => \N__4435\
        );

    \I__937\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4432\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4427\
        );

    \I__935\ : Span4Mux_s0_h
    port map (
            O => \N__4435\,
            I => \N__4427\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4432\,
            I => \counter_3Z0Z_3\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__4427\,
            I => \counter_3Z0Z_3\
        );

    \I__932\ : ClkMux
    port map (
            O => \N__4422\,
            I => \N__4356\
        );

    \I__931\ : ClkMux
    port map (
            O => \N__4421\,
            I => \N__4356\
        );

    \I__930\ : ClkMux
    port map (
            O => \N__4420\,
            I => \N__4356\
        );

    \I__929\ : ClkMux
    port map (
            O => \N__4419\,
            I => \N__4356\
        );

    \I__928\ : ClkMux
    port map (
            O => \N__4418\,
            I => \N__4356\
        );

    \I__927\ : ClkMux
    port map (
            O => \N__4417\,
            I => \N__4356\
        );

    \I__926\ : ClkMux
    port map (
            O => \N__4416\,
            I => \N__4356\
        );

    \I__925\ : ClkMux
    port map (
            O => \N__4415\,
            I => \N__4356\
        );

    \I__924\ : ClkMux
    port map (
            O => \N__4414\,
            I => \N__4356\
        );

    \I__923\ : ClkMux
    port map (
            O => \N__4413\,
            I => \N__4356\
        );

    \I__922\ : ClkMux
    port map (
            O => \N__4412\,
            I => \N__4356\
        );

    \I__921\ : ClkMux
    port map (
            O => \N__4411\,
            I => \N__4356\
        );

    \I__920\ : ClkMux
    port map (
            O => \N__4410\,
            I => \N__4356\
        );

    \I__919\ : ClkMux
    port map (
            O => \N__4409\,
            I => \N__4356\
        );

    \I__918\ : ClkMux
    port map (
            O => \N__4408\,
            I => \N__4356\
        );

    \I__917\ : ClkMux
    port map (
            O => \N__4407\,
            I => \N__4356\
        );

    \I__916\ : ClkMux
    port map (
            O => \N__4406\,
            I => \N__4356\
        );

    \I__915\ : ClkMux
    port map (
            O => \N__4405\,
            I => \N__4356\
        );

    \I__914\ : ClkMux
    port map (
            O => \N__4404\,
            I => \N__4356\
        );

    \I__913\ : ClkMux
    port map (
            O => \N__4403\,
            I => \N__4356\
        );

    \I__912\ : ClkMux
    port map (
            O => \N__4402\,
            I => \N__4356\
        );

    \I__911\ : ClkMux
    port map (
            O => \N__4401\,
            I => \N__4356\
        );

    \I__910\ : GlobalMux
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__909\ : gio2CtrlBuf
    port map (
            O => \N__4353\,
            I => \CLK_27mhz_0_0_c_g\
        );

    \I__908\ : CEMux
    port map (
            O => \N__4350\,
            I => \N__4326\
        );

    \I__907\ : CEMux
    port map (
            O => \N__4349\,
            I => \N__4326\
        );

    \I__906\ : CEMux
    port map (
            O => \N__4348\,
            I => \N__4326\
        );

    \I__905\ : CEMux
    port map (
            O => \N__4347\,
            I => \N__4326\
        );

    \I__904\ : CEMux
    port map (
            O => \N__4346\,
            I => \N__4326\
        );

    \I__903\ : CEMux
    port map (
            O => \N__4345\,
            I => \N__4326\
        );

    \I__902\ : CEMux
    port map (
            O => \N__4344\,
            I => \N__4326\
        );

    \I__901\ : CEMux
    port map (
            O => \N__4343\,
            I => \N__4326\
        );

    \I__900\ : GlobalMux
    port map (
            O => \N__4326\,
            I => \N__4323\
        );

    \I__899\ : gio2CtrlBuf
    port map (
            O => \N__4323\,
            I => \N_67_g\
        );

    \I__898\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4316\
        );

    \I__897\ : InMux
    port map (
            O => \N__4319\,
            I => \N__4313\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4316\,
            I => \counter_3Z0Z_17\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4313\,
            I => \counter_3Z0Z_17\
        );

    \I__894\ : InMux
    port map (
            O => \N__4308\,
            I => \bfn_12_9_0_\
        );

    \I__893\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4301\
        );

    \I__892\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4298\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4301\,
            I => \counter_3Z0Z_18\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4298\,
            I => \counter_3Z0Z_18\
        );

    \I__889\ : InMux
    port map (
            O => \N__4293\,
            I => counter_3_1_cry_17
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__4290\,
            I => \N__4286\
        );

    \I__887\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4283\
        );

    \I__886\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4280\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4283\,
            I => \counter_3Z0Z_19\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4280\,
            I => \counter_3Z0Z_19\
        );

    \I__883\ : InMux
    port map (
            O => \N__4275\,
            I => counter_3_1_cry_18
        );

    \I__882\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4268\
        );

    \I__881\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4265\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4268\,
            I => \counter_3Z0Z_20\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4265\,
            I => \counter_3Z0Z_20\
        );

    \I__878\ : InMux
    port map (
            O => \N__4260\,
            I => counter_3_1_cry_19
        );

    \I__877\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4253\
        );

    \I__876\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4250\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4253\,
            I => \counter_3Z0Z_21\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4250\,
            I => \counter_3Z0Z_21\
        );

    \I__873\ : InMux
    port map (
            O => \N__4245\,
            I => counter_3_1_cry_20
        );

    \I__872\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4238\
        );

    \I__871\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4235\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4238\,
            I => \counter_3Z0Z_22\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4235\,
            I => \counter_3Z0Z_22\
        );

    \I__868\ : InMux
    port map (
            O => \N__4230\,
            I => counter_3_1_cry_21
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__4227\,
            I => \N__4223\
        );

    \I__866\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4220\
        );

    \I__865\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4217\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4220\,
            I => \counter_3Z0Z_23\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4217\,
            I => \counter_3Z0Z_23\
        );

    \I__862\ : InMux
    port map (
            O => \N__4212\,
            I => counter_3_1_cry_22
        );

    \I__861\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4205\
        );

    \I__860\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4202\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4205\,
            I => \counter_3Z0Z_24\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4202\,
            I => \counter_3Z0Z_24\
        );

    \I__857\ : InMux
    port map (
            O => \N__4197\,
            I => counter_3_1_cry_23
        );

    \I__856\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4190\
        );

    \I__855\ : InMux
    port map (
            O => \N__4193\,
            I => \N__4187\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4190\,
            I => \counter_3Z0Z_9\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4187\,
            I => \counter_3Z0Z_9\
        );

    \I__852\ : InMux
    port map (
            O => \N__4182\,
            I => \bfn_12_8_0_\
        );

    \I__851\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4175\
        );

    \I__850\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4172\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4175\,
            I => \N__4169\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4172\,
            I => \counter_3Z0Z_10\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__4169\,
            I => \counter_3Z0Z_10\
        );

    \I__846\ : InMux
    port map (
            O => \N__4164\,
            I => counter_3_1_cry_9
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__4161\,
            I => \N__4157\
        );

    \I__844\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4154\
        );

    \I__843\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4151\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4154\,
            I => \counter_3Z0Z_11\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4151\,
            I => \counter_3Z0Z_11\
        );

    \I__840\ : InMux
    port map (
            O => \N__4146\,
            I => counter_3_1_cry_10
        );

    \I__839\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4139\
        );

    \I__838\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4136\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4139\,
            I => \counter_3Z0Z_12\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4136\,
            I => \counter_3Z0Z_12\
        );

    \I__835\ : InMux
    port map (
            O => \N__4131\,
            I => counter_3_1_cry_11
        );

    \I__834\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4124\
        );

    \I__833\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4121\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4124\,
            I => \counter_3Z0Z_13\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4121\,
            I => \counter_3Z0Z_13\
        );

    \I__830\ : InMux
    port map (
            O => \N__4116\,
            I => counter_3_1_cry_12
        );

    \I__829\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4109\
        );

    \I__828\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4106\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4109\,
            I => \counter_3Z0Z_14\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4106\,
            I => \counter_3Z0Z_14\
        );

    \I__825\ : InMux
    port map (
            O => \N__4101\,
            I => counter_3_1_cry_13
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__823\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4091\
        );

    \I__822\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4088\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4091\,
            I => \N__4085\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4088\,
            I => \counter_3Z0Z_15\
        );

    \I__819\ : Odrv4
    port map (
            O => \N__4085\,
            I => \counter_3Z0Z_15\
        );

    \I__818\ : InMux
    port map (
            O => \N__4080\,
            I => counter_3_1_cry_14
        );

    \I__817\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4073\
        );

    \I__816\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4070\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4073\,
            I => \counter_3Z0Z_16\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4070\,
            I => \counter_3Z0Z_16\
        );

    \I__813\ : InMux
    port map (
            O => \N__4065\,
            I => counter_3_1_cry_15
        );

    \I__812\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4057\
        );

    \I__811\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4054\
        );

    \I__810\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4051\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4057\,
            I => \N__4048\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4054\,
            I => \counter_3Z0Z_1\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4051\,
            I => \counter_3Z0Z_1\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__4048\,
            I => \counter_3Z0Z_1\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4041\,
            I => \N__4037\
        );

    \I__804\ : InMux
    port map (
            O => \N__4040\,
            I => \N__4034\
        );

    \I__803\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4031\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4034\,
            I => \N__4026\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4031\,
            I => \N__4023\
        );

    \I__800\ : InMux
    port map (
            O => \N__4030\,
            I => \N__4020\
        );

    \I__799\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4017\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__4026\,
            I => \N__4010\
        );

    \I__797\ : Span4Mux_s0_h
    port map (
            O => \N__4023\,
            I => \N__4010\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4020\,
            I => \N__4010\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4017\,
            I => \counter_3Z0Z_0\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__4010\,
            I => \counter_3Z0Z_0\
        );

    \I__793\ : InMux
    port map (
            O => \N__4005\,
            I => \N__4001\
        );

    \I__792\ : InMux
    port map (
            O => \N__4004\,
            I => \N__3998\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4001\,
            I => \counter_3Z0Z_2\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3998\,
            I => \counter_3Z0Z_2\
        );

    \I__789\ : InMux
    port map (
            O => \N__3993\,
            I => counter_3_1_cry_1
        );

    \I__788\ : InMux
    port map (
            O => \N__3990\,
            I => counter_3_1_cry_2
        );

    \I__787\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3983\
        );

    \I__786\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3979\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3983\,
            I => \N__3976\
        );

    \I__784\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3973\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__3979\,
            I => \counter_3Z0Z_4\
        );

    \I__782\ : Odrv4
    port map (
            O => \N__3976\,
            I => \counter_3Z0Z_4\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3973\,
            I => \counter_3Z0Z_4\
        );

    \I__780\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3963\,
            I => \N__3960\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__3960\,
            I => \counter_3_1_cry_3_THRU_CO\
        );

    \I__777\ : InMux
    port map (
            O => \N__3957\,
            I => counter_3_1_cry_3
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__775\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3946\
        );

    \I__774\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3943\
        );

    \I__773\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3940\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__3946\,
            I => \N__3937\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3943\,
            I => \counter_3Z0Z_5\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3940\,
            I => \counter_3Z0Z_5\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__3937\,
            I => \counter_3Z0Z_5\
        );

    \I__768\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__3927\,
            I => \counter_3_1_cry_4_THRU_CO\
        );

    \I__766\ : InMux
    port map (
            O => \N__3924\,
            I => counter_3_1_cry_4
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__3921\,
            I => \N__3917\
        );

    \I__764\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3913\
        );

    \I__763\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3910\
        );

    \I__762\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3907\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3913\,
            I => \counter_3Z0Z_6\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3910\,
            I => \counter_3Z0Z_6\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3907\,
            I => \counter_3Z0Z_6\
        );

    \I__758\ : InMux
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3897\,
            I => \counter_3_1_cry_5_THRU_CO\
        );

    \I__756\ : InMux
    port map (
            O => \N__3894\,
            I => counter_3_1_cry_5
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__3891\,
            I => \N__3887\
        );

    \I__754\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3883\
        );

    \I__753\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3880\
        );

    \I__752\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3877\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3883\,
            I => \N__3874\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3880\,
            I => \N__3871\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3877\,
            I => \counter_3Z0Z_7\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__3874\,
            I => \counter_3Z0Z_7\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__3871\,
            I => \counter_3Z0Z_7\
        );

    \I__746\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3861\,
            I => \N__3858\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__3858\,
            I => \counter_3_1_cry_6_THRU_CO\
        );

    \I__743\ : InMux
    port map (
            O => \N__3855\,
            I => counter_3_1_cry_6
        );

    \I__742\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3848\
        );

    \I__741\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3845\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3848\,
            I => \counter_3Z0Z_8\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3845\,
            I => \counter_3Z0Z_8\
        );

    \I__738\ : InMux
    port map (
            O => \N__3840\,
            I => counter_3_1_cry_7
        );

    \I__737\ : InMux
    port map (
            O => \N__3837\,
            I => \bfn_11_9_0_\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__735\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3828\,
            I => un4_counter_3_7_and
        );

    \I__733\ : InMux
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3822\,
            I => un4_counter_3_5_and
        );

    \I__731\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3816\,
            I => un4_counter_3_4_and
        );

    \I__729\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3810\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3810\,
            I => un4_counter_3_0_and
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__3807\,
            I => \N__3804\
        );

    \I__726\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3801\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3801\,
            I => un4_counter_3_6_and
        );

    \I__724\ : InMux
    port map (
            O => \N__3798\,
            I => \N__3795\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3795\,
            I => un4_counter_3_1_and
        );

    \I__722\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3789\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3789\,
            I => un4_counter_3_2_and
        );

    \I__720\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3783\,
            I => un4_counter_3_3_and
        );

    \I__718\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3777\,
            I => \clk_2Hz_cnv_m3_e_1\
        );

    \I__716\ : IoInMux
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3771\,
            I => \N__3767\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__3770\,
            I => \N__3764\
        );

    \I__713\ : Span12Mux_s7_v
    port map (
            O => \N__3767\,
            I => \N__3761\
        );

    \I__712\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3758\
        );

    \I__711\ : Odrv12
    port map (
            O => \N__3761\,
            I => \clk_2Hz_c\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3758\,
            I => \clk_2Hz_c\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__3753\,
            I => \N__3750\
        );

    \I__708\ : InMux
    port map (
            O => \N__3750\,
            I => \N__3743\
        );

    \I__707\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3743\
        );

    \I__706\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3740\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3743\,
            I => \clk_1Khz_i\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3740\,
            I => \clk_1Khz_i\
        );

    \I__703\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3726\
        );

    \I__702\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3726\
        );

    \I__701\ : InMux
    port map (
            O => \N__3733\,
            I => \N__3723\
        );

    \I__700\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3718\
        );

    \I__699\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3718\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3726\,
            I => \clk_1MHz_i\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3723\,
            I => \clk_1MHz_i\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3718\,
            I => \clk_1MHz_i\
        );

    \I__695\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3701\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__3710\,
            I => \N__3697\
        );

    \I__693\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3694\
        );

    \I__692\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3683\
        );

    \I__691\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3683\
        );

    \I__690\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3683\
        );

    \I__689\ : InMux
    port map (
            O => \N__3705\,
            I => \N__3683\
        );

    \I__688\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3683\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3701\,
            I => \N__3680\
        );

    \I__686\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3677\
        );

    \I__685\ : InMux
    port map (
            O => \N__3697\,
            I => \N__3674\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3694\,
            I => \N__3671\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3683\,
            I => \N__3666\
        );

    \I__682\ : Span4Mux_h
    port map (
            O => \N__3680\,
            I => \N__3666\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3677\,
            I => \N__3661\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3674\,
            I => \N__3661\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__3671\,
            I => \un4_counter_2_7_THRU_CO\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__3666\,
            I => \un4_counter_2_7_THRU_CO\
        );

    \I__677\ : Odrv12
    port map (
            O => \N__3661\,
            I => \un4_counter_2_7_THRU_CO\
        );

    \I__676\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3641\
        );

    \I__675\ : InMux
    port map (
            O => \N__3653\,
            I => \N__3641\
        );

    \I__674\ : InMux
    port map (
            O => \N__3652\,
            I => \N__3641\
        );

    \I__673\ : InMux
    port map (
            O => \N__3651\,
            I => \N__3641\
        );

    \I__672\ : InMux
    port map (
            O => \N__3650\,
            I => \N__3635\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3641\,
            I => \N__3632\
        );

    \I__670\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3627\
        );

    \I__669\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3627\
        );

    \I__668\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3624\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3635\,
            I => \un4_counter_1_7_THRU_CO\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__3632\,
            I => \un4_counter_1_7_THRU_CO\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3627\,
            I => \un4_counter_1_7_THRU_CO\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3624\,
            I => \un4_counter_1_7_THRU_CO\
        );

    \I__663\ : IoInMux
    port map (
            O => \N__3615\,
            I => \N__3612\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__661\ : Odrv12
    port map (
            O => \N__3609\,
            I => \clk_1Khz_RNIDQNNZ0\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__659\ : InMux
    port map (
            O => \N__3603\,
            I => \N__3600\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__657\ : Span4Mux_v
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__3594\,
            I => un4_counter_1_1_and
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__654\ : InMux
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__652\ : Span4Mux_v
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__3579\,
            I => un4_counter_1_2_and
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__649\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3570\,
            I => \N__3567\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__3567\,
            I => \N__3564\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__3564\,
            I => un4_counter_1_3_and
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__3561\,
            I => \N__3558\
        );

    \I__644\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3555\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3555\,
            I => \N__3552\
        );

    \I__642\ : Span4Mux_h
    port map (
            O => \N__3552\,
            I => \N__3549\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__3549\,
            I => un4_counter_1_4_and
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3546\,
            I => \N__3543\
        );

    \I__639\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3540\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3540\,
            I => \N__3537\
        );

    \I__637\ : Span4Mux_h
    port map (
            O => \N__3537\,
            I => \N__3534\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__3534\,
            I => un4_counter_1_5_and
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__3531\,
            I => \N__3528\
        );

    \I__634\ : InMux
    port map (
            O => \N__3528\,
            I => \N__3525\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3525\,
            I => \N__3522\
        );

    \I__632\ : Span4Mux_h
    port map (
            O => \N__3522\,
            I => \N__3519\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3519\,
            I => un4_counter_1_6_and
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__3516\,
            I => \N__3513\
        );

    \I__629\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3510\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3510\,
            I => \N__3507\
        );

    \I__627\ : Span4Mux_h
    port map (
            O => \N__3507\,
            I => \N__3504\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__3504\,
            I => un4_counter_1_7_and
        );

    \I__625\ : InMux
    port map (
            O => \N__3501\,
            I => \bfn_5_7_0_\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__3498\,
            I => \un4_counter_1_7_THRU_CO_cascade_\
        );

    \I__623\ : IoInMux
    port map (
            O => \N__3495\,
            I => \N__3492\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3492\,
            I => \N__3489\
        );

    \I__621\ : Span4Mux_s0_h
    port map (
            O => \N__3489\,
            I => \N__3486\
        );

    \I__620\ : Span4Mux_h
    port map (
            O => \N__3486\,
            I => \N__3483\
        );

    \I__619\ : Odrv4
    port map (
            O => \N__3483\,
            I => \clk_1Khz_cnv_0\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__3480\,
            I => \N__3476\
        );

    \I__617\ : InMux
    port map (
            O => \N__3479\,
            I => \N__3473\
        );

    \I__616\ : InMux
    port map (
            O => \N__3476\,
            I => \N__3470\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3473\,
            I => \counter_2Z0Z_30\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3470\,
            I => \counter_2Z0Z_30\
        );

    \I__613\ : InMux
    port map (
            O => \N__3465\,
            I => counter_2_1_cry_29
        );

    \I__612\ : InMux
    port map (
            O => \N__3462\,
            I => counter_2_1_cry_30
        );

    \I__611\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3455\
        );

    \I__610\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3452\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3455\,
            I => \counter_2Z0Z_31\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3452\,
            I => \counter_2Z0Z_31\
        );

    \I__607\ : CEMux
    port map (
            O => \N__3447\,
            I => \N__3429\
        );

    \I__606\ : CEMux
    port map (
            O => \N__3446\,
            I => \N__3429\
        );

    \I__605\ : CEMux
    port map (
            O => \N__3445\,
            I => \N__3429\
        );

    \I__604\ : CEMux
    port map (
            O => \N__3444\,
            I => \N__3429\
        );

    \I__603\ : CEMux
    port map (
            O => \N__3443\,
            I => \N__3429\
        );

    \I__602\ : CEMux
    port map (
            O => \N__3442\,
            I => \N__3429\
        );

    \I__601\ : GlobalMux
    port map (
            O => \N__3429\,
            I => \N__3426\
        );

    \I__600\ : gio2CtrlBuf
    port map (
            O => \N__3426\,
            I => \clk_1Khz_cnv_0_g\
        );

    \I__599\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3420\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3417\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__3417\,
            I => \N__3414\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__3414\,
            I => \counter_1_1_cry_2_THRU_CO\
        );

    \I__595\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3408\,
            I => \N__3405\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__592\ : Odrv4
    port map (
            O => \N__3402\,
            I => \counter_1_1_cry_1_THRU_CO\
        );

    \I__591\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3396\,
            I => \N__3392\
        );

    \I__589\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3388\
        );

    \I__588\ : Span4Mux_s3_h
    port map (
            O => \N__3392\,
            I => \N__3385\
        );

    \I__587\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3382\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3388\,
            I => \counter_1Z0Z_2\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__3385\,
            I => \counter_1Z0Z_2\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3382\,
            I => \counter_1Z0Z_2\
        );

    \I__583\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3372\,
            I => \N__3369\
        );

    \I__581\ : Span4Mux_s3_h
    port map (
            O => \N__3369\,
            I => \N__3364\
        );

    \I__580\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3359\
        );

    \I__579\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3359\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__3364\,
            I => \counter_1Z0Z_3\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3359\,
            I => \counter_1Z0Z_3\
        );

    \I__576\ : InMux
    port map (
            O => \N__3354\,
            I => \N__3351\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3351\,
            I => \N__3347\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__3350\,
            I => \N__3342\
        );

    \I__573\ : Span4Mux_s3_h
    port map (
            O => \N__3347\,
            I => \N__3339\
        );

    \I__572\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3332\
        );

    \I__571\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3332\
        );

    \I__570\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3332\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__3339\,
            I => \counter_1Z0Z_0\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3332\,
            I => \counter_1Z0Z_0\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__566\ : InMux
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3321\,
            I => \N__3317\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3320\,
            I => \N__3314\
        );

    \I__563\ : Span12Mux_s4_v
    port map (
            O => \N__3317\,
            I => \N__3310\
        );

    \I__562\ : InMux
    port map (
            O => \N__3314\,
            I => \N__3305\
        );

    \I__561\ : InMux
    port map (
            O => \N__3313\,
            I => \N__3305\
        );

    \I__560\ : Odrv12
    port map (
            O => \N__3310\,
            I => \counter_1Z0Z_1\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3305\,
            I => \counter_1Z0Z_1\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__3300\,
            I => \N__3297\
        );

    \I__557\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3294\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3294\,
            I => un4_counter_1_0_and
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__3291\,
            I => \N__3287\
        );

    \I__554\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3284\
        );

    \I__553\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3281\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3284\,
            I => \counter_2Z0Z_21\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3281\,
            I => \counter_2Z0Z_21\
        );

    \I__550\ : InMux
    port map (
            O => \N__3276\,
            I => counter_2_1_cry_20
        );

    \I__549\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3269\
        );

    \I__548\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3266\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3269\,
            I => \counter_2Z0Z_22\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3266\,
            I => \counter_2Z0Z_22\
        );

    \I__545\ : InMux
    port map (
            O => \N__3261\,
            I => counter_2_1_cry_21
        );

    \I__544\ : InMux
    port map (
            O => \N__3258\,
            I => \N__3254\
        );

    \I__543\ : InMux
    port map (
            O => \N__3257\,
            I => \N__3251\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3254\,
            I => \counter_2Z0Z_23\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3251\,
            I => \counter_2Z0Z_23\
        );

    \I__540\ : InMux
    port map (
            O => \N__3246\,
            I => counter_2_1_cry_22
        );

    \I__539\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3239\
        );

    \I__538\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3236\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3239\,
            I => \counter_2Z0Z_24\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3236\,
            I => \counter_2Z0Z_24\
        );

    \I__535\ : InMux
    port map (
            O => \N__3231\,
            I => counter_2_1_cry_23
        );

    \I__534\ : InMux
    port map (
            O => \N__3228\,
            I => \N__3224\
        );

    \I__533\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3221\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3224\,
            I => \counter_2Z0Z_25\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3221\,
            I => \counter_2Z0Z_25\
        );

    \I__530\ : InMux
    port map (
            O => \N__3216\,
            I => \bfn_2_10_0_\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__3213\,
            I => \N__3209\
        );

    \I__528\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3206\
        );

    \I__527\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3203\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3206\,
            I => \counter_2Z0Z_26\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3203\,
            I => \counter_2Z0Z_26\
        );

    \I__524\ : InMux
    port map (
            O => \N__3198\,
            I => counter_2_1_cry_25
        );

    \I__523\ : InMux
    port map (
            O => \N__3195\,
            I => \N__3191\
        );

    \I__522\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3188\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3191\,
            I => \counter_2Z0Z_27\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3188\,
            I => \counter_2Z0Z_27\
        );

    \I__519\ : InMux
    port map (
            O => \N__3183\,
            I => counter_2_1_cry_26
        );

    \I__518\ : InMux
    port map (
            O => \N__3180\,
            I => \N__3176\
        );

    \I__517\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3173\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3176\,
            I => \counter_2Z0Z_28\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3173\,
            I => \counter_2Z0Z_28\
        );

    \I__514\ : InMux
    port map (
            O => \N__3168\,
            I => counter_2_1_cry_27
        );

    \I__513\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3161\
        );

    \I__512\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3158\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3161\,
            I => \counter_2Z0Z_29\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3158\,
            I => \counter_2Z0Z_29\
        );

    \I__509\ : InMux
    port map (
            O => \N__3153\,
            I => counter_2_1_cry_28
        );

    \I__508\ : InMux
    port map (
            O => \N__3150\,
            I => \N__3146\
        );

    \I__507\ : InMux
    port map (
            O => \N__3149\,
            I => \N__3143\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3146\,
            I => \counter_2Z0Z_13\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3143\,
            I => \counter_2Z0Z_13\
        );

    \I__504\ : InMux
    port map (
            O => \N__3138\,
            I => counter_2_1_cry_12
        );

    \I__503\ : CascadeMux
    port map (
            O => \N__3135\,
            I => \N__3131\
        );

    \I__502\ : InMux
    port map (
            O => \N__3134\,
            I => \N__3128\
        );

    \I__501\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3125\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3128\,
            I => \counter_2Z0Z_14\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3125\,
            I => \counter_2Z0Z_14\
        );

    \I__498\ : InMux
    port map (
            O => \N__3120\,
            I => counter_2_1_cry_13
        );

    \I__497\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3113\
        );

    \I__496\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3110\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3113\,
            I => \counter_2Z0Z_15\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3110\,
            I => \counter_2Z0Z_15\
        );

    \I__493\ : InMux
    port map (
            O => \N__3105\,
            I => counter_2_1_cry_14
        );

    \I__492\ : InMux
    port map (
            O => \N__3102\,
            I => \N__3098\
        );

    \I__491\ : InMux
    port map (
            O => \N__3101\,
            I => \N__3095\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3098\,
            I => \counter_2Z0Z_16\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3095\,
            I => \counter_2Z0Z_16\
        );

    \I__488\ : InMux
    port map (
            O => \N__3090\,
            I => counter_2_1_cry_15
        );

    \I__487\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3083\
        );

    \I__486\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3080\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3083\,
            I => \counter_2Z0Z_17\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3080\,
            I => \counter_2Z0Z_17\
        );

    \I__483\ : InMux
    port map (
            O => \N__3075\,
            I => \bfn_2_9_0_\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__3072\,
            I => \N__3069\
        );

    \I__481\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3065\
        );

    \I__480\ : InMux
    port map (
            O => \N__3068\,
            I => \N__3062\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3065\,
            I => \N__3059\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3062\,
            I => \counter_2Z0Z_18\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__3059\,
            I => \counter_2Z0Z_18\
        );

    \I__476\ : InMux
    port map (
            O => \N__3054\,
            I => counter_2_1_cry_17
        );

    \I__475\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3047\
        );

    \I__474\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3044\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3047\,
            I => \N__3041\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3044\,
            I => \counter_2Z0Z_19\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__3041\,
            I => \counter_2Z0Z_19\
        );

    \I__470\ : InMux
    port map (
            O => \N__3036\,
            I => counter_2_1_cry_18
        );

    \I__469\ : InMux
    port map (
            O => \N__3033\,
            I => \N__3029\
        );

    \I__468\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3026\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3029\,
            I => \counter_2Z0Z_20\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3026\,
            I => \counter_2Z0Z_20\
        );

    \I__465\ : InMux
    port map (
            O => \N__3021\,
            I => counter_2_1_cry_19
        );

    \I__464\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3014\
        );

    \I__463\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3010\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3014\,
            I => \N__3007\
        );

    \I__461\ : InMux
    port map (
            O => \N__3013\,
            I => \N__3004\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3010\,
            I => \counter_2Z0Z_5\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__3007\,
            I => \counter_2Z0Z_5\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3004\,
            I => \counter_2Z0Z_5\
        );

    \I__457\ : InMux
    port map (
            O => \N__2997\,
            I => \N__2994\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2994\,
            I => \N__2991\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__2991\,
            I => \counter_2_1_cry_4_THRU_CO\
        );

    \I__454\ : InMux
    port map (
            O => \N__2988\,
            I => counter_2_1_cry_4
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__2985\,
            I => \N__2980\
        );

    \I__452\ : InMux
    port map (
            O => \N__2984\,
            I => \N__2977\
        );

    \I__451\ : InMux
    port map (
            O => \N__2983\,
            I => \N__2974\
        );

    \I__450\ : InMux
    port map (
            O => \N__2980\,
            I => \N__2971\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2977\,
            I => \counter_2Z0Z_6\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2974\,
            I => \counter_2Z0Z_6\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2971\,
            I => \counter_2Z0Z_6\
        );

    \I__446\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2961\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2961\,
            I => \counter_2_1_cry_5_THRU_CO\
        );

    \I__444\ : InMux
    port map (
            O => \N__2958\,
            I => counter_2_1_cry_5
        );

    \I__443\ : InMux
    port map (
            O => \N__2955\,
            I => \N__2950\
        );

    \I__442\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2947\
        );

    \I__441\ : InMux
    port map (
            O => \N__2953\,
            I => \N__2944\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2950\,
            I => \counter_2Z0Z_7\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2947\,
            I => \counter_2Z0Z_7\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2944\,
            I => \counter_2Z0Z_7\
        );

    \I__437\ : InMux
    port map (
            O => \N__2937\,
            I => \N__2934\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2934\,
            I => \counter_2_1_cry_6_THRU_CO\
        );

    \I__435\ : InMux
    port map (
            O => \N__2931\,
            I => counter_2_1_cry_6
        );

    \I__434\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2923\
        );

    \I__433\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2920\
        );

    \I__432\ : InMux
    port map (
            O => \N__2926\,
            I => \N__2917\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2923\,
            I => \counter_2Z0Z_8\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2920\,
            I => \counter_2Z0Z_8\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2917\,
            I => \counter_2Z0Z_8\
        );

    \I__428\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2907\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2907\,
            I => \counter_2_1_cry_7_THRU_CO\
        );

    \I__426\ : InMux
    port map (
            O => \N__2904\,
            I => counter_2_1_cry_7
        );

    \I__425\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2897\
        );

    \I__424\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2894\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2897\,
            I => \counter_2Z0Z_9\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2894\,
            I => \counter_2Z0Z_9\
        );

    \I__421\ : InMux
    port map (
            O => \N__2889\,
            I => \bfn_2_8_0_\
        );

    \I__420\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2882\
        );

    \I__419\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2879\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2882\,
            I => \counter_2Z0Z_10\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2879\,
            I => \counter_2Z0Z_10\
        );

    \I__416\ : InMux
    port map (
            O => \N__2874\,
            I => counter_2_1_cry_9
        );

    \I__415\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2867\
        );

    \I__414\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2864\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2867\,
            I => \counter_2Z0Z_11\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2864\,
            I => \counter_2Z0Z_11\
        );

    \I__411\ : InMux
    port map (
            O => \N__2859\,
            I => counter_2_1_cry_10
        );

    \I__410\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2852\
        );

    \I__409\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2849\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2852\,
            I => \counter_2Z0Z_12\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2849\,
            I => \counter_2Z0Z_12\
        );

    \I__406\ : InMux
    port map (
            O => \N__2844\,
            I => counter_2_1_cry_11
        );

    \I__405\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2833\
        );

    \I__404\ : InMux
    port map (
            O => \N__2840\,
            I => \N__2833\
        );

    \I__403\ : InMux
    port map (
            O => \N__2839\,
            I => \N__2830\
        );

    \I__402\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2827\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2833\,
            I => \counter_2Z0Z_0\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2830\,
            I => \counter_2Z0Z_0\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2827\,
            I => \counter_2Z0Z_0\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__2820\,
            I => \N__2815\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__2819\,
            I => \N__2812\
        );

    \I__396\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2809\
        );

    \I__395\ : InMux
    port map (
            O => \N__2815\,
            I => \N__2806\
        );

    \I__394\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2803\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2809\,
            I => \counter_2Z0Z_1\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2806\,
            I => \counter_2Z0Z_1\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2803\,
            I => \counter_2Z0Z_1\
        );

    \I__390\ : InMux
    port map (
            O => \N__2796\,
            I => \N__2791\
        );

    \I__389\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2788\
        );

    \I__388\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2785\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2791\,
            I => \counter_2Z0Z_2\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2788\,
            I => \counter_2Z0Z_2\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2785\,
            I => \counter_2Z0Z_2\
        );

    \I__384\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2775\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2775\,
            I => \counter_2_1_cry_1_THRU_CO\
        );

    \I__382\ : InMux
    port map (
            O => \N__2772\,
            I => counter_2_1_cry_1
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__2769\,
            I => \N__2765\
        );

    \I__380\ : InMux
    port map (
            O => \N__2768\,
            I => \N__2762\
        );

    \I__379\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2759\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2762\,
            I => \counter_2Z0Z_3\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2759\,
            I => \counter_2Z0Z_3\
        );

    \I__376\ : InMux
    port map (
            O => \N__2754\,
            I => counter_2_1_cry_2
        );

    \I__375\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2746\
        );

    \I__374\ : InMux
    port map (
            O => \N__2750\,
            I => \N__2743\
        );

    \I__373\ : InMux
    port map (
            O => \N__2749\,
            I => \N__2740\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2746\,
            I => \counter_2Z0Z_4\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2743\,
            I => \counter_2Z0Z_4\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2740\,
            I => \counter_2Z0Z_4\
        );

    \I__369\ : CascadeMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__368\ : InMux
    port map (
            O => \N__2730\,
            I => \N__2727\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2727\,
            I => \counter_2_1_cry_3_THRU_CO\
        );

    \I__366\ : InMux
    port map (
            O => \N__2724\,
            I => counter_2_1_cry_3
        );

    \I__365\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2717\
        );

    \I__364\ : InMux
    port map (
            O => \N__2720\,
            I => \N__2714\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2717\,
            I => \counter_1Z0Z_5\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2714\,
            I => \counter_1Z0Z_5\
        );

    \I__361\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2705\
        );

    \I__360\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2702\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2705\,
            I => \counter_1Z0Z_7\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2702\,
            I => \counter_1Z0Z_7\
        );

    \I__357\ : CascadeMux
    port map (
            O => \N__2697\,
            I => \N__2693\
        );

    \I__356\ : InMux
    port map (
            O => \N__2696\,
            I => \N__2690\
        );

    \I__355\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2687\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2690\,
            I => \counter_1Z0Z_6\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2687\,
            I => \counter_1Z0Z_6\
        );

    \I__352\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2678\
        );

    \I__351\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2675\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2678\,
            I => \counter_1Z0Z_4\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2675\,
            I => \counter_1Z0Z_4\
        );

    \I__348\ : InMux
    port map (
            O => \N__2670\,
            I => \N__2666\
        );

    \I__347\ : InMux
    port map (
            O => \N__2669\,
            I => \N__2663\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2666\,
            I => \counter_1Z0Z_8\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2663\,
            I => \counter_1Z0Z_8\
        );

    \I__344\ : InMux
    port map (
            O => \N__2658\,
            I => \N__2654\
        );

    \I__343\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2651\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2654\,
            I => \counter_1Z0Z_10\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2651\,
            I => \counter_1Z0Z_10\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__2646\,
            I => \N__2642\
        );

    \I__339\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2639\
        );

    \I__338\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2636\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2639\,
            I => \counter_1Z0Z_9\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2636\,
            I => \counter_1Z0Z_9\
        );

    \I__335\ : InMux
    port map (
            O => \N__2631\,
            I => \N__2627\
        );

    \I__334\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2624\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2627\,
            I => \counter_1Z0Z_11\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2624\,
            I => \counter_1Z0Z_11\
        );

    \I__331\ : InMux
    port map (
            O => \N__2619\,
            I => \N__2615\
        );

    \I__330\ : InMux
    port map (
            O => \N__2618\,
            I => \N__2612\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2615\,
            I => \counter_1Z0Z_13\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2612\,
            I => \counter_1Z0Z_13\
        );

    \I__327\ : InMux
    port map (
            O => \N__2607\,
            I => \N__2603\
        );

    \I__326\ : InMux
    port map (
            O => \N__2606\,
            I => \N__2600\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2603\,
            I => \counter_1Z0Z_12\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2600\,
            I => \counter_1Z0Z_12\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__2595\,
            I => \N__2591\
        );

    \I__322\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2588\
        );

    \I__321\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2585\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2588\,
            I => \counter_1Z0Z_15\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2585\,
            I => \counter_1Z0Z_15\
        );

    \I__318\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2576\
        );

    \I__317\ : InMux
    port map (
            O => \N__2579\,
            I => \N__2573\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2576\,
            I => \counter_1Z0Z_14\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2573\,
            I => \counter_1Z0Z_14\
        );

    \I__314\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2564\
        );

    \I__313\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2561\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2564\,
            I => \counter_1Z0Z_18\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2561\,
            I => \counter_1Z0Z_18\
        );

    \I__310\ : InMux
    port map (
            O => \N__2556\,
            I => \N__2552\
        );

    \I__309\ : InMux
    port map (
            O => \N__2555\,
            I => \N__2549\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2552\,
            I => \counter_1Z0Z_19\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2549\,
            I => \counter_1Z0Z_19\
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2544\,
            I => \N__2540\
        );

    \I__305\ : InMux
    port map (
            O => \N__2543\,
            I => \N__2537\
        );

    \I__304\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2534\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2537\,
            I => \counter_1Z0Z_17\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2534\,
            I => \counter_1Z0Z_17\
        );

    \I__301\ : InMux
    port map (
            O => \N__2529\,
            I => \N__2525\
        );

    \I__300\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2522\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2525\,
            I => \counter_1Z0Z_16\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2522\,
            I => \counter_1Z0Z_16\
        );

    \I__297\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2513\
        );

    \I__296\ : InMux
    port map (
            O => \N__2516\,
            I => \N__2510\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2513\,
            I => \counter_1Z0Z_20\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2510\,
            I => \counter_1Z0Z_20\
        );

    \I__293\ : InMux
    port map (
            O => \N__2505\,
            I => \N__2501\
        );

    \I__292\ : InMux
    port map (
            O => \N__2504\,
            I => \N__2498\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2501\,
            I => \counter_1Z0Z_21\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2498\,
            I => \counter_1Z0Z_21\
        );

    \I__289\ : CascadeMux
    port map (
            O => \N__2493\,
            I => \N__2489\
        );

    \I__288\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2486\
        );

    \I__287\ : InMux
    port map (
            O => \N__2489\,
            I => \N__2483\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2486\,
            I => \counter_1Z0Z_23\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2483\,
            I => \counter_1Z0Z_23\
        );

    \I__284\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2474\
        );

    \I__283\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2471\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2474\,
            I => \counter_1Z0Z_22\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2471\,
            I => \counter_1Z0Z_22\
        );

    \I__280\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2462\
        );

    \I__279\ : InMux
    port map (
            O => \N__2465\,
            I => \N__2459\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2462\,
            I => \counter_1Z0Z_27\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2459\,
            I => \counter_1Z0Z_27\
        );

    \I__276\ : InMux
    port map (
            O => \N__2454\,
            I => \N__2450\
        );

    \I__275\ : InMux
    port map (
            O => \N__2453\,
            I => \N__2447\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2450\,
            I => \counter_1Z0Z_24\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2447\,
            I => \counter_1Z0Z_24\
        );

    \I__272\ : CascadeMux
    port map (
            O => \N__2442\,
            I => \N__2438\
        );

    \I__271\ : InMux
    port map (
            O => \N__2441\,
            I => \N__2435\
        );

    \I__270\ : InMux
    port map (
            O => \N__2438\,
            I => \N__2432\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2435\,
            I => \counter_1Z0Z_25\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2432\,
            I => \counter_1Z0Z_25\
        );

    \I__267\ : InMux
    port map (
            O => \N__2427\,
            I => \N__2423\
        );

    \I__266\ : InMux
    port map (
            O => \N__2426\,
            I => \N__2420\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2423\,
            I => \counter_1Z0Z_26\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2420\,
            I => \counter_1Z0Z_26\
        );

    \I__263\ : InMux
    port map (
            O => \N__2415\,
            I => \bfn_1_8_0_\
        );

    \I__262\ : CascadeMux
    port map (
            O => \N__2412\,
            I => \N__2409\
        );

    \I__261\ : InMux
    port map (
            O => \N__2409\,
            I => \N__2406\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2406\,
            I => un4_counter_2_5_and
        );

    \I__259\ : CascadeMux
    port map (
            O => \N__2403\,
            I => \N__2400\
        );

    \I__258\ : InMux
    port map (
            O => \N__2400\,
            I => \N__2397\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2397\,
            I => un4_counter_2_4_and
        );

    \I__256\ : CascadeMux
    port map (
            O => \N__2394\,
            I => \N__2391\
        );

    \I__255\ : InMux
    port map (
            O => \N__2391\,
            I => \N__2388\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2388\,
            I => un4_counter_2_2_and
        );

    \I__253\ : CascadeMux
    port map (
            O => \N__2385\,
            I => \N__2382\
        );

    \I__252\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2379\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2379\,
            I => un4_counter_2_3_and
        );

    \I__250\ : CascadeMux
    port map (
            O => \N__2376\,
            I => \N__2373\
        );

    \I__249\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2370\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__2370\,
            I => \N__2367\
        );

    \I__247\ : Odrv4
    port map (
            O => \N__2367\,
            I => un4_counter_2_7_and
        );

    \I__246\ : CascadeMux
    port map (
            O => \N__2364\,
            I => \N__2361\
        );

    \I__245\ : InMux
    port map (
            O => \N__2361\,
            I => \N__2358\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2358\,
            I => \N__2355\
        );

    \I__243\ : Odrv4
    port map (
            O => \N__2355\,
            I => un4_counter_2_6_and
        );

    \I__242\ : InMux
    port map (
            O => \N__2352\,
            I => \N__2349\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2349\,
            I => un4_counter_2_0_and
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__2346\,
            I => \N__2343\
        );

    \I__239\ : InMux
    port map (
            O => \N__2343\,
            I => \N__2340\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2340\,
            I => un4_counter_2_1_and
        );

    \I__237\ : InMux
    port map (
            O => \N__2337\,
            I => counter_1_1_cry_23
        );

    \I__236\ : InMux
    port map (
            O => \N__2334\,
            I => \bfn_1_4_0_\
        );

    \I__235\ : InMux
    port map (
            O => \N__2331\,
            I => counter_1_1_cry_25
        );

    \I__234\ : InMux
    port map (
            O => \N__2328\,
            I => counter_1_1_cry_26
        );

    \I__233\ : InMux
    port map (
            O => \N__2325\,
            I => counter_1_1_cry_27
        );

    \I__232\ : InMux
    port map (
            O => \N__2322\,
            I => counter_1_1_cry_28
        );

    \I__231\ : InMux
    port map (
            O => \N__2319\,
            I => counter_1_1_cry_29
        );

    \I__230\ : InMux
    port map (
            O => \N__2316\,
            I => counter_1_1_cry_30
        );

    \I__229\ : InMux
    port map (
            O => \N__2313\,
            I => \N__2307\
        );

    \I__228\ : InMux
    port map (
            O => \N__2312\,
            I => \N__2307\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2307\,
            I => \counter_1Z0Z_29\
        );

    \I__226\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2298\
        );

    \I__225\ : InMux
    port map (
            O => \N__2303\,
            I => \N__2298\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2298\,
            I => \counter_1Z0Z_28\
        );

    \I__223\ : CascadeMux
    port map (
            O => \N__2295\,
            I => \N__2291\
        );

    \I__222\ : CascadeMux
    port map (
            O => \N__2294\,
            I => \N__2288\
        );

    \I__221\ : InMux
    port map (
            O => \N__2291\,
            I => \N__2283\
        );

    \I__220\ : InMux
    port map (
            O => \N__2288\,
            I => \N__2283\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__2283\,
            I => \counter_1Z0Z_30\
        );

    \I__218\ : InMux
    port map (
            O => \N__2280\,
            I => \N__2274\
        );

    \I__217\ : InMux
    port map (
            O => \N__2279\,
            I => \N__2274\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__2274\,
            I => \counter_1Z0Z_31\
        );

    \I__215\ : InMux
    port map (
            O => \N__2271\,
            I => counter_1_1_cry_14
        );

    \I__214\ : InMux
    port map (
            O => \N__2268\,
            I => counter_1_1_cry_15
        );

    \I__213\ : InMux
    port map (
            O => \N__2265\,
            I => \bfn_1_3_0_\
        );

    \I__212\ : InMux
    port map (
            O => \N__2262\,
            I => counter_1_1_cry_17
        );

    \I__211\ : InMux
    port map (
            O => \N__2259\,
            I => counter_1_1_cry_18
        );

    \I__210\ : InMux
    port map (
            O => \N__2256\,
            I => counter_1_1_cry_19
        );

    \I__209\ : InMux
    port map (
            O => \N__2253\,
            I => counter_1_1_cry_20
        );

    \I__208\ : InMux
    port map (
            O => \N__2250\,
            I => counter_1_1_cry_21
        );

    \I__207\ : InMux
    port map (
            O => \N__2247\,
            I => counter_1_1_cry_22
        );

    \I__206\ : InMux
    port map (
            O => \N__2244\,
            I => counter_1_1_cry_5
        );

    \I__205\ : InMux
    port map (
            O => \N__2241\,
            I => counter_1_1_cry_6
        );

    \I__204\ : InMux
    port map (
            O => \N__2238\,
            I => counter_1_1_cry_7
        );

    \I__203\ : InMux
    port map (
            O => \N__2235\,
            I => \bfn_1_2_0_\
        );

    \I__202\ : InMux
    port map (
            O => \N__2232\,
            I => counter_1_1_cry_9
        );

    \I__201\ : InMux
    port map (
            O => \N__2229\,
            I => counter_1_1_cry_10
        );

    \I__200\ : InMux
    port map (
            O => \N__2226\,
            I => counter_1_1_cry_11
        );

    \I__199\ : InMux
    port map (
            O => \N__2223\,
            I => counter_1_1_cry_12
        );

    \I__198\ : InMux
    port map (
            O => \N__2220\,
            I => counter_1_1_cry_13
        );

    \I__197\ : InMux
    port map (
            O => \N__2217\,
            I => counter_1_1_cry_1
        );

    \I__196\ : InMux
    port map (
            O => \N__2214\,
            I => counter_1_1_cry_2
        );

    \I__195\ : InMux
    port map (
            O => \N__2211\,
            I => counter_1_1_cry_3
        );

    \I__194\ : InMux
    port map (
            O => \N__2208\,
            I => counter_1_1_cry_4
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_counter_3_7,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_counter_2_7,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_counter_1_7,
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_3_1_cry_8,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_3_1_cry_16,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_3_1_cry_24,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_2_1_cry_8,
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_2_1_cry_16,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_2_1_cry_24,
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_1_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_1_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_1_1_cry_8,
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_1_1_cry_16,
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_1_1_cry_24,
            carryinitout => \bfn_1_4_0_\
        );

    \clk_1MHz_RNINCP9_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3495\,
            GLOBALBUFFEROUTPUT => \clk_1Khz_cnv_0_g\
        );

    \clk_1Khz_RNIDQNN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3615\,
            GLOBALBUFFEROUTPUT => \N_67_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \counter_1_1_cry_1_c_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3354\,
            in2 => \N__3327\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_1_0_\,
            carryout => counter_1_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_1_cry_1_THRU_LUT4_0_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3399\,
            in2 => \_gnd_net_\,
            in3 => \N__2217\,
            lcout => \counter_1_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => counter_1_1_cry_1,
            carryout => counter_1_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_1_cry_2_THRU_LUT4_0_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3375\,
            in2 => \_gnd_net_\,
            in3 => \N__2214\,
            lcout => \counter_1_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => counter_1_1_cry_2,
            carryout => counter_1_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_4_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2682\,
            in2 => \_gnd_net_\,
            in3 => \N__2211\,
            lcout => \counter_1Z0Z_4\,
            ltout => OPEN,
            carryin => counter_1_1_cry_3,
            carryout => counter_1_1_cry_4,
            clk => \N__4414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_5_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2721\,
            in2 => \_gnd_net_\,
            in3 => \N__2208\,
            lcout => \counter_1Z0Z_5\,
            ltout => OPEN,
            carryin => counter_1_1_cry_4,
            carryout => counter_1_1_cry_5,
            clk => \N__4414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_6_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2696\,
            in2 => \_gnd_net_\,
            in3 => \N__2244\,
            lcout => \counter_1Z0Z_6\,
            ltout => OPEN,
            carryin => counter_1_1_cry_5,
            carryout => counter_1_1_cry_6,
            clk => \N__4414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_7_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2709\,
            in2 => \_gnd_net_\,
            in3 => \N__2241\,
            lcout => \counter_1Z0Z_7\,
            ltout => OPEN,
            carryin => counter_1_1_cry_6,
            carryout => counter_1_1_cry_7,
            clk => \N__4414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_8_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2670\,
            in2 => \_gnd_net_\,
            in3 => \N__2238\,
            lcout => \counter_1Z0Z_8\,
            ltout => OPEN,
            carryin => counter_1_1_cry_7,
            carryout => counter_1_1_cry_8,
            clk => \N__4414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_9_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2645\,
            in2 => \_gnd_net_\,
            in3 => \N__2235\,
            lcout => \counter_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => counter_1_1_cry_9,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_10_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2658\,
            in2 => \_gnd_net_\,
            in3 => \N__2232\,
            lcout => \counter_1Z0Z_10\,
            ltout => OPEN,
            carryin => counter_1_1_cry_9,
            carryout => counter_1_1_cry_10,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_11_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2631\,
            in2 => \_gnd_net_\,
            in3 => \N__2229\,
            lcout => \counter_1Z0Z_11\,
            ltout => OPEN,
            carryin => counter_1_1_cry_10,
            carryout => counter_1_1_cry_11,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_12_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2607\,
            in2 => \_gnd_net_\,
            in3 => \N__2226\,
            lcout => \counter_1Z0Z_12\,
            ltout => OPEN,
            carryin => counter_1_1_cry_11,
            carryout => counter_1_1_cry_12,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_13_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2619\,
            in2 => \_gnd_net_\,
            in3 => \N__2223\,
            lcout => \counter_1Z0Z_13\,
            ltout => OPEN,
            carryin => counter_1_1_cry_12,
            carryout => counter_1_1_cry_13,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_14_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2580\,
            in2 => \_gnd_net_\,
            in3 => \N__2220\,
            lcout => \counter_1Z0Z_14\,
            ltout => OPEN,
            carryin => counter_1_1_cry_13,
            carryout => counter_1_1_cry_14,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_15_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2594\,
            in2 => \_gnd_net_\,
            in3 => \N__2271\,
            lcout => \counter_1Z0Z_15\,
            ltout => OPEN,
            carryin => counter_1_1_cry_14,
            carryout => counter_1_1_cry_15,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_16_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2529\,
            in2 => \_gnd_net_\,
            in3 => \N__2268\,
            lcout => \counter_1Z0Z_16\,
            ltout => OPEN,
            carryin => counter_1_1_cry_15,
            carryout => counter_1_1_cry_16,
            clk => \N__4412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_17_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2543\,
            in2 => \_gnd_net_\,
            in3 => \N__2265\,
            lcout => \counter_1Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => counter_1_1_cry_17,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_18_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2568\,
            in2 => \_gnd_net_\,
            in3 => \N__2262\,
            lcout => \counter_1Z0Z_18\,
            ltout => OPEN,
            carryin => counter_1_1_cry_17,
            carryout => counter_1_1_cry_18,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_19_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2556\,
            in2 => \_gnd_net_\,
            in3 => \N__2259\,
            lcout => \counter_1Z0Z_19\,
            ltout => OPEN,
            carryin => counter_1_1_cry_18,
            carryout => counter_1_1_cry_19,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_20_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2517\,
            in2 => \_gnd_net_\,
            in3 => \N__2256\,
            lcout => \counter_1Z0Z_20\,
            ltout => OPEN,
            carryin => counter_1_1_cry_19,
            carryout => counter_1_1_cry_20,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_21_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2505\,
            in2 => \_gnd_net_\,
            in3 => \N__2253\,
            lcout => \counter_1Z0Z_21\,
            ltout => OPEN,
            carryin => counter_1_1_cry_20,
            carryout => counter_1_1_cry_21,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_22_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2478\,
            in2 => \_gnd_net_\,
            in3 => \N__2250\,
            lcout => \counter_1Z0Z_22\,
            ltout => OPEN,
            carryin => counter_1_1_cry_21,
            carryout => counter_1_1_cry_22,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_23_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2492\,
            in2 => \_gnd_net_\,
            in3 => \N__2247\,
            lcout => \counter_1Z0Z_23\,
            ltout => OPEN,
            carryin => counter_1_1_cry_22,
            carryout => counter_1_1_cry_23,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_24_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2454\,
            in2 => \_gnd_net_\,
            in3 => \N__2337\,
            lcout => \counter_1Z0Z_24\,
            ltout => OPEN,
            carryin => counter_1_1_cry_23,
            carryout => counter_1_1_cry_24,
            clk => \N__4409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_25_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2441\,
            in2 => \_gnd_net_\,
            in3 => \N__2334\,
            lcout => \counter_1Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => counter_1_1_cry_25,
            clk => \N__4408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_26_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2427\,
            in2 => \_gnd_net_\,
            in3 => \N__2331\,
            lcout => \counter_1Z0Z_26\,
            ltout => OPEN,
            carryin => counter_1_1_cry_25,
            carryout => counter_1_1_cry_26,
            clk => \N__4408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_27_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2466\,
            in2 => \_gnd_net_\,
            in3 => \N__2328\,
            lcout => \counter_1Z0Z_27\,
            ltout => OPEN,
            carryin => counter_1_1_cry_26,
            carryout => counter_1_1_cry_27,
            clk => \N__4408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_28_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2304\,
            in2 => \_gnd_net_\,
            in3 => \N__2325\,
            lcout => \counter_1Z0Z_28\,
            ltout => OPEN,
            carryin => counter_1_1_cry_27,
            carryout => counter_1_1_cry_28,
            clk => \N__4408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_29_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2313\,
            in2 => \_gnd_net_\,
            in3 => \N__2322\,
            lcout => \counter_1Z0Z_29\,
            ltout => OPEN,
            carryin => counter_1_1_cry_28,
            carryout => counter_1_1_cry_29,
            clk => \N__4408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_30_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2295\,
            in3 => \N__2319\,
            lcout => \counter_1Z0Z_30\,
            ltout => OPEN,
            carryin => counter_1_1_cry_29,
            carryout => counter_1_1_cry_30,
            clk => \N__4408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_31_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__2280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2316\,
            lcout => \counter_1Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_7_c_RNO_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2312\,
            in1 => \N__2303\,
            in2 => \N__2294\,
            in3 => \N__2279\,
            lcout => un4_counter_1_7_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_5_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__2997\,
            in1 => \N__3017\,
            in2 => \_gnd_net_\,
            in3 => \N__3709\,
            lcout => \counter_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4404\,
            ce => \N__3446\,
            sr => \_gnd_net_\
        );

    \un4_counter_2_0_c_RNO_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3013\,
            in1 => \N__2794\,
            in2 => \N__2985\,
            in3 => \N__2749\,
            lcout => un4_counter_2_0_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_1_c_RNO_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__2838\,
            in1 => \N__2953\,
            in2 => \N__2819\,
            in3 => \N__2926\,
            lcout => un4_counter_2_1_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_0_c_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2352\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => un4_counter_2_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_1_c_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2346\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_2_0,
            carryout => un4_counter_2_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_2_c_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2394\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_2_1,
            carryout => un4_counter_2_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_3_c_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2385\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_2_2,
            carryout => un4_counter_2_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_4_c_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2403\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_2_3,
            carryout => un4_counter_2_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_5_c_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_2_4,
            carryout => un4_counter_2_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_6_c_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2364\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_2_5,
            carryout => un4_counter_2_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_7_c_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2376\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_2_6,
            carryout => un4_counter_2_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_7_THRU_LUT4_0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2415\,
            lcout => \un4_counter_2_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_5_c_RNO_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3272\,
            in1 => \N__3032\,
            in2 => \N__3291\,
            in3 => \N__3257\,
            lcout => un4_counter_2_5_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_4_c_RNO_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3101\,
            in1 => \N__3086\,
            in2 => \N__3072\,
            in3 => \N__3051\,
            lcout => un4_counter_2_4_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_2_c_RNO_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2870\,
            in1 => \N__2900\,
            in2 => \N__2769\,
            in3 => \N__2885\,
            lcout => un4_counter_2_2_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_3_c_RNO_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3149\,
            in1 => \N__3116\,
            in2 => \N__3135\,
            in3 => \N__2855\,
            lcout => un4_counter_2_3_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_7_c_RNO_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3164\,
            in1 => \N__3179\,
            in2 => \N__3480\,
            in3 => \N__3458\,
            lcout => un4_counter_2_7_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_2_6_c_RNO_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3227\,
            in1 => \N__3194\,
            in2 => \N__3213\,
            in3 => \N__3242\,
            lcout => un4_counter_2_6_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_1_c_RNO_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2720\,
            in1 => \N__2708\,
            in2 => \N__2697\,
            in3 => \N__2681\,
            lcout => un4_counter_1_1_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_2_c_RNO_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2669\,
            in1 => \N__2657\,
            in2 => \N__2646\,
            in3 => \N__2630\,
            lcout => un4_counter_1_2_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_3_c_RNO_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2618\,
            in1 => \N__2606\,
            in2 => \N__2595\,
            in3 => \N__2579\,
            lcout => un4_counter_1_3_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_4_c_RNO_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2567\,
            in1 => \N__2555\,
            in2 => \N__2544\,
            in3 => \N__2528\,
            lcout => un4_counter_1_4_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_5_c_RNO_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2516\,
            in1 => \N__2504\,
            in2 => \N__2493\,
            in3 => \N__2477\,
            lcout => un4_counter_1_5_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_6_c_RNO_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2465\,
            in1 => \N__2453\,
            in2 => \N__2442\,
            in3 => \N__2426\,
            lcout => un4_counter_1_6_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_6_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__2984\,
            in1 => \N__2964\,
            in2 => \_gnd_net_\,
            in3 => \N__3706\,
            lcout => \counter_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => \N__3447\,
            sr => \_gnd_net_\
        );

    \counter_2_1_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2818\,
            in2 => \_gnd_net_\,
            in3 => \N__2841\,
            lcout => \counter_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => \N__3447\,
            sr => \_gnd_net_\
        );

    \counter_2_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__2778\,
            in1 => \N__3705\,
            in2 => \_gnd_net_\,
            in3 => \N__2796\,
            lcout => \counter_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => \N__3447\,
            sr => \_gnd_net_\
        );

    \counter_2_4_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__3704\,
            in1 => \_gnd_net_\,
            in2 => \N__2733\,
            in3 => \N__2751\,
            lcout => \counter_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => \N__3447\,
            sr => \_gnd_net_\
        );

    \counter_2_7_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__2937\,
            in1 => \N__2955\,
            in2 => \_gnd_net_\,
            in3 => \N__3707\,
            lcout => \counter_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => \N__3447\,
            sr => \_gnd_net_\
        );

    \counter_2_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2840\,
            lcout => \counter_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => \N__3447\,
            sr => \_gnd_net_\
        );

    \counter_2_8_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__2910\,
            in1 => \N__2928\,
            in2 => \_gnd_net_\,
            in3 => \N__3708\,
            lcout => \counter_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => \N__3447\,
            sr => \_gnd_net_\
        );

    \counter_2_1_cry_1_c_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2839\,
            in2 => \N__2820\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => counter_2_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_1_cry_1_THRU_LUT4_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2795\,
            in2 => \_gnd_net_\,
            in3 => \N__2772\,
            lcout => \counter_2_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => counter_2_1_cry_1,
            carryout => counter_2_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_3_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2768\,
            in2 => \_gnd_net_\,
            in3 => \N__2754\,
            lcout => \counter_2Z0Z_3\,
            ltout => OPEN,
            carryin => counter_2_1_cry_2,
            carryout => counter_2_1_cry_3,
            clk => \N__4402\,
            ce => \N__3445\,
            sr => \_gnd_net_\
        );

    \counter_2_1_cry_3_THRU_LUT4_0_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2750\,
            in2 => \_gnd_net_\,
            in3 => \N__2724\,
            lcout => \counter_2_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => counter_2_1_cry_3,
            carryout => counter_2_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_1_cry_4_THRU_LUT4_0_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3018\,
            in2 => \_gnd_net_\,
            in3 => \N__2988\,
            lcout => \counter_2_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => counter_2_1_cry_4,
            carryout => counter_2_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_1_cry_5_THRU_LUT4_0_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2983\,
            in2 => \_gnd_net_\,
            in3 => \N__2958\,
            lcout => \counter_2_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => counter_2_1_cry_5,
            carryout => counter_2_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_1_cry_6_THRU_LUT4_0_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2954\,
            in2 => \_gnd_net_\,
            in3 => \N__2931\,
            lcout => \counter_2_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => counter_2_1_cry_6,
            carryout => counter_2_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_1_cry_7_THRU_LUT4_0_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2927\,
            in2 => \_gnd_net_\,
            in3 => \N__2904\,
            lcout => \counter_2_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => counter_2_1_cry_7,
            carryout => counter_2_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_9_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2901\,
            in2 => \_gnd_net_\,
            in3 => \N__2889\,
            lcout => \counter_2Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => counter_2_1_cry_9,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_10_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2886\,
            in2 => \_gnd_net_\,
            in3 => \N__2874\,
            lcout => \counter_2Z0Z_10\,
            ltout => OPEN,
            carryin => counter_2_1_cry_9,
            carryout => counter_2_1_cry_10,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_11_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2871\,
            in2 => \_gnd_net_\,
            in3 => \N__2859\,
            lcout => \counter_2Z0Z_11\,
            ltout => OPEN,
            carryin => counter_2_1_cry_10,
            carryout => counter_2_1_cry_11,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_12_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2856\,
            in2 => \_gnd_net_\,
            in3 => \N__2844\,
            lcout => \counter_2Z0Z_12\,
            ltout => OPEN,
            carryin => counter_2_1_cry_11,
            carryout => counter_2_1_cry_12,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_13_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3150\,
            in2 => \_gnd_net_\,
            in3 => \N__3138\,
            lcout => \counter_2Z0Z_13\,
            ltout => OPEN,
            carryin => counter_2_1_cry_12,
            carryout => counter_2_1_cry_13,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_14_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3134\,
            in2 => \_gnd_net_\,
            in3 => \N__3120\,
            lcout => \counter_2Z0Z_14\,
            ltout => OPEN,
            carryin => counter_2_1_cry_13,
            carryout => counter_2_1_cry_14,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_15_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3117\,
            in2 => \_gnd_net_\,
            in3 => \N__3105\,
            lcout => \counter_2Z0Z_15\,
            ltout => OPEN,
            carryin => counter_2_1_cry_14,
            carryout => counter_2_1_cry_15,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_16_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3102\,
            in2 => \_gnd_net_\,
            in3 => \N__3090\,
            lcout => \counter_2Z0Z_16\,
            ltout => OPEN,
            carryin => counter_2_1_cry_15,
            carryout => counter_2_1_cry_16,
            clk => \N__4401\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \counter_2_17_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3087\,
            in2 => \_gnd_net_\,
            in3 => \N__3075\,
            lcout => \counter_2Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => counter_2_1_cry_17,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_18_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3068\,
            in2 => \_gnd_net_\,
            in3 => \N__3054\,
            lcout => \counter_2Z0Z_18\,
            ltout => OPEN,
            carryin => counter_2_1_cry_17,
            carryout => counter_2_1_cry_18,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_19_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3050\,
            in2 => \_gnd_net_\,
            in3 => \N__3036\,
            lcout => \counter_2Z0Z_19\,
            ltout => OPEN,
            carryin => counter_2_1_cry_18,
            carryout => counter_2_1_cry_19,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_20_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3033\,
            in2 => \_gnd_net_\,
            in3 => \N__3021\,
            lcout => \counter_2Z0Z_20\,
            ltout => OPEN,
            carryin => counter_2_1_cry_19,
            carryout => counter_2_1_cry_20,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_21_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3290\,
            in2 => \_gnd_net_\,
            in3 => \N__3276\,
            lcout => \counter_2Z0Z_21\,
            ltout => OPEN,
            carryin => counter_2_1_cry_20,
            carryout => counter_2_1_cry_21,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_22_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3273\,
            in2 => \_gnd_net_\,
            in3 => \N__3261\,
            lcout => \counter_2Z0Z_22\,
            ltout => OPEN,
            carryin => counter_2_1_cry_21,
            carryout => counter_2_1_cry_22,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_23_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3258\,
            in2 => \_gnd_net_\,
            in3 => \N__3246\,
            lcout => \counter_2Z0Z_23\,
            ltout => OPEN,
            carryin => counter_2_1_cry_22,
            carryout => counter_2_1_cry_23,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_24_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3243\,
            in2 => \_gnd_net_\,
            in3 => \N__3231\,
            lcout => \counter_2Z0Z_24\,
            ltout => OPEN,
            carryin => counter_2_1_cry_23,
            carryout => counter_2_1_cry_24,
            clk => \N__4403\,
            ce => \N__3442\,
            sr => \_gnd_net_\
        );

    \counter_2_25_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3228\,
            in2 => \_gnd_net_\,
            in3 => \N__3216\,
            lcout => \counter_2Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => counter_2_1_cry_25,
            clk => \N__4405\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \counter_2_26_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3212\,
            in2 => \_gnd_net_\,
            in3 => \N__3198\,
            lcout => \counter_2Z0Z_26\,
            ltout => OPEN,
            carryin => counter_2_1_cry_25,
            carryout => counter_2_1_cry_26,
            clk => \N__4405\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \counter_2_27_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3195\,
            in2 => \_gnd_net_\,
            in3 => \N__3183\,
            lcout => \counter_2Z0Z_27\,
            ltout => OPEN,
            carryin => counter_2_1_cry_26,
            carryout => counter_2_1_cry_27,
            clk => \N__4405\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \counter_2_28_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3180\,
            in2 => \_gnd_net_\,
            in3 => \N__3168\,
            lcout => \counter_2Z0Z_28\,
            ltout => OPEN,
            carryin => counter_2_1_cry_27,
            carryout => counter_2_1_cry_28,
            clk => \N__4405\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \counter_2_29_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3165\,
            in2 => \_gnd_net_\,
            in3 => \N__3153\,
            lcout => \counter_2Z0Z_29\,
            ltout => OPEN,
            carryin => counter_2_1_cry_28,
            carryout => counter_2_1_cry_29,
            clk => \N__4405\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \counter_2_30_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3479\,
            in2 => \_gnd_net_\,
            in3 => \N__3465\,
            lcout => \counter_2Z0Z_30\,
            ltout => OPEN,
            carryin => counter_2_1_cry_29,
            carryout => counter_2_1_cry_30,
            clk => \N__4405\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \counter_2_31_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3459\,
            in2 => \_gnd_net_\,
            in3 => \N__3462\,
            lcout => \counter_2Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4405\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \counter_1_3_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3651\,
            in1 => \N__3423\,
            in2 => \_gnd_net_\,
            in3 => \N__3368\,
            lcout => \counter_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_2_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3395\,
            in1 => \N__3652\,
            in2 => \_gnd_net_\,
            in3 => \N__3411\,
            lcout => \counter_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_0_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3653\,
            in2 => \_gnd_net_\,
            in3 => \N__3345\,
            lcout => \counter_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_0_c_RNO_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3391\,
            in1 => \N__3367\,
            in2 => \N__3350\,
            in3 => \N__3313\,
            lcout => un4_counter_1_0_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_1_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3654\,
            in2 => \N__3320\,
            in3 => \N__3346\,
            lcout => \counter_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_0_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3300\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => un4_counter_1_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_1_c_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3606\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_1_0,
            carryout => un4_counter_1_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_2_c_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_1_1,
            carryout => un4_counter_1_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_3_c_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3576\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_1_2,
            carryout => un4_counter_1_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_4_c_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3561\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_1_3,
            carryout => un4_counter_1_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_5_c_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3546\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_1_4,
            carryout => un4_counter_1_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_6_c_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3531\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_1_5,
            carryout => un4_counter_1_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_7_c_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3516\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_1_6,
            carryout => un4_counter_1_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_1_7_THRU_LUT4_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3501\,
            lcout => \un4_counter_1_7_THRU_CO\,
            ltout => \un4_counter_1_7_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_1MHz_RNINCP9_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3498\,
            in3 => \N__3731\,
            lcout => \clk_1Khz_cnv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_1MHz_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__3732\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3650\,
            lcout => \clk_1MHz_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_2Hz_RNO_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__3749\,
            in1 => \N__3734\,
            in2 => \_gnd_net_\,
            in3 => \N__3639\,
            lcout => \clk_2Hz_cnv_m3_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_1Khz_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001011110000"
        )
    port map (
            in0 => \N__3700\,
            in1 => \N__3735\,
            in2 => \N__3753\,
            in3 => \N__3640\,
            lcout => \clk_1Khz_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_2HzZ0_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__4491\,
            in1 => \N__3780\,
            in2 => \N__3770\,
            in3 => \N__3711\,
            lcout => \clk_2Hz_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_1Khz_RNIDQNN_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3748\,
            in1 => \N__3733\,
            in2 => \N__3710\,
            in3 => \N__3638\,
            lcout => \clk_1Khz_RNIDQNNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4029\,
            lcout => \counter_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4415\,
            ce => \N__4350\,
            sr => \_gnd_net_\
        );

    \counter_3_6_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4485\,
            in1 => \N__3900\,
            in2 => \_gnd_net_\,
            in3 => \N__3920\,
            lcout => \counter_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4418\,
            ce => \N__4348\,
            sr => \_gnd_net_\
        );

    \counter_3_5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3950\,
            in1 => \N__3930\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => \counter_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4418\,
            ce => \N__4348\,
            sr => \_gnd_net_\
        );

    \counter_3_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4486\,
            in1 => \N__4040\,
            in2 => \_gnd_net_\,
            in3 => \N__4061\,
            lcout => \counter_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4418\,
            ce => \N__4348\,
            sr => \_gnd_net_\
        );

    \un4_counter_3_3_c_RNO_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4112\,
            in1 => \N__4127\,
            in2 => \N__4098\,
            in3 => \N__4142\,
            lcout => un4_counter_3_3_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_1_c_RNO_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3916\,
            in1 => \N__4004\,
            in2 => \N__3891\,
            in3 => \N__4030\,
            lcout => un4_counter_3_1_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_2_c_RNO_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4179\,
            in1 => \N__4193\,
            in2 => \N__4161\,
            in3 => \N__3851\,
            lcout => un4_counter_3_2_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_0_c_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3813\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => un4_counter_3_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_1_c_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3798\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_3_0,
            carryout => un4_counter_3_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_2_c_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3792\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_3_1,
            carryout => un4_counter_3_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_3_c_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3786\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_3_2,
            carryout => un4_counter_3_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_4_c_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3819\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_3_3,
            carryout => un4_counter_3_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_5_c_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3825\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_3_4,
            carryout => un4_counter_3_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_6_c_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3807\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_3_5,
            carryout => un4_counter_3_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_7_c_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3834\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_counter_3_6,
            carryout => un4_counter_3_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_7_THRU_LUT4_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3837\,
            lcout => \un4_counter_3_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_7_c_RNO_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4532\,
            in1 => \N__4547\,
            in2 => \N__4515\,
            in3 => \N__4562\,
            lcout => un4_counter_3_7_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_5_c_RNO_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4241\,
            in1 => \N__4256\,
            in2 => \N__4227\,
            in3 => \N__4271\,
            lcout => un4_counter_3_5_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_4_c_RNO_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4076\,
            in1 => \N__4304\,
            in2 => \N__4290\,
            in3 => \N__4319\,
            lcout => un4_counter_3_4_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_0_c_RNO_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3982\,
            in1 => \N__4062\,
            in2 => \N__3954\,
            in3 => \N__4445\,
            lcout => un4_counter_3_0_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_counter_3_6_c_RNO_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4610\,
            in1 => \N__4577\,
            in2 => \N__4596\,
            in3 => \N__4208\,
            lcout => un4_counter_3_6_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_4_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3966\,
            in1 => \N__3986\,
            in2 => \_gnd_net_\,
            in3 => \N__4469\,
            lcout => \counter_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4417\,
            ce => \N__4347\,
            sr => \_gnd_net_\
        );

    \counter_3_7_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3886\,
            in1 => \N__3864\,
            in2 => \_gnd_net_\,
            in3 => \N__4470\,
            lcout => \counter_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4417\,
            ce => \N__4347\,
            sr => \_gnd_net_\
        );

    \counter_3_1_cry_1_c_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4060\,
            in2 => \N__4041\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => counter_3_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4005\,
            in2 => \_gnd_net_\,
            in3 => \N__3993\,
            lcout => \counter_3Z0Z_2\,
            ltout => OPEN,
            carryin => counter_3_1_cry_1,
            carryout => counter_3_1_cry_2,
            clk => \N__4419\,
            ce => \N__4344\,
            sr => \_gnd_net_\
        );

    \counter_3_1_cry_2_THRU_LUT4_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4446\,
            in2 => \_gnd_net_\,
            in3 => \N__3990\,
            lcout => \counter_3_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => counter_3_1_cry_2,
            carryout => counter_3_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_1_cry_3_THRU_LUT4_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3987\,
            in2 => \_gnd_net_\,
            in3 => \N__3957\,
            lcout => \counter_3_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => counter_3_1_cry_3,
            carryout => counter_3_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_1_cry_4_THRU_LUT4_0_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3949\,
            in2 => \_gnd_net_\,
            in3 => \N__3924\,
            lcout => \counter_3_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => counter_3_1_cry_4,
            carryout => counter_3_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_1_cry_5_THRU_LUT4_0_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3921\,
            in3 => \N__3894\,
            lcout => \counter_3_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => counter_3_1_cry_5,
            carryout => counter_3_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_1_cry_6_THRU_LUT4_0_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3890\,
            in2 => \_gnd_net_\,
            in3 => \N__3855\,
            lcout => \counter_3_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => counter_3_1_cry_6,
            carryout => counter_3_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_8_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3852\,
            in2 => \_gnd_net_\,
            in3 => \N__3840\,
            lcout => \counter_3Z0Z_8\,
            ltout => OPEN,
            carryin => counter_3_1_cry_7,
            carryout => counter_3_1_cry_8,
            clk => \N__4419\,
            ce => \N__4344\,
            sr => \_gnd_net_\
        );

    \counter_3_9_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4194\,
            in2 => \_gnd_net_\,
            in3 => \N__4182\,
            lcout => \counter_3Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => counter_3_1_cry_9,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_10_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4178\,
            in2 => \_gnd_net_\,
            in3 => \N__4164\,
            lcout => \counter_3Z0Z_10\,
            ltout => OPEN,
            carryin => counter_3_1_cry_9,
            carryout => counter_3_1_cry_10,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_11_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4160\,
            in2 => \_gnd_net_\,
            in3 => \N__4146\,
            lcout => \counter_3Z0Z_11\,
            ltout => OPEN,
            carryin => counter_3_1_cry_10,
            carryout => counter_3_1_cry_11,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_12_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4143\,
            in2 => \_gnd_net_\,
            in3 => \N__4131\,
            lcout => \counter_3Z0Z_12\,
            ltout => OPEN,
            carryin => counter_3_1_cry_11,
            carryout => counter_3_1_cry_12,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_13_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4128\,
            in2 => \_gnd_net_\,
            in3 => \N__4116\,
            lcout => \counter_3Z0Z_13\,
            ltout => OPEN,
            carryin => counter_3_1_cry_12,
            carryout => counter_3_1_cry_13,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_14_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4113\,
            in2 => \_gnd_net_\,
            in3 => \N__4101\,
            lcout => \counter_3Z0Z_14\,
            ltout => OPEN,
            carryin => counter_3_1_cry_13,
            carryout => counter_3_1_cry_14,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_15_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4094\,
            in2 => \_gnd_net_\,
            in3 => \N__4080\,
            lcout => \counter_3Z0Z_15\,
            ltout => OPEN,
            carryin => counter_3_1_cry_14,
            carryout => counter_3_1_cry_15,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_16_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4077\,
            in2 => \_gnd_net_\,
            in3 => \N__4065\,
            lcout => \counter_3Z0Z_16\,
            ltout => OPEN,
            carryin => counter_3_1_cry_15,
            carryout => counter_3_1_cry_16,
            clk => \N__4416\,
            ce => \N__4343\,
            sr => \_gnd_net_\
        );

    \counter_3_17_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4320\,
            in2 => \_gnd_net_\,
            in3 => \N__4308\,
            lcout => \counter_3Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => counter_3_1_cry_17,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_18_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4305\,
            in2 => \_gnd_net_\,
            in3 => \N__4293\,
            lcout => \counter_3Z0Z_18\,
            ltout => OPEN,
            carryin => counter_3_1_cry_17,
            carryout => counter_3_1_cry_18,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_19_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4289\,
            in2 => \_gnd_net_\,
            in3 => \N__4275\,
            lcout => \counter_3Z0Z_19\,
            ltout => OPEN,
            carryin => counter_3_1_cry_18,
            carryout => counter_3_1_cry_19,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_20_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4272\,
            in2 => \_gnd_net_\,
            in3 => \N__4260\,
            lcout => \counter_3Z0Z_20\,
            ltout => OPEN,
            carryin => counter_3_1_cry_19,
            carryout => counter_3_1_cry_20,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_21_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4257\,
            in2 => \_gnd_net_\,
            in3 => \N__4245\,
            lcout => \counter_3Z0Z_21\,
            ltout => OPEN,
            carryin => counter_3_1_cry_20,
            carryout => counter_3_1_cry_21,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_22_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4242\,
            in2 => \_gnd_net_\,
            in3 => \N__4230\,
            lcout => \counter_3Z0Z_22\,
            ltout => OPEN,
            carryin => counter_3_1_cry_21,
            carryout => counter_3_1_cry_22,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_23_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4226\,
            in2 => \_gnd_net_\,
            in3 => \N__4212\,
            lcout => \counter_3Z0Z_23\,
            ltout => OPEN,
            carryin => counter_3_1_cry_22,
            carryout => counter_3_1_cry_23,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_24_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4209\,
            in2 => \_gnd_net_\,
            in3 => \N__4197\,
            lcout => \counter_3Z0Z_24\,
            ltout => OPEN,
            carryin => counter_3_1_cry_23,
            carryout => counter_3_1_cry_24,
            clk => \N__4420\,
            ce => \N__4345\,
            sr => \_gnd_net_\
        );

    \counter_3_25_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4611\,
            in2 => \_gnd_net_\,
            in3 => \N__4599\,
            lcout => \counter_3Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => counter_3_1_cry_25,
            clk => \N__4421\,
            ce => \N__4346\,
            sr => \_gnd_net_\
        );

    \counter_3_26_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4595\,
            in2 => \_gnd_net_\,
            in3 => \N__4581\,
            lcout => \counter_3Z0Z_26\,
            ltout => OPEN,
            carryin => counter_3_1_cry_25,
            carryout => counter_3_1_cry_26,
            clk => \N__4421\,
            ce => \N__4346\,
            sr => \_gnd_net_\
        );

    \counter_3_27_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4578\,
            in2 => \_gnd_net_\,
            in3 => \N__4566\,
            lcout => \counter_3Z0Z_27\,
            ltout => OPEN,
            carryin => counter_3_1_cry_26,
            carryout => counter_3_1_cry_27,
            clk => \N__4421\,
            ce => \N__4346\,
            sr => \_gnd_net_\
        );

    \counter_3_28_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4563\,
            in2 => \_gnd_net_\,
            in3 => \N__4551\,
            lcout => \counter_3Z0Z_28\,
            ltout => OPEN,
            carryin => counter_3_1_cry_27,
            carryout => counter_3_1_cry_28,
            clk => \N__4421\,
            ce => \N__4346\,
            sr => \_gnd_net_\
        );

    \counter_3_29_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4548\,
            in2 => \_gnd_net_\,
            in3 => \N__4536\,
            lcout => \counter_3Z0Z_29\,
            ltout => OPEN,
            carryin => counter_3_1_cry_28,
            carryout => counter_3_1_cry_29,
            clk => \N__4421\,
            ce => \N__4346\,
            sr => \_gnd_net_\
        );

    \counter_3_30_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4533\,
            in2 => \_gnd_net_\,
            in3 => \N__4521\,
            lcout => \counter_3Z0Z_30\,
            ltout => OPEN,
            carryin => counter_3_1_cry_29,
            carryout => counter_3_1_cry_30,
            clk => \N__4421\,
            ce => \N__4346\,
            sr => \_gnd_net_\
        );

    \counter_3_31_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4514\,
            in2 => \_gnd_net_\,
            in3 => \N__4518\,
            lcout => \counter_3Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4421\,
            ce => \N__4346\,
            sr => \_gnd_net_\
        );

    \counter_3_3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4500\,
            in1 => \N__4441\,
            in2 => \_gnd_net_\,
            in3 => \N__4487\,
            lcout => \counter_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4422\,
            ce => \N__4349\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
