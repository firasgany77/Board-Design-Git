-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 14 2022 09:26:23

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : in std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \VCCG0\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal v33a_enn : std_logic;
signal v5s_enn : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \VPP_VDDQ.un1_curr_state12_0_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state11\ : std_logic;
signal \VPP_VDDQ.un1_vddq_pwrgdZ0_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_curr_state13_0\ : std_logic;
signal \VPP_VDDQ.un1_vddq_pwrgdZ0\ : std_logic;
signal slp_s4n : std_logic;
signal vccst_en : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \vccst_en_cascade_\ : std_logic;
signal vpp_en : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un6_count_8_cascade_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un6_count_9\ : std_logic;
signal \PCH_PWRGD.un4_count_11\ : std_logic;
signal \PCH_PWRGD.un4_count_10\ : std_logic;
signal \PCH_PWRGD.un4_count_8_cascade_\ : std_logic;
signal \PCH_PWRGD.un4_count_9\ : std_logic;
signal \PCH_PWRGD_un1_delayed_vccin_ok_0_sqmuxa_0_cascade_\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.N_3_i_cascade_\ : std_logic;
signal \VPP_VDDQ.N_15_0\ : std_logic;
signal \PCH_PWRGD.N_6_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_RNI0TJM7Z0Z_0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_1_sqmuxa\ : std_logic;
signal \VPP_VDDQ.un6_count\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_s_1_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_okZ0\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_stateZ1Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state12\ : std_logic;
signal \PCH_PWRGD.N_3_i\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.i3_mux_0_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal pch_pwrok : std_logic;
signal vccst_pwrgd : std_logic;
signal \PCH_PWRGD.un1_curr_state10_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_2\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.countZ0Z_10\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.N_15_2\ : std_logic;
signal \G_12\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_0\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \VPP_VDDQ.g0_3_a3_0_1_cascade_\ : std_logic;
signal \VPP_VDDQ.N_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_6_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_12\ : std_logic;
signal \VPP_VDDQ.count_2_1_11_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \VPP_VDDQ.count_2_1_6\ : std_logic;
signal \VPP_VDDQ.count_2_RNI25V3Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIZ0_cascade_\ : std_logic;
signal \VPP_VDDQ.m4_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_4\ : std_logic;
signal \VPP_VDDQ.count_2_1_4_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_en_0_tz_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_en_cascade_\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \VPP_VDDQ.un1_clk_100khz_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIRZ0Z9731\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVFZ0Z931\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\ : std_logic;
signal \VPP_VDDQ.count_2_1_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_1_12\ : std_logic;
signal \VPP_VDDQ.count_2_1_13_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.count_2_1_14_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_14\ : std_logic;
signal \VPP_VDDQ.count_2_0_2\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal v5a_ok : std_logic;
signal v33a_ok : std_logic;
signal slp_susn : std_logic;
signal v1p8a_ok : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \VPP_VDDQ.m4_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.m6_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_e_0Z0Z_1\ : std_logic;
signal \VPP_VDDQ.GZ0Z_76\ : std_logic;
signal \VPP_VDDQ.count_2_1_3_cascade_\ : std_logic;
signal vddq_ok : std_logic;
signal \clk_100Khz_signalkeep\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_RNOZ0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un5_clk_100khz_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_4_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_8_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.N_1_i_12\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_14_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_RNI_0Z0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.count_2_1_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_10_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_10\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state10_0\ : std_logic;
signal \RSMRST_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\ : std_logic;
signal \G_29\ : std_logic;
signal \G_29_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_15_1\ : std_logic;
signal slp_s3n : std_logic;
signal \RSMRST_PWRGD.curr_state10_cascade_\ : std_logic;
signal rsmrstn : std_logic;
signal \VPP_VDDQ.g0_0_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \VPP_VDDQ.count_2_en\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_1\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_7_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_8\ : std_logic;
signal \VPP_VDDQ.N_10\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_9_cascade_\ : std_logic;
signal \VPP_VDDQ.N_9\ : std_logic;
signal \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\ : std_logic;
signal \VPP_VDDQ.m4_1\ : std_logic;
signal \VPP_VDDQ.un5_clk_100khz\ : std_logic;
signal \VPP_VDDQ.count_2_1_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.un4_count_11\ : std_logic;
signal \RSMRST_PWRGD.un4_count_10\ : std_logic;
signal \RSMRST_PWRGD.un4_count_8_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un4_count_9\ : std_logic;
signal \RSMRST_PWRGD.i3_mux_0_cascade_\ : std_logic;
signal v33s_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal v5s_ok : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_1\ : std_logic;
signal vccin_en : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal \RSMRST_PWRGD.N_1_i\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.N_6_cascade_\ : std_logic;
signal \G_10\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal fpga_osc : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    \SUSWARN_N_wire\ <= SUSWARN_N;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9794\,
            DIN => \N__9793\,
            DOUT => \N__9792\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9794\,
            PADOUT => \N__9793\,
            PADIN => \N__9792\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9785\,
            DIN => \N__9784\,
            DOUT => \N__9783\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9785\,
            PADOUT => \N__9784\,
            PADIN => \N__9783\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4045\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9776\,
            DIN => \N__9775\,
            DOUT => \N__9774\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9776\,
            PADOUT => \N__9775\,
            PADIN => \N__9774\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__6297\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9767\,
            DIN => \N__9766\,
            DOUT => \N__9765\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9767\,
            PADOUT => \N__9766\,
            PADIN => \N__9765\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4054\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9758\,
            DIN => \N__9757\,
            DOUT => \N__9756\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9758\,
            PADOUT => \N__9757\,
            PADIN => \N__9756\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9749\,
            DIN => \N__9748\,
            DOUT => \N__9747\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9749\,
            PADOUT => \N__9748\,
            PADIN => \N__9747\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9740\,
            DIN => \N__9739\,
            DOUT => \N__9738\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9740\,
            PADOUT => \N__9739\,
            PADIN => \N__9738\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9731\,
            DIN => \N__9730\,
            DOUT => \N__9729\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9731\,
            PADOUT => \N__9730\,
            PADIN => \N__9729\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9722\,
            DIN => \N__9721\,
            DOUT => \N__9720\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9722\,
            PADOUT => \N__9721\,
            PADIN => \N__9720\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4036\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9713\,
            DIN => \N__9712\,
            DOUT => \N__9711\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9713\,
            PADOUT => \N__9712\,
            PADIN => \N__9711\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9704\,
            DIN => \N__9703\,
            DOUT => \N__9702\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9704\,
            PADOUT => \N__9703\,
            PADIN => \N__9702\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9695\,
            DIN => \N__9694\,
            DOUT => \N__9693\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9695\,
            PADOUT => \N__9694\,
            PADIN => \N__9693\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9686\,
            DIN => \N__9685\,
            DOUT => \N__9684\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9686\,
            PADOUT => \N__9685\,
            PADIN => \N__9684\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9677\,
            DIN => \N__9676\,
            DOUT => \N__9675\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9677\,
            PADOUT => \N__9676\,
            PADIN => \N__9675\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9668\,
            DIN => \N__9667\,
            DOUT => \N__9666\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9668\,
            PADOUT => \N__9667\,
            PADIN => \N__9666\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9659\,
            DIN => \N__9658\,
            DOUT => \N__9657\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9659\,
            PADOUT => \N__9658\,
            PADIN => \N__9657\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9650\,
            DIN => \N__9649\,
            DOUT => \N__9648\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9650\,
            PADOUT => \N__9649\,
            PADIN => \N__9648\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4267\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9641\,
            DIN => \N__9640\,
            DOUT => \N__9639\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9641\,
            PADOUT => \N__9640\,
            PADIN => \N__9639\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9632\,
            DIN => \N__9631\,
            DOUT => \N__9630\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9632\,
            PADOUT => \N__9631\,
            PADIN => \N__9630\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9623\,
            DIN => \N__9622\,
            DOUT => \N__9621\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9623\,
            PADOUT => \N__9622\,
            PADIN => \N__9621\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9614\,
            DIN => \N__9613\,
            DOUT => \N__9612\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9614\,
            PADOUT => \N__9613\,
            PADIN => \N__9612\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9605\,
            DIN => \N__9604\,
            DOUT => \N__9603\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9605\,
            PADOUT => \N__9604\,
            PADIN => \N__9603\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9596\,
            DIN => \N__9595\,
            DOUT => \N__9594\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9596\,
            PADOUT => \N__9595\,
            PADIN => \N__9594\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9587\,
            DIN => \N__9586\,
            DOUT => \N__9585\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9587\,
            PADOUT => \N__9586\,
            PADIN => \N__9585\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9578\,
            DIN => \N__9577\,
            DOUT => \N__9576\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9578\,
            PADOUT => \N__9577\,
            PADIN => \N__9576\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__7813\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9569\,
            DIN => \N__9568\,
            DOUT => \N__9567\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9569\,
            PADOUT => \N__9568\,
            PADIN => \N__9567\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9560\,
            DIN => \N__9559\,
            DOUT => \N__9558\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9560\,
            PADOUT => \N__9559\,
            PADIN => \N__9558\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4624\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9551\,
            DIN => \N__9550\,
            DOUT => \N__9549\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9551\,
            PADOUT => \N__9550\,
            PADIN => \N__9549\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4663\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9542\,
            DIN => \N__9541\,
            DOUT => \N__9540\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9542\,
            PADOUT => \N__9541\,
            PADIN => \N__9540\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9533\,
            DIN => \N__9532\,
            DOUT => \N__9531\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9533\,
            PADOUT => \N__9532\,
            PADIN => \N__9531\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9524\,
            DIN => \N__9523\,
            DOUT => \N__9522\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9524\,
            PADOUT => \N__9523\,
            PADIN => \N__9522\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9515\,
            DIN => \N__9514\,
            DOUT => \N__9513\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9515\,
            PADOUT => \N__9514\,
            PADIN => \N__9513\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9506\,
            DIN => \N__9505\,
            DOUT => \N__9504\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9506\,
            PADOUT => \N__9505\,
            PADIN => \N__9504\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__7234\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9497\,
            DIN => \N__9496\,
            DOUT => \N__9495\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9497\,
            PADOUT => \N__9496\,
            PADIN => \N__9495\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9488\,
            DIN => \N__9487\,
            DOUT => \N__9486\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9488\,
            PADOUT => \N__9487\,
            PADIN => \N__9486\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9479\,
            DIN => \N__9478\,
            DOUT => \N__9477\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9479\,
            PADOUT => \N__9478\,
            PADIN => \N__9477\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4231\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9470\,
            DIN => \N__9469\,
            DOUT => \N__9468\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9470\,
            PADOUT => \N__9469\,
            PADIN => \N__9468\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9461\,
            DIN => \N__9460\,
            DOUT => \N__9459\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9461\,
            PADOUT => \N__9460\,
            PADIN => \N__9459\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9452\,
            DIN => \N__9451\,
            DOUT => \N__9450\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9452\,
            PADOUT => \N__9451\,
            PADIN => \N__9450\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9443\,
            DIN => \N__9442\,
            DOUT => \N__9441\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9443\,
            PADOUT => \N__9442\,
            PADIN => \N__9441\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9434\,
            DIN => \N__9433\,
            DOUT => \N__9432\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9434\,
            PADOUT => \N__9433\,
            PADIN => \N__9432\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__6232\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9425\,
            DIN => \N__9424\,
            DOUT => \N__9423\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9425\,
            PADOUT => \N__9424\,
            PADIN => \N__9423\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9416\,
            DIN => \N__9415\,
            DOUT => \N__9414\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9416\,
            PADOUT => \N__9415\,
            PADIN => \N__9414\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4032\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9407\,
            DIN => \N__9406\,
            DOUT => \N__9405\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9407\,
            PADOUT => \N__9406\,
            PADIN => \N__9405\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9398\,
            DIN => \N__9397\,
            DOUT => \N__9396\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9398\,
            PADOUT => \N__9397\,
            PADIN => \N__9396\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__7219\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9389\,
            DIN => \N__9388\,
            DOUT => \N__9387\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9389\,
            PADOUT => \N__9388\,
            PADIN => \N__9387\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__6301\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9380\,
            DIN => \N__9379\,
            DOUT => \N__9378\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9380\,
            PADOUT => \N__9379\,
            PADIN => \N__9378\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9371\,
            DIN => \N__9370\,
            DOUT => \N__9369\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9371\,
            PADOUT => \N__9370\,
            PADIN => \N__9369\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9362\,
            DIN => \N__9361\,
            DOUT => \N__9360\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9362\,
            PADOUT => \N__9361\,
            PADIN => \N__9360\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9353\,
            DIN => \N__9352\,
            DOUT => \N__9351\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9353\,
            PADOUT => \N__9352\,
            PADIN => \N__9351\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__7233\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9344\,
            DIN => \N__9343\,
            DOUT => \N__9342\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9344\,
            PADOUT => \N__9343\,
            PADIN => \N__9342\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__9202\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9335\,
            DIN => \N__9334\,
            DOUT => \N__9333\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9335\,
            PADOUT => \N__9334\,
            PADIN => \N__9333\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9326\,
            DIN => \N__9325\,
            DOUT => \N__9324\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9326\,
            PADOUT => \N__9325\,
            PADIN => \N__9324\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9317\,
            DIN => \N__9316\,
            DOUT => \N__9315\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9317\,
            PADOUT => \N__9316\,
            PADIN => \N__9315\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9308\,
            DIN => \N__9307\,
            DOUT => \N__9306\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9308\,
            PADOUT => \N__9307\,
            PADIN => \N__9306\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9299\,
            DIN => \N__9298\,
            DOUT => \N__9297\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9299\,
            PADOUT => \N__9298\,
            PADIN => \N__9297\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9290\,
            DIN => \N__9289\,
            DOUT => \N__9288\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9290\,
            PADOUT => \N__9289\,
            PADIN => \N__9288\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9281\,
            DIN => \N__9280\,
            DOUT => \N__9279\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9281\,
            PADOUT => \N__9280\,
            PADIN => \N__9279\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4662\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9272\,
            DIN => \N__9271\,
            DOUT => \N__9270\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9272\,
            PADOUT => \N__9271\,
            PADIN => \N__9270\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__2092\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9250\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9250\,
            I => \N__9247\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__9247\,
            I => \N__9244\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__9244\,
            I => v33s_ok
        );

    \I__2088\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9238\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__2086\ : Span4Mux_v
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__9229\,
            I => vccst_cpu_ok
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9220\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9220\,
            I => \N__9217\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__2079\ : Span4Mux_v
    port map (
            O => \N__9214\,
            I => \N__9211\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__9211\,
            I => v5s_ok
        );

    \I__2077\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9205\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9205\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_1\
        );

    \I__2075\ : IoInMux
    port map (
            O => \N__9202\,
            I => \N__9199\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9199\,
            I => \N__9196\
        );

    \I__2073\ : Span4Mux_s1_v
    port map (
            O => \N__9196\,
            I => \N__9193\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__9190\,
            I => vccin_en
        );

    \I__2070\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9177\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9186\,
            I => \N__9177\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9172\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9172\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9167\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9167\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9177\,
            I => \N__9164\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9172\,
            I => \N__9159\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9167\,
            I => \N__9159\
        );

    \I__2061\ : Odrv12
    port map (
            O => \N__9164\,
            I => rsmrst_pwrgd_signal
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__9159\,
            I => rsmrst_pwrgd_signal
        );

    \I__2059\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9147\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9147\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9144\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9147\,
            I => \N__9139\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9144\,
            I => \N__9139\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__9139\,
            I => \RSMRST_PWRGD.N_1_i\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9126\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9126\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9123\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9133\,
            I => \N__9116\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9116\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9116\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9126\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9123\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9116\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__9109\,
            I => \RSMRST_PWRGD.N_6_cascade_\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9085\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9085\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9085\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9085\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__9102\,
            I => \N__9081\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9056\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9056\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9056\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9056\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9029\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9029\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9029\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9029\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9026\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9019\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9019\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9019\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9079\,
            I => \N__9010\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9010\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9010\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9010\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9003\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9003\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9003\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9072\,
            I => \N__8994\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9071\,
            I => \N__8994\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9070\,
            I => \N__8994\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9069\,
            I => \N__8994\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9068\,
            I => \N__8985\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9067\,
            I => \N__8985\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9066\,
            I => \N__8985\
        );

    \I__2012\ : InMux
    port map (
            O => \N__9065\,
            I => \N__8985\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9056\,
            I => \N__8976\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9055\,
            I => \N__8967\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9054\,
            I => \N__8967\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9053\,
            I => \N__8967\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9052\,
            I => \N__8967\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9051\,
            I => \N__8958\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9050\,
            I => \N__8958\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9049\,
            I => \N__8958\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9048\,
            I => \N__8958\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9047\,
            I => \N__8951\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9046\,
            I => \N__8951\
        );

    \I__2000\ : InMux
    port map (
            O => \N__9045\,
            I => \N__8951\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9044\,
            I => \N__8944\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9043\,
            I => \N__8944\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9042\,
            I => \N__8944\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9041\,
            I => \N__8935\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9040\,
            I => \N__8935\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9039\,
            I => \N__8935\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9038\,
            I => \N__8935\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9029\,
            I => \N__8932\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9026\,
            I => \N__8927\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9019\,
            I => \N__8927\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__8922\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9003\,
            I => \N__8922\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__8994\,
            I => \N__8917\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8917\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8908\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8908\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8908\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8908\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8896\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8896\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__8976\,
            I => \N__8893\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8967\,
            I => \N__8890\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__8958\,
            I => \N__8885\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__8951\,
            I => \N__8885\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8944\,
            I => \N__8882\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8935\,
            I => \N__8873\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__8932\,
            I => \N__8873\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__8927\,
            I => \N__8873\
        );

    \I__1971\ : Span4Mux_h
    port map (
            O => \N__8922\,
            I => \N__8873\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__8917\,
            I => \N__8868\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8868\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8861\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8906\,
            I => \N__8861\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8861\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8852\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8852\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8852\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8852\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8896\,
            I => \N__8849\
        );

    \I__1960\ : Span4Mux_s1_h
    port map (
            O => \N__8893\,
            I => \N__8844\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__8890\,
            I => \N__8844\
        );

    \I__1958\ : Span4Mux_s2_h
    port map (
            O => \N__8885\,
            I => \N__8841\
        );

    \I__1957\ : Span4Mux_h
    port map (
            O => \N__8882\,
            I => \N__8836\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__8873\,
            I => \N__8836\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__8868\,
            I => \N__8833\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8861\,
            I => \N__8828\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8852\,
            I => \N__8828\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__8849\,
            I => \G_10\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__8844\,
            I => \G_10\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__8841\,
            I => \G_10\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__8836\,
            I => \G_10\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__8833\,
            I => \G_10\
        );

    \I__1947\ : Odrv12
    port map (
            O => \N__8828\,
            I => \G_10\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__8815\,
            I => \N__8808\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8800\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8800\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8800\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8811\,
            I => \N__8793\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8808\,
            I => \N__8793\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8793\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8800\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8793\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__1937\ : ClkMux
    port map (
            O => \N__8788\,
            I => \N__8784\
        );

    \I__1936\ : ClkMux
    port map (
            O => \N__8787\,
            I => \N__8781\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8784\,
            I => \N__8770\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8781\,
            I => \N__8767\
        );

    \I__1933\ : ClkMux
    port map (
            O => \N__8780\,
            I => \N__8764\
        );

    \I__1932\ : ClkMux
    port map (
            O => \N__8779\,
            I => \N__8760\
        );

    \I__1931\ : ClkMux
    port map (
            O => \N__8778\,
            I => \N__8755\
        );

    \I__1930\ : ClkMux
    port map (
            O => \N__8777\,
            I => \N__8749\
        );

    \I__1929\ : ClkMux
    port map (
            O => \N__8776\,
            I => \N__8744\
        );

    \I__1928\ : ClkMux
    port map (
            O => \N__8775\,
            I => \N__8741\
        );

    \I__1927\ : ClkMux
    port map (
            O => \N__8774\,
            I => \N__8738\
        );

    \I__1926\ : ClkMux
    port map (
            O => \N__8773\,
            I => \N__8734\
        );

    \I__1925\ : Span4Mux_s1_h
    port map (
            O => \N__8770\,
            I => \N__8726\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__8767\,
            I => \N__8726\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8764\,
            I => \N__8726\
        );

    \I__1922\ : ClkMux
    port map (
            O => \N__8763\,
            I => \N__8723\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8760\,
            I => \N__8720\
        );

    \I__1920\ : ClkMux
    port map (
            O => \N__8759\,
            I => \N__8717\
        );

    \I__1919\ : ClkMux
    port map (
            O => \N__8758\,
            I => \N__8714\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8755\,
            I => \N__8711\
        );

    \I__1917\ : ClkMux
    port map (
            O => \N__8754\,
            I => \N__8708\
        );

    \I__1916\ : ClkMux
    port map (
            O => \N__8753\,
            I => \N__8705\
        );

    \I__1915\ : ClkMux
    port map (
            O => \N__8752\,
            I => \N__8702\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8749\,
            I => \N__8699\
        );

    \I__1913\ : ClkMux
    port map (
            O => \N__8748\,
            I => \N__8696\
        );

    \I__1912\ : ClkMux
    port map (
            O => \N__8747\,
            I => \N__8693\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8690\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8741\,
            I => \N__8687\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8684\
        );

    \I__1908\ : ClkMux
    port map (
            O => \N__8737\,
            I => \N__8673\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8734\,
            I => \N__8670\
        );

    \I__1906\ : ClkMux
    port map (
            O => \N__8733\,
            I => \N__8667\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__8726\,
            I => \N__8662\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8723\,
            I => \N__8662\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__8720\,
            I => \N__8654\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8654\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8654\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__8711\,
            I => \N__8651\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8708\,
            I => \N__8648\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8705\,
            I => \N__8645\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8702\,
            I => \N__8642\
        );

    \I__1896\ : Span4Mux_h
    port map (
            O => \N__8699\,
            I => \N__8639\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8636\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8693\,
            I => \N__8633\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__8690\,
            I => \N__8626\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__8687\,
            I => \N__8626\
        );

    \I__1891\ : Span4Mux_h
    port map (
            O => \N__8684\,
            I => \N__8626\
        );

    \I__1890\ : ClkMux
    port map (
            O => \N__8683\,
            I => \N__8623\
        );

    \I__1889\ : ClkMux
    port map (
            O => \N__8682\,
            I => \N__8620\
        );

    \I__1888\ : ClkMux
    port map (
            O => \N__8681\,
            I => \N__8616\
        );

    \I__1887\ : ClkMux
    port map (
            O => \N__8680\,
            I => \N__8613\
        );

    \I__1886\ : ClkMux
    port map (
            O => \N__8679\,
            I => \N__8610\
        );

    \I__1885\ : ClkMux
    port map (
            O => \N__8678\,
            I => \N__8607\
        );

    \I__1884\ : ClkMux
    port map (
            O => \N__8677\,
            I => \N__8604\
        );

    \I__1883\ : ClkMux
    port map (
            O => \N__8676\,
            I => \N__8601\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__8673\,
            I => \N__8598\
        );

    \I__1881\ : Span4Mux_h
    port map (
            O => \N__8670\,
            I => \N__8591\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8591\
        );

    \I__1879\ : Span4Mux_h
    port map (
            O => \N__8662\,
            I => \N__8591\
        );

    \I__1878\ : ClkMux
    port map (
            O => \N__8661\,
            I => \N__8588\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__8654\,
            I => \N__8585\
        );

    \I__1876\ : Span4Mux_v
    port map (
            O => \N__8651\,
            I => \N__8576\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__8648\,
            I => \N__8576\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__8645\,
            I => \N__8576\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__8642\,
            I => \N__8576\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__8639\,
            I => \N__8563\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__8636\,
            I => \N__8563\
        );

    \I__1870\ : Span4Mux_h
    port map (
            O => \N__8633\,
            I => \N__8563\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__8626\,
            I => \N__8563\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8623\,
            I => \N__8563\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8620\,
            I => \N__8563\
        );

    \I__1866\ : ClkMux
    port map (
            O => \N__8619\,
            I => \N__8560\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8616\,
            I => \N__8551\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8613\,
            I => \N__8551\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8551\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8607\,
            I => \N__8551\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8546\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8601\,
            I => \N__8546\
        );

    \I__1859\ : Span4Mux_h
    port map (
            O => \N__8598\,
            I => \N__8539\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__8591\,
            I => \N__8539\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8588\,
            I => \N__8539\
        );

    \I__1856\ : Span4Mux_h
    port map (
            O => \N__8585\,
            I => \N__8533\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__8576\,
            I => \N__8533\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__8563\,
            I => \N__8530\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8560\,
            I => \N__8527\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__8551\,
            I => \N__8522\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__8546\,
            I => \N__8522\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__8539\,
            I => \N__8519\
        );

    \I__1849\ : ClkMux
    port map (
            O => \N__8538\,
            I => \N__8516\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__8533\,
            I => \N__8513\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__8530\,
            I => \N__8510\
        );

    \I__1846\ : Span12Mux_s5_h
    port map (
            O => \N__8527\,
            I => \N__8501\
        );

    \I__1845\ : Sp12to4
    port map (
            O => \N__8522\,
            I => \N__8501\
        );

    \I__1844\ : Sp12to4
    port map (
            O => \N__8519\,
            I => \N__8501\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8516\,
            I => \N__8501\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__8513\,
            I => fpga_osc
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__8510\,
            I => fpga_osc
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__8501\,
            I => fpga_osc
        );

    \I__1839\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8491\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8491\,
            I => \N__8485\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8482\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8479\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8488\,
            I => \N__8475\
        );

    \I__1834\ : Span4Mux_s3_v
    port map (
            O => \N__8485\,
            I => \N__8472\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8482\,
            I => \N__8469\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8479\,
            I => \N__8466\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8463\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8475\,
            I => \N__8460\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__8472\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__1828\ : Odrv12
    port map (
            O => \N__8469\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__1827\ : Odrv12
    port map (
            O => \N__8466\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8463\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__8460\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__8449\,
            I => \N__8445\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8442\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8439\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8442\,
            I => \N__8436\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8439\,
            I => \N__8433\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__8436\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__8433\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__8428\,
            I => \N__8425\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8406\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8402\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8395\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8395\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8395\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8387\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8381\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8378\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8365\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8365\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8365\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8365\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8365\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8365\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8360\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8360\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__8409\,
            I => \N__8355\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8406\,
            I => \N__8350\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8347\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8402\,
            I => \N__8342\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8395\,
            I => \N__8342\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__8394\,
            I => \N__8337\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8326\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8392\,
            I => \N__8326\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8326\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8326\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8387\,
            I => \N__8323\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8316\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8316\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8316\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8381\,
            I => \N__8307\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8307\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8307\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8360\,
            I => \N__8307\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8300\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8300\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8300\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8295\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8295\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__8350\,
            I => \N__8290\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8290\
        );

    \I__1775\ : Span4Mux_s3_v
    port map (
            O => \N__8342\,
            I => \N__8287\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8282\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8282\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8277\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8277\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8274\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8269\
        );

    \I__1768\ : Span4Mux_s2_v
    port map (
            O => \N__8323\,
            I => \N__8269\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8316\,
            I => \N__8262\
        );

    \I__1766\ : Span4Mux_s2_v
    port map (
            O => \N__8307\,
            I => \N__8262\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8262\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8295\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__8290\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__8287\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8282\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8277\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8274\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__8269\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__8262\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__8245\,
            I => \N__8219\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8214\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__8243\,
            I => \N__8211\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__8242\,
            I => \N__8208\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8202\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8193\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8193\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8193\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8184\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8184\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8184\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8184\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8233\,
            I => \N__8171\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8232\,
            I => \N__8171\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8171\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8171\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8171\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8171\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8168\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8165\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8162\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8159\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8156\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8153\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8145\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8145\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8145\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8214\,
            I => \N__8142\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8137\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8208\,
            I => \N__8137\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8130\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8130\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8130\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8127\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8122\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8122\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8193\,
            I => \N__8111\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8184\,
            I => \N__8111\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8171\,
            I => \N__8111\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8168\,
            I => \N__8111\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8165\,
            I => \N__8111\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8162\,
            I => \N__8105\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8159\,
            I => \N__8098\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8156\,
            I => \N__8098\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8153\,
            I => \N__8098\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8095\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8086\
        );

    \I__1709\ : Span12Mux_s8_h
    port map (
            O => \N__8142\,
            I => \N__8086\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8137\,
            I => \N__8086\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__8130\,
            I => \N__8086\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__8127\,
            I => \N__8079\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8122\,
            I => \N__8079\
        );

    \I__1704\ : Span4Mux_s3_v
    port map (
            O => \N__8111\,
            I => \N__8079\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8072\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8072\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8072\
        );

    \I__1700\ : Span4Mux_s2_h
    port map (
            O => \N__8105\,
            I => \N__8069\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__8098\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8095\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__8086\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__1696\ : Odrv4
    port map (
            O => \N__8079\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8072\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__8069\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__8050\,
            I => \N__8047\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__8047\,
            I => \VPP_VDDQ.count_2_1_2\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8040\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8037\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8040\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8037\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8028\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8025\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8028\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8025\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__8020\,
            I => \N__8016\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8019\,
            I => \N__8013\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8016\,
            I => \N__8010\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8013\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8010\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8005\,
            I => \N__8001\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7998\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8001\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7998\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7993\,
            I => \N__7989\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7986\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__7989\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__7986\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7977\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7974\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7977\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7974\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__7969\,
            I => \N__7965\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7962\
        );

    \I__1662\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7959\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7962\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7959\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7950\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7947\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__7950\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__7947\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7938\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7938\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7935\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7930\,
            I => \N__7926\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7923\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7926\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7923\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__7918\,
            I => \N__7914\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7911\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7908\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7911\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7908\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7899\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7896\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7899\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7896\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1638\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7887\
        );

    \I__1637\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7884\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7887\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__7884\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7875\
        );

    \I__1633\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7872\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7875\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7872\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__7867\,
            I => \N__7863\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7860\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7863\,
            I => \N__7857\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7860\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7857\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7848\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7845\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7848\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7845\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7837\,
            I => \RSMRST_PWRGD.un4_count_11\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7831\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7831\,
            I => \RSMRST_PWRGD.un4_count_10\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__7828\,
            I => \RSMRST_PWRGD.un4_count_8_cascade_\
        );

    \I__1616\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7822\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7822\,
            I => \RSMRST_PWRGD.un4_count_9\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \RSMRST_PWRGD.i3_mux_0_cascade_\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__7816\,
            I => \RSMRST_PWRGD.curr_state10_cascade_\
        );

    \I__1612\ : IoInMux
    port map (
            O => \N__7813\,
            I => \N__7810\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7810\,
            I => \N__7806\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7802\
        );

    \I__1609\ : IoSpan4Mux
    port map (
            O => \N__7806\,
            I => \N__7797\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7794\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7802\,
            I => \N__7790\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7787\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7784\
        );

    \I__1604\ : Span4Mux_s1_v
    port map (
            O => \N__7797\,
            I => \N__7779\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7779\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7776\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__7790\,
            I => \N__7769\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7787\,
            I => \N__7769\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__7784\,
            I => \N__7769\
        );

    \I__1598\ : Span4Mux_v
    port map (
            O => \N__7779\,
            I => \N__7762\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7776\,
            I => \N__7762\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__7769\,
            I => \N__7759\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7754\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7754\
        );

    \I__1593\ : Span4Mux_h
    port map (
            O => \N__7762\,
            I => \N__7751\
        );

    \I__1592\ : Span4Mux_h
    port map (
            O => \N__7759\,
            I => \N__7748\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7754\,
            I => rsmrstn
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__7751\,
            I => rsmrstn
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__7748\,
            I => rsmrstn
        );

    \I__1588\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7738\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7738\,
            I => \N__7735\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__7735\,
            I => \VPP_VDDQ.g0_0_0\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__7732\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__7729\,
            I => \N__7726\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7723\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7723\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__1581\ : CEMux
    port map (
            O => \N__7720\,
            I => \N__7714\
        );

    \I__1580\ : CEMux
    port map (
            O => \N__7719\,
            I => \N__7711\
        );

    \I__1579\ : CEMux
    port map (
            O => \N__7718\,
            I => \N__7694\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7691\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7714\,
            I => \N__7688\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7685\
        );

    \I__1575\ : CEMux
    port map (
            O => \N__7710\,
            I => \N__7674\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7674\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7674\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7671\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7666\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7705\,
            I => \N__7666\
        );

    \I__1569\ : CEMux
    port map (
            O => \N__7704\,
            I => \N__7663\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7660\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7653\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7653\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7700\,
            I => \N__7653\
        );

    \I__1564\ : CEMux
    port map (
            O => \N__7699\,
            I => \N__7646\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7646\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7646\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7694\,
            I => \N__7641\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7691\,
            I => \N__7641\
        );

    \I__1559\ : Span4Mux_s2_v
    port map (
            O => \N__7688\,
            I => \N__7636\
        );

    \I__1558\ : Span4Mux_s3_v
    port map (
            O => \N__7685\,
            I => \N__7633\
        );

    \I__1557\ : CEMux
    port map (
            O => \N__7684\,
            I => \N__7628\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7628\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7625\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7622\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7674\,
            I => \N__7615\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7615\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7666\,
            I => \N__7615\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7663\,
            I => \N__7604\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7660\,
            I => \N__7604\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7653\,
            I => \N__7604\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7604\
        );

    \I__1546\ : Span4Mux_s3_h
    port map (
            O => \N__7641\,
            I => \N__7604\
        );

    \I__1545\ : CEMux
    port map (
            O => \N__7640\,
            I => \N__7599\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7599\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__7636\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__7633\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7628\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7625\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7622\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__7615\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__7604\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7599\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7576\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7573\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__7580\,
            I => \N__7570\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7566\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7576\,
            I => \N__7563\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7573\,
            I => \N__7560\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7557\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7554\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7566\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__1526\ : Odrv12
    port map (
            O => \N__7563\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__7560\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7557\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7554\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7540\,
            I => \N__7535\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__7539\,
            I => \N__7532\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__7538\,
            I => \N__7528\
        );

    \I__1518\ : Span4Mux_v
    port map (
            O => \N__7535\,
            I => \N__7525\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7522\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7519\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7516\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__7525\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7522\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7519\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7516\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__7507\,
            I => \N__7502\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7499\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7495\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7502\,
            I => \N__7492\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7499\,
            I => \N__7488\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7498\,
            I => \N__7485\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7495\,
            I => \N__7482\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7492\,
            I => \N__7479\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7491\,
            I => \N__7476\
        );

    \I__1501\ : Span4Mux_h
    port map (
            O => \N__7488\,
            I => \N__7469\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7469\
        );

    \I__1499\ : Span4Mux_h
    port map (
            O => \N__7482\,
            I => \N__7469\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__7479\,
            I => \N__7466\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7476\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__7469\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__7466\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__7459\,
            I => \N__7456\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7453\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7453\,
            I => \N__7446\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7443\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7440\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__7450\,
            I => \N__7437\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7434\
        );

    \I__1487\ : Span4Mux_s3_h
    port map (
            O => \N__7446\,
            I => \N__7427\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7443\,
            I => \N__7427\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7440\,
            I => \N__7427\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7424\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7434\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__7427\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7424\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7413\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7410\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7413\,
            I => \N__7405\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7410\,
            I => \N__7402\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__7409\,
            I => \N__7399\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__7408\,
            I => \N__7395\
        );

    \I__1474\ : Span4Mux_h
    port map (
            O => \N__7405\,
            I => \N__7392\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__7402\,
            I => \N__7389\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7386\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7398\,
            I => \N__7383\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7380\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__7392\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__7389\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7386\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7383\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7380\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7366\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7366\,
            I => \N__7362\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__7365\,
            I => \N__7357\
        );

    \I__1461\ : Span4Mux_v
    port map (
            O => \N__7362\,
            I => \N__7354\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7361\,
            I => \N__7351\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7348\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7345\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__7354\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7351\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7348\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7345\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7333\,
            I => \VPP_VDDQ.g0_2_a2_1\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__7330\,
            I => \VPP_VDDQ.g0_2_a2_7_cascade_\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7323\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7317\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7314\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7311\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7308\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7305\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7302\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__7314\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7311\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7308\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7305\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__7302\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7288\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7288\,
            I => \N__7285\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__7285\,
            I => \N__7282\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__7282\,
            I => \VPP_VDDQ.g0_2_a2_8\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7276\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7273\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__7273\,
            I => \N__7270\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__7270\,
            I => \VPP_VDDQ.N_10\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__7267\,
            I => \VPP_VDDQ.g0_2_a2_9_cascade_\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7261\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7261\,
            I => \N__7258\
        );

    \I__1427\ : Odrv12
    port map (
            O => \N__7258\,
            I => \VPP_VDDQ.N_9\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7249\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7249\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__1423\ : Span4Mux_h
    port map (
            O => \N__7246\,
            I => \N__7243\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__7243\,
            I => \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7240\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7237\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__1419\ : IoInMux
    port map (
            O => \N__7234\,
            I => \N__7230\
        );

    \I__1418\ : IoInMux
    port map (
            O => \N__7233\,
            I => \N__7227\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__7230\,
            I => \N__7224\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7227\,
            I => \N__7221\
        );

    \I__1415\ : IoSpan4Mux
    port map (
            O => \N__7224\,
            I => \N__7214\
        );

    \I__1414\ : IoSpan4Mux
    port map (
            O => \N__7221\,
            I => \N__7214\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7211\
        );

    \I__1412\ : IoInMux
    port map (
            O => \N__7219\,
            I => \N__7208\
        );

    \I__1411\ : Span4Mux_s0_h
    port map (
            O => \N__7214\,
            I => \N__7202\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7202\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7199\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7196\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__7202\,
            I => \N__7192\
        );

    \I__1406\ : Span4Mux_s1_h
    port map (
            O => \N__7199\,
            I => \N__7187\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7196\,
            I => \N__7187\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7195\,
            I => \N__7184\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__7192\,
            I => \N__7181\
        );

    \I__1402\ : Span4Mux_h
    port map (
            O => \N__7187\,
            I => \N__7176\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7184\,
            I => \N__7176\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__7181\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__7176\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7171\,
            I => \bfn_11_10_0_\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__7168\,
            I => \N__7164\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7161\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7158\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7161\,
            I => \N__7155\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7158\,
            I => \N__7152\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__7155\,
            I => \RSMRST_PWRGD.un1_curr_state10_0\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__7152\,
            I => \RSMRST_PWRGD.un1_curr_state10_0\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \RSMRST_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\
        );

    \I__1389\ : SRMux
    port map (
            O => \N__7144\,
            I => \N__7140\
        );

    \I__1388\ : SRMux
    port map (
            O => \N__7143\,
            I => \N__7136\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7140\,
            I => \N__7133\
        );

    \I__1386\ : SRMux
    port map (
            O => \N__7139\,
            I => \N__7130\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7136\,
            I => \N__7127\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__7133\,
            I => \N__7122\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7130\,
            I => \N__7122\
        );

    \I__1382\ : Span4Mux_h
    port map (
            O => \N__7127\,
            I => \N__7119\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__7122\,
            I => \G_29\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__7119\,
            I => \G_29\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__7114\,
            I => \G_29_cascade_\
        );

    \I__1378\ : CEMux
    port map (
            O => \N__7111\,
            I => \N__7108\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7108\,
            I => \RSMRST_PWRGD.N_15_1\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7105\,
            I => \N__7102\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7102\,
            I => \N__7097\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7094\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7091\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__7097\,
            I => \N__7088\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7083\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7091\,
            I => \N__7083\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__7088\,
            I => \N__7078\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__7083\,
            I => \N__7078\
        );

    \I__1367\ : Sp12to4
    port map (
            O => \N__7078\,
            I => \N__7074\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7077\,
            I => \N__7071\
        );

    \I__1365\ : Span12Mux_s10_h
    port map (
            O => \N__7074\,
            I => \N__7066\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7071\,
            I => \N__7066\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__7066\,
            I => slp_s3n
        );

    \I__1362\ : InMux
    port map (
            O => \N__7063\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7060\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7057\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7054\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7051\,
            I => \bfn_11_9_0_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7048\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7045\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7042\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7039\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7032\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7035\,
            I => \N__7029\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7032\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_THRU_CO\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7029\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_THRU_CO\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7021\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__7018\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__7015\,
            I => \VPP_VDDQ.count_2_1_9_cascade_\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__7012\,
            I => \VPP_VDDQ.count_2_1_10_cascade_\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7009\,
            I => \N__7003\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7008\,
            I => \N__7003\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7003\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_THRU_CO\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__7000\,
            I => \VPP_VDDQ.count_2Z0Z_10_cascade_\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6994\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6994\,
            I => \VPP_VDDQ.count_2_0_10\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6991\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6988\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6985\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6975\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6972\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6975\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6972\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6964\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6964\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__6961\,
            I => \N__6955\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__6960\,
            I => \N__6952\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__6959\,
            I => \N__6949\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6946\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6943\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6940\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6937\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6946\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6943\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6940\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6937\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__6928\,
            I => \N__6925\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6921\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__6924\,
            I => \N__6918\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6915\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6910\
        );

    \I__1312\ : Span4Mux_s3_h
    port map (
            O => \N__6915\,
            I => \N__6907\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6904\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6901\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6910\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__6907\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6904\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6901\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__6892\,
            I => \N__6886\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__6891\,
            I => \N__6883\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6880\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6877\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6874\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6883\,
            I => \N__6871\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6880\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6877\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6874\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6871\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6859\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6859\,
            I => \N__6856\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__6856\,
            I => \N__6853\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__6853\,
            I => \VPP_VDDQ.N_1_i_12\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__6850\,
            I => \VPP_VDDQ.un9_clk_100khz_14_1_cascade_\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__6847\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_3_cascade_\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6841\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6841\,
            I => \N__6838\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__6838\,
            I => \VPP_VDDQ.count_2_RNI_0Z0Z_2\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6832\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6832\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6826\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6826\,
            I => \N__6822\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__6825\,
            I => \N__6819\
        );

    \I__1281\ : Span4Mux_s1_v
    port map (
            O => \N__6822\,
            I => \N__6815\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6812\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6809\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__6815\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6812\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6809\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__6802\,
            I => \VPP_VDDQ.count_2Z0Z_15_cascade_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6795\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6792\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6795\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6792\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6784\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6784\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__6781\,
            I => \VPP_VDDQ.un5_clk_100khz_cascade_\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__6778\,
            I => \VPP_VDDQ.count_2_1_5_cascade_\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6772\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6772\,
            I => \N__6769\
        );

    \I__1264\ : Span4Mux_v
    port map (
            O => \N__6769\,
            I => \N__6764\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6761\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6758\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__6764\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6761\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6758\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6748\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6748\,
            I => \N__6744\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__6747\,
            I => \N__6740\
        );

    \I__1255\ : Span4Mux_v
    port map (
            O => \N__6744\,
            I => \N__6737\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6734\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6731\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__6737\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6734\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6731\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6719\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6716\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6713\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6719\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6716\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6713\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6706\,
            I => \N__6703\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6703\,
            I => \N__6699\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6702\,
            I => \N__6695\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__6699\,
            I => \N__6692\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6689\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6695\,
            I => \N__6686\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__6692\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6689\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__6686\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__6679\,
            I => \VPP_VDDQ.un9_clk_100khz_4_1_cascade_\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__6676\,
            I => \VPP_VDDQ.count_2_1_8_cascade_\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6667\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6667\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6667\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__6664\,
            I => \VPP_VDDQ.count_2Z0Z_8_cascade_\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6658\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__6655\,
            I => \N__6651\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6648\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6645\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6648\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6645\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6637\,
            I => \VPP_VDDQ.count_2_0_5\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__6634\,
            I => \VPP_VDDQ.m4_cascade_\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6628\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6616\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6616\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6616\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__6613\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__6610\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0_cascade_\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__6607\,
            I => \VPP_VDDQ.m6_cascade_\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__6604\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6598\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6598\,
            I => \VPP_VDDQ.curr_state_2_e_0Z0Z_1\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6592\,
            I => \N__6588\
        );

    \I__1204\ : CEMux
    port map (
            O => \N__6591\,
            I => \N__6585\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__6588\,
            I => \N__6582\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6585\,
            I => \VPP_VDDQ.GZ0Z_76\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__6582\,
            I => \VPP_VDDQ.GZ0Z_76\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__6577\,
            I => \VPP_VDDQ.count_2_1_3_cascade_\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__6574\,
            I => \N__6570\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6562\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6570\,
            I => \N__6562\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6559\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6556\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__6567\,
            I => \N__6551\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6562\,
            I => \N__6541\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6541\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6538\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6535\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6532\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6527\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6527\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6520\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6520\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6520\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6517\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__6541\,
            I => \N__6514\
        );

    \I__1181\ : Span4Mux_v
    port map (
            O => \N__6538\,
            I => \N__6511\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6535\,
            I => \N__6500\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6532\,
            I => \N__6500\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6527\,
            I => \N__6500\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6500\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6517\,
            I => \N__6500\
        );

    \I__1175\ : Span4Mux_h
    port map (
            O => \N__6514\,
            I => \N__6497\
        );

    \I__1174\ : Span4Mux_h
    port map (
            O => \N__6511\,
            I => \N__6492\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__6500\,
            I => \N__6492\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__6497\,
            I => vddq_ok
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__6492\,
            I => vddq_ok
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__6487\,
            I => \N__6483\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6480\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6477\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6480\,
            I => \N__6470\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6477\,
            I => \N__6465\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6462\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6455\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6455\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6455\
        );

    \I__1161\ : Span4Mux_h
    port map (
            O => \N__6470\,
            I => \N__6452\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6469\,
            I => \N__6447\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6447\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__6465\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6462\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6455\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__6452\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6447\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1153\ : SRMux
    port map (
            O => \N__6436\,
            I => \N__6433\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1151\ : Span4Mux_h
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__6427\,
            I => \VPP_VDDQ.delayed_vddq_ok_RNOZ0\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6419\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__6423\,
            I => \N__6412\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6409\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6406\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6403\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6400\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6416\,
            I => \N__6395\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6395\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6392\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6409\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__6406\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6403\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6400\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6395\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6392\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__6379\,
            I => \N__6375\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__6378\,
            I => \N__6370\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6365\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6374\,
            I => \N__6362\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6355\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6355\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6355\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6352\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6365\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6362\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6355\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6352\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6340\,
            I => \N__6337\
        );

    \I__1120\ : Span4Mux_s3_h
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6334\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6325\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__6325\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6322\,
            I => \bfn_9_11_0_\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__1110\ : Sp12to4
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__6304\,
            I => v5a_ok
        );

    \I__1108\ : IoInMux
    port map (
            O => \N__6301\,
            I => \N__6298\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6298\,
            I => \N__6294\
        );

    \I__1106\ : IoInMux
    port map (
            O => \N__6297\,
            I => \N__6291\
        );

    \I__1105\ : IoSpan4Mux
    port map (
            O => \N__6294\,
            I => \N__6288\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6291\,
            I => \N__6285\
        );

    \I__1103\ : IoSpan4Mux
    port map (
            O => \N__6288\,
            I => \N__6280\
        );

    \I__1102\ : IoSpan4Mux
    port map (
            O => \N__6285\,
            I => \N__6280\
        );

    \I__1101\ : Span4Mux_s3_h
    port map (
            O => \N__6280\,
            I => \N__6276\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6273\
        );

    \I__1099\ : Span4Mux_h
    port map (
            O => \N__6276\,
            I => \N__6268\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6273\,
            I => \N__6268\
        );

    \I__1097\ : Span4Mux_h
    port map (
            O => \N__6268\,
            I => \N__6265\
        );

    \I__1096\ : Span4Mux_v
    port map (
            O => \N__6265\,
            I => \N__6262\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__6262\,
            I => v33a_ok
        );

    \I__1094\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__6253\,
            I => \N__6249\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__6252\,
            I => \N__6246\
        );

    \I__1090\ : Sp12to4
    port map (
            O => \N__6249\,
            I => \N__6243\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6240\
        );

    \I__1088\ : Span12Mux_s8_h
    port map (
            O => \N__6243\,
            I => \N__6235\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6235\
        );

    \I__1086\ : Odrv12
    port map (
            O => \N__6235\,
            I => slp_susn
        );

    \I__1085\ : IoInMux
    port map (
            O => \N__6232\,
            I => \N__6229\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6229\,
            I => \N__6226\
        );

    \I__1083\ : IoSpan4Mux
    port map (
            O => \N__6226\,
            I => \N__6222\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6219\
        );

    \I__1081\ : Span4Mux_s3_h
    port map (
            O => \N__6222\,
            I => \N__6214\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6219\,
            I => \N__6214\
        );

    \I__1079\ : Span4Mux_v
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__1078\ : Span4Mux_h
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__1077\ : Span4Mux_h
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__6205\,
            I => v1p8a_ok
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__6202\,
            I => \N__6198\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__6201\,
            I => \N__6195\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6188\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6188\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6182\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6182\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6188\,
            I => \N__6178\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__6187\,
            I => \N__6168\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6164\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6161\
        );

    \I__1065\ : Span4Mux_v
    port map (
            O => \N__6178\,
            I => \N__6158\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6151\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6151\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6151\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6174\,
            I => \N__6146\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6146\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6143\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6136\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6136\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6136\
        );

    \I__1055\ : Span4Mux_h
    port map (
            O => \N__6164\,
            I => \N__6131\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6161\,
            I => \N__6131\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__6158\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6151\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6146\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6143\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6136\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__6131\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__6118\,
            I => \VPP_VDDQ.count_2Z0Z_14_cascade_\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6109\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6109\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6109\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_THRU_CO\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6103\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6103\,
            I => \VPP_VDDQ.count_2_0_14\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6097\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1039\ : Odrv12
    port map (
            O => \N__6094\,
            I => \VPP_VDDQ.count_2_0_2\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6088\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6088\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6082\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6082\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6076\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6076\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6070\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6070\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6064\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6064\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6058\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__6058\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6055\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6052\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6044\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6041\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6038\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6044\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6041\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6038\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6028\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6028\,
            I => \N__6024\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6021\
        );

    \I__1015\ : Odrv12
    port map (
            O => \N__6024\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6021\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6012\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6009\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__6012\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6009\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6004\,
            I => \N__6001\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6001\,
            I => \VPP_VDDQ.count_2_1_12\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__5998\,
            I => \VPP_VDDQ.count_2_1_13_cascade_\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__5995\,
            I => \VPP_VDDQ.count_2Z0Z_13_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5986\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5986\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5986\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_THRU_CO\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5980\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__5977\,
            I => \VPP_VDDQ.count_2_1_14_cascade_\
        );

    \I__999\ : InMux
    port map (
            O => \N__5974\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__998\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5968\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5968\,
            I => \VPP_VDDQ.un1_count_2_1_axb_6\
        );

    \I__996\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5956\
        );

    \I__995\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5956\
        );

    \I__994\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5956\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5956\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVFZ0Z931\
        );

    \I__992\ : InMux
    port map (
            O => \N__5953\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__5950\,
            I => \N__5947\
        );

    \I__990\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5944\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__988\ : InMux
    port map (
            O => \N__5941\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__987\ : InMux
    port map (
            O => \N__5938\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__986\ : InMux
    port map (
            O => \N__5935\,
            I => \bfn_8_15_0_\
        );

    \I__985\ : InMux
    port map (
            O => \N__5932\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__983\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5922\
        );

    \I__982\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5919\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5922\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5919\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\
        );

    \I__979\ : InMux
    port map (
            O => \N__5914\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__978\ : InMux
    port map (
            O => \N__5911\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__977\ : InMux
    port map (
            O => \N__5908\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__5905\,
            I => \VPP_VDDQ.count_2_en_0_tz_cascade_\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__5902\,
            I => \VPP_VDDQ.count_2_en_cascade_\
        );

    \I__974\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5895\
        );

    \I__973\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5892\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5895\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5892\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__970\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5883\
        );

    \I__969\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5880\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5883\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__5880\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__5875\,
            I => \N__5871\
        );

    \I__965\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5868\
        );

    \I__964\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5865\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5868\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5865\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__961\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5856\
        );

    \I__960\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5853\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5856\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5853\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__957\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5844\
        );

    \I__956\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5841\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5844\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5841\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__953\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5832\
        );

    \I__952\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5829\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5832\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5829\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__5824\,
            I => \N__5820\
        );

    \I__948\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5817\
        );

    \I__947\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5814\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5817\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5814\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__944\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5805\
        );

    \I__943\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5802\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5805\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5802\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__940\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5790\
        );

    \I__938\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5787\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__5790\,
            I => \N__5782\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5787\,
            I => \N__5782\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__5782\,
            I => \VPP_VDDQ.un1_clk_100khz_1\
        );

    \I__934\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5772\
        );

    \I__932\ : InMux
    port map (
            O => \N__5775\,
            I => \N__5769\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__5772\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5769\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__929\ : InMux
    port map (
            O => \N__5764\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__928\ : InMux
    port map (
            O => \N__5761\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__927\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5755\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5755\,
            I => \VPP_VDDQ.un1_count_2_1_axb_4\
        );

    \I__925\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5749\,
            I => \N__5744\
        );

    \I__923\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5739\
        );

    \I__922\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5739\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__5744\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIRZ0Z9731\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5739\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIRZ0Z9731\
        );

    \I__919\ : InMux
    port map (
            O => \N__5734\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__918\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__5725\,
            I => \VPP_VDDQ.count_2_1_6\
        );

    \I__915\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5719\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5719\,
            I => \VPP_VDDQ.count_2_RNI25V3Z0Z_1\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5716\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIZ0_cascade_\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__5713\,
            I => \VPP_VDDQ.m4_1_cascade_\
        );

    \I__911\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5707\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5707\,
            I => \N__5702\
        );

    \I__909\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5697\
        );

    \I__908\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5697\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__5702\,
            I => \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5697\,
            I => \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__5692\,
            I => \N__5689\
        );

    \I__904\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5686\,
            I => \VPP_VDDQ.count_2_1_1\
        );

    \I__902\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__901\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5677\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__899\ : Span4Mux_s3_v
    port map (
            O => \N__5674\,
            I => \N__5670\
        );

    \I__898\ : InMux
    port map (
            O => \N__5673\,
            I => \N__5667\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__5670\,
            I => \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5667\,
            I => \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__5662\,
            I => \VPP_VDDQ.count_2_1_1_cascade_\
        );

    \I__894\ : InMux
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5656\,
            I => \VPP_VDDQ.count_2_1_4\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__5653\,
            I => \VPP_VDDQ.count_2_1_4_cascade_\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__5650\,
            I => \N__5646\
        );

    \I__890\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5642\
        );

    \I__889\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5637\
        );

    \I__888\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5637\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5642\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5637\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \N__5628\
        );

    \I__884\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5625\
        );

    \I__883\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5622\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5625\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5622\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__5617\,
            I => \N__5613\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__5616\,
            I => \N__5610\
        );

    \I__878\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5606\
        );

    \I__877\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5601\
        );

    \I__876\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5601\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5606\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5601\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__873\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5593\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__5590\,
            I => \N__5586\
        );

    \I__870\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5582\
        );

    \I__869\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5577\
        );

    \I__868\ : InMux
    port map (
            O => \N__5585\,
            I => \N__5577\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5582\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5577\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__865\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5568\
        );

    \I__864\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5565\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5568\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5565\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__861\ : InMux
    port map (
            O => \N__5560\,
            I => \N__5556\
        );

    \I__860\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5553\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5556\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5553\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__5548\,
            I => \N__5544\
        );

    \I__856\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5541\
        );

    \I__855\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5538\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5541\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5538\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__852\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5529\
        );

    \I__851\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5526\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5529\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5526\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__848\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5517\
        );

    \I__847\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5514\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5517\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5514\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__844\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5505\
        );

    \I__843\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5502\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5505\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5502\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__5497\,
            I => \N__5493\
        );

    \I__839\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5490\
        );

    \I__838\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5487\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5490\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5487\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__835\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5478\
        );

    \I__834\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5475\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5478\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5475\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__831\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5466\
        );

    \I__830\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5463\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5466\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5463\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__827\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5454\
        );

    \I__826\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5451\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5454\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5451\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__5446\,
            I => \N__5442\
        );

    \I__822\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5439\
        );

    \I__821\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5436\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5439\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5436\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__818\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5427\
        );

    \I__817\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5424\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5427\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5424\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__814\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5415\
        );

    \I__813\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5412\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5415\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5412\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__810\ : InMux
    port map (
            O => \N__5407\,
            I => \N__5403\
        );

    \I__809\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5400\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5403\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5400\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__5395\,
            I => \N__5391\
        );

    \I__805\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5388\
        );

    \I__804\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5385\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5388\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5385\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__801\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5376\
        );

    \I__800\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5373\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5376\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5373\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__5368\,
            I => \VPP_VDDQ.count_2_1_11_cascade_\
        );

    \I__796\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5362\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__794\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5356\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__792\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5350\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__790\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5342\
        );

    \I__789\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5337\
        );

    \I__788\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5337\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5342\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5337\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__785\ : InMux
    port map (
            O => \N__5332\,
            I => \N__5327\
        );

    \I__784\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5324\
        );

    \I__783\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5321\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5327\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5324\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5321\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__779\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5308\
        );

    \I__778\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5305\
        );

    \I__777\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5300\
        );

    \I__776\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5300\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5308\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5305\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5300\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__772\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__5287\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__5284\,
            I => \N__5279\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__5283\,
            I => \N__5276\
        );

    \I__767\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5273\
        );

    \I__766\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5268\
        );

    \I__765\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5268\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5273\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5268\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__762\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5260\,
            I => \VPP_VDDQ.N_6\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__5257\,
            I => \VPP_VDDQ.count_2_1_6_cascade_\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__5254\,
            I => \VPP_VDDQ.count_2Z0Z_12_cascade_\
        );

    \I__758\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5248\,
            I => \VPP_VDDQ.count_2_0_12\
        );

    \I__756\ : InMux
    port map (
            O => \N__5245\,
            I => \bfn_7_13_0_\
        );

    \I__755\ : InMux
    port map (
            O => \N__5242\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__754\ : InMux
    port map (
            O => \N__5239\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__753\ : InMux
    port map (
            O => \N__5236\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__752\ : InMux
    port map (
            O => \N__5233\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__751\ : InMux
    port map (
            O => \N__5230\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__750\ : InMux
    port map (
            O => \N__5227\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__5224\,
            I => \VPP_VDDQ.g0_3_a3_0_1_cascade_\
        );

    \I__748\ : InMux
    port map (
            O => \N__5221\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__747\ : InMux
    port map (
            O => \N__5218\,
            I => \bfn_7_12_0_\
        );

    \I__746\ : InMux
    port map (
            O => \N__5215\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__745\ : InMux
    port map (
            O => \N__5212\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__744\ : InMux
    port map (
            O => \N__5209\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__743\ : InMux
    port map (
            O => \N__5206\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__742\ : InMux
    port map (
            O => \N__5203\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__741\ : InMux
    port map (
            O => \N__5200\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__740\ : InMux
    port map (
            O => \N__5197\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__739\ : InMux
    port map (
            O => \N__5194\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__738\ : InMux
    port map (
            O => \N__5191\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__737\ : InMux
    port map (
            O => \N__5188\,
            I => \bfn_7_11_0_\
        );

    \I__736\ : InMux
    port map (
            O => \N__5185\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__735\ : InMux
    port map (
            O => \N__5182\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__734\ : InMux
    port map (
            O => \N__5179\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__733\ : InMux
    port map (
            O => \N__5176\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__732\ : InMux
    port map (
            O => \N__5173\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__731\ : InMux
    port map (
            O => \N__5170\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__730\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5164\,
            I => \VPP_VDDQ.delayed_vddq_ok_en\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__5161\,
            I => \N__5157\
        );

    \I__727\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5154\
        );

    \I__726\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5151\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5154\,
            I => \VPP_VDDQ.delayed_vddq_ok_0\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5151\,
            I => \VPP_VDDQ.delayed_vddq_ok_0\
        );

    \I__723\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5143\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5143\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__721\ : InMux
    port map (
            O => \N__5140\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__720\ : InMux
    port map (
            O => \N__5137\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__719\ : InMux
    port map (
            O => \N__5134\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__718\ : InMux
    port map (
            O => \N__5131\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__717\ : InMux
    port map (
            O => \N__5128\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__716\ : InMux
    port map (
            O => \N__5125\,
            I => \PCH_PWRGD.un1_count_1_cry_9\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__5122\,
            I => \N__5118\
        );

    \I__714\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5115\
        );

    \I__713\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5112\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5115\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5112\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__710\ : InMux
    port map (
            O => \N__5107\,
            I => \PCH_PWRGD.un1_count_1_cry_10\
        );

    \I__709\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5100\
        );

    \I__708\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5097\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5100\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5097\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__705\ : InMux
    port map (
            O => \N__5092\,
            I => \PCH_PWRGD.un1_count_1_cry_11\
        );

    \I__704\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5085\
        );

    \I__703\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5082\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5085\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5082\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__700\ : InMux
    port map (
            O => \N__5077\,
            I => \PCH_PWRGD.un1_count_1_cry_12\
        );

    \I__699\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5070\
        );

    \I__698\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5067\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5070\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5067\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__695\ : InMux
    port map (
            O => \N__5062\,
            I => \PCH_PWRGD.un1_count_1_cry_13\
        );

    \I__694\ : InMux
    port map (
            O => \N__5059\,
            I => \bfn_6_11_0_\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__5056\,
            I => \N__5052\
        );

    \I__692\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__691\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5046\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5049\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5046\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__688\ : CEMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5038\,
            I => \N__5035\
        );

    \I__686\ : Odrv12
    port map (
            O => \N__5035\,
            I => \PCH_PWRGD.N_15_2\
        );

    \I__685\ : SRMux
    port map (
            O => \N__5032\,
            I => \N__5028\
        );

    \I__684\ : SRMux
    port map (
            O => \N__5031\,
            I => \N__5024\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5028\,
            I => \N__5021\
        );

    \I__682\ : SRMux
    port map (
            O => \N__5027\,
            I => \N__5018\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__5014\
        );

    \I__680\ : Span4Mux_h
    port map (
            O => \N__5021\,
            I => \N__5009\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5018\,
            I => \N__5009\
        );

    \I__678\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5006\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__5014\,
            I => \G_12\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__5009\,
            I => \G_12\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5006\,
            I => \G_12\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__4999\,
            I => \VPP_VDDQ.delayed_vddq_ok_en_cascade_\
        );

    \I__673\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4993\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4993\,
            I => \N__4990\
        );

    \I__671\ : Odrv12
    port map (
            O => \N__4990\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__670\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4983\
        );

    \I__669\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4980\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4983\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4980\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__666\ : InMux
    port map (
            O => \N__4975\,
            I => \PCH_PWRGD.un1_count_1_cry_1\
        );

    \I__665\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4968\
        );

    \I__664\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4965\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4968\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4965\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__661\ : InMux
    port map (
            O => \N__4960\,
            I => \PCH_PWRGD.un1_count_1_cry_2\
        );

    \I__660\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4953\
        );

    \I__659\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4950\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4953\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4950\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__656\ : InMux
    port map (
            O => \N__4945\,
            I => \PCH_PWRGD.un1_count_1_cry_3\
        );

    \I__655\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4938\
        );

    \I__654\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4935\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4938\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4935\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__651\ : InMux
    port map (
            O => \N__4930\,
            I => \PCH_PWRGD.un1_count_1_cry_4\
        );

    \I__650\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4923\
        );

    \I__649\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4920\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4923\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4920\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__646\ : InMux
    port map (
            O => \N__4915\,
            I => \PCH_PWRGD.un1_count_1_cry_5\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__4912\,
            I => \N__4908\
        );

    \I__644\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4905\
        );

    \I__643\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4902\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4905\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4902\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__640\ : InMux
    port map (
            O => \N__4897\,
            I => \PCH_PWRGD.un1_count_1_cry_6\
        );

    \I__639\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4890\
        );

    \I__638\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4887\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4890\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__4887\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__635\ : InMux
    port map (
            O => \N__4882\,
            I => \bfn_6_10_0_\
        );

    \I__634\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4875\
        );

    \I__633\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4872\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4869\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4872\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__4869\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__629\ : InMux
    port map (
            O => \N__4864\,
            I => \PCH_PWRGD.un1_count_1_cry_8\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__4861\,
            I => \N__4857\
        );

    \I__627\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4854\
        );

    \I__626\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4851\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4854\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4851\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__4846\,
            I => \PCH_PWRGD.delayed_vccin_ok_s_1_cascade_\
        );

    \I__622\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4834\
        );

    \I__621\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4834\
        );

    \I__620\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4834\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4834\,
            I => \PCH_PWRGD.delayed_vccin_okZ0\
        );

    \I__618\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4814\
        );

    \I__617\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4814\
        );

    \I__616\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4814\
        );

    \I__615\ : InMux
    port map (
            O => \N__4828\,
            I => \N__4814\
        );

    \I__614\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4814\
        );

    \I__613\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4809\
        );

    \I__612\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4809\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4814\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4809\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__609\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4788\
        );

    \I__608\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4788\
        );

    \I__607\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4788\
        );

    \I__606\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4788\
        );

    \I__605\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4788\
        );

    \I__604\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4785\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4788\,
            I => \VPP_VDDQ.curr_stateZ1Z_0\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4785\,
            I => \VPP_VDDQ.curr_stateZ1Z_0\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__600\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4774\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4774\,
            I => \VPP_VDDQ.curr_state12\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__4771\,
            I => \N__4766\
        );

    \I__597\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4760\
        );

    \I__596\ : InMux
    port map (
            O => \N__4769\,
            I => \N__4760\
        );

    \I__595\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4755\
        );

    \I__594\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4755\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4760\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4755\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__591\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4747\,
            I => \N__4742\
        );

    \I__589\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4737\
        );

    \I__588\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4737\
        );

    \I__587\ : Odrv4
    port map (
            O => \N__4742\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4737\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__585\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4726\
        );

    \I__584\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4723\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__4730\,
            I => \N__4718\
        );

    \I__582\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4715\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4726\,
            I => \N__4710\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4723\,
            I => \N__4710\
        );

    \I__579\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4703\
        );

    \I__578\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4703\
        );

    \I__577\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4703\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4715\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__4710\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4703\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__4696\,
            I => \PCH_PWRGD.i3_mux_0_cascade_\
        );

    \I__572\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4685\
        );

    \I__571\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4682\
        );

    \I__570\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4677\
        );

    \I__569\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4677\
        );

    \I__568\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4672\
        );

    \I__567\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4672\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4685\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4682\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4677\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4672\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__562\ : IoInMux
    port map (
            O => \N__4663\,
            I => \N__4659\
        );

    \I__561\ : IoInMux
    port map (
            O => \N__4662\,
            I => \N__4655\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4659\,
            I => \N__4652\
        );

    \I__559\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4649\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4655\,
            I => \N__4646\
        );

    \I__557\ : Span4Mux_s3_h
    port map (
            O => \N__4652\,
            I => \N__4643\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4640\
        );

    \I__555\ : Span12Mux_s4_h
    port map (
            O => \N__4646\,
            I => \N__4637\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__4643\,
            I => \N__4634\
        );

    \I__553\ : Span4Mux_v
    port map (
            O => \N__4640\,
            I => \N__4631\
        );

    \I__552\ : Odrv12
    port map (
            O => \N__4637\,
            I => pch_pwrok
        );

    \I__551\ : Odrv4
    port map (
            O => \N__4634\,
            I => pch_pwrok
        );

    \I__550\ : Odrv4
    port map (
            O => \N__4631\,
            I => pch_pwrok
        );

    \I__549\ : IoInMux
    port map (
            O => \N__4624\,
            I => \N__4621\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__547\ : Odrv12
    port map (
            O => \N__4618\,
            I => vccst_pwrgd
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__545\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4608\
        );

    \I__544\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4605\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4608\,
            I => \N__4602\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4605\,
            I => \N__4599\
        );

    \I__541\ : Span4Mux_h
    port map (
            O => \N__4602\,
            I => \N__4596\
        );

    \I__540\ : Odrv4
    port map (
            O => \N__4599\,
            I => \PCH_PWRGD.un1_curr_state10_0\
        );

    \I__539\ : Odrv4
    port map (
            O => \N__4596\,
            I => \PCH_PWRGD.un1_curr_state10_0\
        );

    \I__538\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4587\
        );

    \I__537\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4584\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4587\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4584\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__534\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4575\
        );

    \I__533\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4572\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4575\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4572\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__530\ : InMux
    port map (
            O => \N__4567\,
            I => \PCH_PWRGD.un1_count_1_cry_0\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__4564\,
            I => \PCH_PWRGD_un1_delayed_vccin_ok_0_sqmuxa_0_cascade_\
        );

    \I__528\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4558\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__526\ : Span4Mux_v
    port map (
            O => \N__4555\,
            I => \N__4552\
        );

    \I__525\ : Span4Mux_h
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__524\ : Odrv4
    port map (
            O => \N__4549\,
            I => vr_ready_vccin
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__4546\,
            I => \PCH_PWRGD.N_3_i_cascade_\
        );

    \I__522\ : CEMux
    port map (
            O => \N__4543\,
            I => \N__4540\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__520\ : Odrv4
    port map (
            O => \N__4537\,
            I => \VPP_VDDQ.N_15_0\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__4534\,
            I => \PCH_PWRGD.N_6_cascade_\
        );

    \I__518\ : SRMux
    port map (
            O => \N__4531\,
            I => \N__4527\
        );

    \I__517\ : SRMux
    port map (
            O => \N__4530\,
            I => \N__4524\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4527\,
            I => \N__4520\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4517\
        );

    \I__514\ : SRMux
    port map (
            O => \N__4523\,
            I => \N__4514\
        );

    \I__513\ : Span4Mux_v
    port map (
            O => \N__4520\,
            I => \N__4506\
        );

    \I__512\ : Span4Mux_h
    port map (
            O => \N__4517\,
            I => \N__4506\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4514\,
            I => \N__4506\
        );

    \I__510\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4503\
        );

    \I__509\ : Odrv4
    port map (
            O => \N__4506\,
            I => \VPP_VDDQ.curr_state_RNI0TJM7Z0Z_0\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4503\,
            I => \VPP_VDDQ.curr_state_RNI0TJM7Z0Z_0\
        );

    \I__507\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4493\
        );

    \I__506\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4488\
        );

    \I__505\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4488\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4493\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_1_sqmuxa\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4488\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_1_sqmuxa\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__501\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4474\
        );

    \I__500\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4474\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__4471\,
            I => \VPP_VDDQ.un6_count\
        );

    \I__497\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4464\
        );

    \I__496\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4461\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4464\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4461\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__493\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4452\
        );

    \I__492\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4449\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4452\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4449\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__4444\,
            I => \N__4440\
        );

    \I__488\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4437\
        );

    \I__487\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4434\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4437\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4434\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__484\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4425\
        );

    \I__483\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4422\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4425\,
            I => \N__4419\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4422\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__480\ : Odrv4
    port map (
            O => \N__4419\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__479\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4411\,
            I => \N__4408\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__4408\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__476\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4401\
        );

    \I__475\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4398\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4401\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4398\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__472\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4389\
        );

    \I__471\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4386\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4389\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4386\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__4381\,
            I => \N__4378\
        );

    \I__467\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4374\
        );

    \I__466\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4371\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4374\,
            I => \N__4368\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4371\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__463\ : Odrv4
    port map (
            O => \N__4368\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__462\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4359\
        );

    \I__461\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4356\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4359\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4356\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__458\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4348\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4348\,
            I => \VPP_VDDQ.un6_count_9\
        );

    \I__456\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4342\,
            I => \PCH_PWRGD.un4_count_11\
        );

    \I__454\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4336\,
            I => \PCH_PWRGD.un4_count_10\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__4333\,
            I => \PCH_PWRGD.un4_count_8_cascade_\
        );

    \I__451\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4327\,
            I => \PCH_PWRGD.un4_count_9\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4324\,
            I => \VPP_VDDQ.un1_vddq_pwrgdZ0_cascade_\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__4321\,
            I => \N__4317\
        );

    \I__447\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4314\
        );

    \I__446\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4311\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4314\,
            I => \N__4306\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4311\,
            I => \N__4306\
        );

    \I__443\ : Odrv12
    port map (
            O => \N__4306\,
            I => \VPP_VDDQ.un1_curr_state13_0\
        );

    \I__442\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4295\
        );

    \I__441\ : InMux
    port map (
            O => \N__4302\,
            I => \N__4295\
        );

    \I__440\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4290\
        );

    \I__439\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4290\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4295\,
            I => \VPP_VDDQ.un1_vddq_pwrgdZ0\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4290\,
            I => \VPP_VDDQ.un1_vddq_pwrgdZ0\
        );

    \I__436\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4282\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4282\,
            I => \N__4278\
        );

    \I__434\ : InMux
    port map (
            O => \N__4281\,
            I => \N__4275\
        );

    \I__433\ : Sp12to4
    port map (
            O => \N__4278\,
            I => \N__4270\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4275\,
            I => \N__4270\
        );

    \I__431\ : Odrv12
    port map (
            O => \N__4270\,
            I => slp_s4n
        );

    \I__430\ : IoInMux
    port map (
            O => \N__4267\,
            I => \N__4264\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4264\,
            I => \N__4261\
        );

    \I__428\ : IoSpan4Mux
    port map (
            O => \N__4261\,
            I => \N__4257\
        );

    \I__427\ : InMux
    port map (
            O => \N__4260\,
            I => \N__4254\
        );

    \I__426\ : Span4Mux_s0_h
    port map (
            O => \N__4257\,
            I => \N__4249\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__4254\,
            I => \N__4249\
        );

    \I__424\ : Odrv4
    port map (
            O => \N__4249\,
            I => vccst_en
        );

    \I__423\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4242\
        );

    \I__422\ : InMux
    port map (
            O => \N__4245\,
            I => \N__4239\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4242\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4239\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__4234\,
            I => \vccst_en_cascade_\
        );

    \I__418\ : IoInMux
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__416\ : Odrv12
    port map (
            O => \N__4225\,
            I => vpp_en
        );

    \I__415\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4218\
        );

    \I__414\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4215\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4218\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4215\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__411\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4206\
        );

    \I__410\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4203\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4206\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4203\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__4198\,
            I => \N__4194\
        );

    \I__406\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4191\
        );

    \I__405\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4188\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4191\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4188\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__402\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4179\
        );

    \I__401\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4176\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4179\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4176\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__398\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4167\
        );

    \I__397\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4164\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4167\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4164\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__394\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4155\
        );

    \I__393\ : InMux
    port map (
            O => \N__4158\,
            I => \N__4152\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__4155\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__4152\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__389\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4140\
        );

    \I__388\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4137\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4134\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4137\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__385\ : Odrv4
    port map (
            O => \N__4134\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__384\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4125\
        );

    \I__383\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4122\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__4125\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__4122\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__380\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4114\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4114\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__4111\,
            I => \VPP_VDDQ.un6_count_8_cascade_\
        );

    \I__377\ : InMux
    port map (
            O => \N__4108\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__376\ : InMux
    port map (
            O => \N__4105\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__375\ : InMux
    port map (
            O => \N__4102\,
            I => \bfn_4_11_0_\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__4099\,
            I => \VPP_VDDQ.un1_curr_state12_0_cascade_\
        );

    \I__373\ : CascadeMux
    port map (
            O => \N__4096\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\
        );

    \I__372\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__4090\,
            I => \VPP_VDDQ.curr_state11\
        );

    \I__370\ : InMux
    port map (
            O => \N__4087\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__369\ : InMux
    port map (
            O => \N__4084\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__368\ : InMux
    port map (
            O => \N__4081\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__367\ : InMux
    port map (
            O => \N__4078\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__366\ : InMux
    port map (
            O => \N__4075\,
            I => \bfn_4_10_0_\
        );

    \I__365\ : InMux
    port map (
            O => \N__4072\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__364\ : InMux
    port map (
            O => \N__4069\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__363\ : InMux
    port map (
            O => \N__4066\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__362\ : InMux
    port map (
            O => \N__4063\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__361\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4057\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__4057\,
            I => vpp_ok
        );

    \I__359\ : IoInMux
    port map (
            O => \N__4054\,
            I => \N__4051\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__4051\,
            I => \N__4048\
        );

    \I__357\ : Odrv12
    port map (
            O => \N__4048\,
            I => vddq_en
        );

    \I__356\ : IoInMux
    port map (
            O => \N__4045\,
            I => \N__4042\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__4039\,
            I => v33a_enn
        );

    \I__353\ : IoInMux
    port map (
            O => \N__4036\,
            I => \N__4033\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__4033\,
            I => \N__4029\
        );

    \I__351\ : IoInMux
    port map (
            O => \N__4032\,
            I => \N__4026\
        );

    \I__350\ : Span4Mux_s1_h
    port map (
            O => \N__4029\,
            I => \N__4023\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__4026\,
            I => \N__4020\
        );

    \I__348\ : Odrv4
    port map (
            O => \N__4023\,
            I => v5s_enn
        );

    \I__347\ : Odrv4
    port map (
            O => \N__4020\,
            I => v5s_enn
        );

    \I__346\ : InMux
    port map (
            O => \N__4015\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__345\ : InMux
    port map (
            O => \N__4012\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__344\ : InMux
    port map (
            O => \N__4009\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_6_11_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4060\,
            in2 => \_gnd_net_\,
            in3 => \N__4260\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_SUSn_RNIN4K9_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6259\,
            lcout => v33a_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.slp_s3n_signal_i_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__7105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7809\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9103\,
            in1 => \N__4428\,
            in2 => \N__4321\,
            in3 => \N__4320\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_1_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9094\,
            in1 => \N__4159\,
            in2 => \_gnd_net_\,
            in3 => \N__4015\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9104\,
            in1 => \N__4129\,
            in2 => \_gnd_net_\,
            in3 => \N__4012\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_3_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9095\,
            in1 => \N__4222\,
            in2 => \_gnd_net_\,
            in3 => \N__4009\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_4_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9105\,
            in1 => \N__4183\,
            in2 => \_gnd_net_\,
            in3 => \N__4087\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_5_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9096\,
            in1 => \N__4210\,
            in2 => \_gnd_net_\,
            in3 => \N__4084\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_6_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9106\,
            in1 => \N__4171\,
            in2 => \_gnd_net_\,
            in3 => \N__4081\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_7_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9097\,
            in1 => \N__4197\,
            in2 => \_gnd_net_\,
            in3 => \N__4078\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__8677\,
            ce => 'H',
            sr => \N__4531\
        );

    \VPP_VDDQ.count_8_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9079\,
            in1 => \N__4456\,
            in2 => \_gnd_net_\,
            in3 => \N__4075\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__4530\
        );

    \VPP_VDDQ.count_9_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9075\,
            in1 => \N__4468\,
            in2 => \_gnd_net_\,
            in3 => \N__4072\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__4530\
        );

    \VPP_VDDQ.count_10_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9076\,
            in1 => \N__4143\,
            in2 => \_gnd_net_\,
            in3 => \N__4069\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__4530\
        );

    \VPP_VDDQ.count_11_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9073\,
            in1 => \N__4443\,
            in2 => \_gnd_net_\,
            in3 => \N__4066\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__4530\
        );

    \VPP_VDDQ.count_12_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9077\,
            in1 => \N__4363\,
            in2 => \_gnd_net_\,
            in3 => \N__4063\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__4530\
        );

    \VPP_VDDQ.count_13_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9074\,
            in1 => \N__4393\,
            in2 => \_gnd_net_\,
            in3 => \N__4108\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__4530\
        );

    \VPP_VDDQ.count_14_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9078\,
            in1 => \N__4405\,
            in2 => \_gnd_net_\,
            in3 => \N__4105\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__4530\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7207\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4377\,
            in2 => \_gnd_net_\,
            in3 => \N__4102\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8737\,
            ce => \N__4543\,
            sr => \N__4523\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_2_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__4829\,
            in1 => \N__4802\,
            in2 => \_gnd_net_\,
            in3 => \N__4301\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_curr_state12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001110"
        )
    port map (
            in0 => \N__9080\,
            in1 => \N__4245\,
            in2 => \N__4099\,
            in3 => \N__4498\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__4303\,
            in1 => \N__4093\,
            in2 => \N__4096\,
            in3 => \N__9084\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4803\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4830\,
            lcout => \VPP_VDDQ.curr_state11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIDNTT1_0_0_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4827\,
            in1 => \N__4800\,
            in2 => \_gnd_net_\,
            in3 => \N__4300\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgd_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_pwrgd_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6568\,
            in1 => \N__4285\,
            in2 => \_gnd_net_\,
            in3 => \N__7800\,
            lcout => \VPP_VDDQ.un1_vddq_pwrgdZ0\,
            ltout => \VPP_VDDQ.un1_vddq_pwrgdZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__4828\,
            in1 => \_gnd_net_\,
            in2 => \N__4324\,
            in3 => \N__4801\,
            lcout => \VPP_VDDQ.un1_curr_state13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__4804\,
            in1 => \N__4831\,
            in2 => \N__9102\,
            in3 => \N__4302\,
            lcout => \VPP_VDDQ.curr_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.VCCST_EN_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7805\,
            lcout => vccst_en,
            ltout => \vccst_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__4246\,
            in1 => \_gnd_net_\,
            in2 => \N__4234\,
            in3 => \_gnd_net_\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4221\,
            in1 => \N__4209\,
            in2 => \N__4198\,
            in3 => \N__4182\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4170\,
            in1 => \N__4158\,
            in2 => \N__4147\,
            in3 => \N__4128\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4414\,
            in1 => \N__4117\,
            in2 => \N__4111\,
            in3 => \N__4351\,
            lcout => \VPP_VDDQ.un6_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI7J2B_3_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4941\,
            in1 => \N__4956\,
            in2 => \N__4912\,
            in3 => \N__4971\,
            lcout => \PCH_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIESHJ_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4926\,
            in1 => \N__4986\,
            in2 => \N__4861\,
            in3 => \N__4578\,
            lcout => \PCH_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIN5IJ_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4879\,
            in1 => \N__4590\,
            in2 => \N__5122\,
            in3 => \N__4893\,
            lcout => \PCH_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4467\,
            in1 => \N__4455\,
            in2 => \N__4444\,
            in3 => \N__4429\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4404\,
            in1 => \N__4392\,
            in2 => \N__4381\,
            in3 => \N__4362\,
            lcout => \VPP_VDDQ.un6_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIFR521_15_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5073\,
            in1 => \N__5088\,
            in2 => \N__5056\,
            in3 => \N__5103\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un4_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4345\,
            in1 => \N__4339\,
            in2 => \N__4333\,
            in3 => \N__4330\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNO_0_15_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8902\,
            in2 => \_gnd_net_\,
            in3 => \N__5017\,
            lcout => \PCH_PWRGD.N_15_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI1LNN4_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__4688\,
            in1 => \N__4765\,
            in2 => \N__4730\,
            in3 => \N__4745\,
            lcout => OPEN,
            ltout => \PCH_PWRGD_un1_delayed_vccin_ok_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.G_12_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4564\,
            in3 => \N__8901\,
            lcout => \G_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_vccin_ok_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4561\,
            in1 => \N__7101\,
            in2 => \_gnd_net_\,
            in3 => \N__7793\,
            lcout => \PCH_PWRGD.N_3_i\,
            ltout => \PCH_PWRGD.N_3_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI64B32_0_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4721\,
            in2 => \N__4546\,
            in3 => \N__4689\,
            lcout => \PCH_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__8903\,
            in1 => \N__4513\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.N_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m5_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__4746\,
            in1 => \_gnd_net_\,
            in2 => \N__4771\,
            in3 => \N__4722\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__8904\,
            in1 => \N__4729\,
            in2 => \N__4534\,
            in3 => \N__4693\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI0TJM7_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__4496\,
            in1 => \N__4479\,
            in2 => \N__4780\,
            in3 => \N__8981\,
            lcout => \VPP_VDDQ.curr_state_RNI0TJM7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001000"
        )
    port map (
            in0 => \N__8983\,
            in1 => \N__4497\,
            in2 => \N__4483\,
            in3 => \N__4826\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI6LSN_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4843\,
            in1 => \N__7100\,
            in2 => \_gnd_net_\,
            in3 => \N__7801\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNO_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110111011"
        )
    port map (
            in0 => \N__4691\,
            in1 => \N__4841\,
            in2 => \_gnd_net_\,
            in3 => \N__4769\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.delayed_vccin_ok_s_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__4842\,
            in1 => \N__4731\,
            in2 => \N__4846\,
            in3 => \N__8984\,
            lcout => \PCH_PWRGD.delayed_vccin_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNID2IU_0_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4825\,
            in2 => \_gnd_net_\,
            in3 => \N__4799\,
            lcout => \VPP_VDDQ.curr_state12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m3_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4770\,
            in1 => \N__4690\,
            in2 => \_gnd_net_\,
            in3 => \N__4750\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.i3_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010110000000"
        )
    port map (
            in0 => \N__8982\,
            in1 => \N__4732\,
            in2 => \N__4696\,
            in3 => \N__4692\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNIQST72_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4658\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4996\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9065\,
            in1 => \N__4591\,
            in2 => \N__4615\,
            in3 => \N__4611\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_0\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9069\,
            in1 => \N__4579\,
            in2 => \_gnd_net_\,
            in3 => \N__4567\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_0\,
            carryout => \PCH_PWRGD.un1_count_1_cry_1\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9066\,
            in1 => \N__4987\,
            in2 => \_gnd_net_\,
            in3 => \N__4975\,
            lcout => \PCH_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_1\,
            carryout => \PCH_PWRGD.un1_count_1_cry_2\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9070\,
            in1 => \N__4972\,
            in2 => \_gnd_net_\,
            in3 => \N__4960\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_2\,
            carryout => \PCH_PWRGD.un1_count_1_cry_3\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_4_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9067\,
            in1 => \N__4957\,
            in2 => \_gnd_net_\,
            in3 => \N__4945\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_3\,
            carryout => \PCH_PWRGD.un1_count_1_cry_4\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_5_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9071\,
            in1 => \N__4942\,
            in2 => \_gnd_net_\,
            in3 => \N__4930\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_4\,
            carryout => \PCH_PWRGD.un1_count_1_cry_5\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_6_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9068\,
            in1 => \N__4927\,
            in2 => \_gnd_net_\,
            in3 => \N__4915\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_5\,
            carryout => \PCH_PWRGD.un1_count_1_cry_6\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_7_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9072\,
            in1 => \N__4911\,
            in2 => \_gnd_net_\,
            in3 => \N__4897\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_6\,
            carryout => \PCH_PWRGD.un1_count_1_cry_7\,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__5031\
        );

    \PCH_PWRGD.count_8_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9041\,
            in1 => \N__4894\,
            in2 => \_gnd_net_\,
            in3 => \N__4882\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_8\,
            clk => \N__8682\,
            ce => 'H',
            sr => \N__5032\
        );

    \PCH_PWRGD.count_9_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9044\,
            in1 => \N__4878\,
            in2 => \_gnd_net_\,
            in3 => \N__4864\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_8\,
            carryout => \PCH_PWRGD.un1_count_1_cry_9\,
            clk => \N__8682\,
            ce => 'H',
            sr => \N__5032\
        );

    \PCH_PWRGD.count_10_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9038\,
            in1 => \N__4860\,
            in2 => \_gnd_net_\,
            in3 => \N__5125\,
            lcout => \PCH_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_9\,
            carryout => \PCH_PWRGD.un1_count_1_cry_10\,
            clk => \N__8682\,
            ce => 'H',
            sr => \N__5032\
        );

    \PCH_PWRGD.count_11_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9042\,
            in1 => \N__5121\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_10\,
            carryout => \PCH_PWRGD.un1_count_1_cry_11\,
            clk => \N__8682\,
            ce => 'H',
            sr => \N__5032\
        );

    \PCH_PWRGD.count_12_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9039\,
            in1 => \N__5104\,
            in2 => \_gnd_net_\,
            in3 => \N__5092\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_11\,
            carryout => \PCH_PWRGD.un1_count_1_cry_12\,
            clk => \N__8682\,
            ce => 'H',
            sr => \N__5032\
        );

    \PCH_PWRGD.count_13_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9043\,
            in1 => \N__5089\,
            in2 => \_gnd_net_\,
            in3 => \N__5077\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_12\,
            carryout => \PCH_PWRGD.un1_count_1_cry_13\,
            clk => \N__8682\,
            ce => 'H',
            sr => \N__5032\
        );

    \PCH_PWRGD.count_14_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9040\,
            in1 => \N__5074\,
            in2 => \_gnd_net_\,
            in3 => \N__5062\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_13\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14\,
            clk => \N__8682\,
            ce => 'H',
            sr => \N__5032\
        );

    \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7195\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_14\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_15_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5055\,
            in2 => \_gnd_net_\,
            in3 => \N__5059\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8679\,
            ce => \N__5041\,
            sr => \N__5027\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIJCTQ_1_1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__6595\,
            in1 => \N__6424\,
            in2 => \N__6574\,
            in3 => \N__8244\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_en\,
            ltout => \VPP_VDDQ.delayed_vddq_ok_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNIK71G1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__5160\,
            in1 => \N__6573\,
            in2 => \N__4999\,
            in3 => \N__5797\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__6569\,
            in1 => \N__5793\,
            in2 => \N__5161\,
            in3 => \N__5167\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8681\,
            ce => 'H',
            sr => \N__6436\
        );

    \COUNTER.counter_2_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5146\,
            in1 => \N__5332\,
            in2 => \_gnd_net_\,
            in3 => \N__6193\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5314\,
            in2 => \_gnd_net_\,
            in3 => \N__6194\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5313\,
            in2 => \N__5617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5331\,
            in2 => \_gnd_net_\,
            in3 => \N__5140\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5347\,
            in2 => \_gnd_net_\,
            in3 => \N__5137\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5282\,
            in2 => \_gnd_net_\,
            in3 => \N__5134\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5589\,
            in2 => \_gnd_net_\,
            in3 => \N__5131\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5649\,
            in2 => \_gnd_net_\,
            in3 => \N__5128\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5631\,
            in2 => \_gnd_net_\,
            in3 => \N__5194\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__8661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5431\,
            in2 => \_gnd_net_\,
            in3 => \N__5191\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__8661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5458\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5470\,
            in2 => \_gnd_net_\,
            in3 => \N__5185\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5445\,
            in2 => \_gnd_net_\,
            in3 => \N__5182\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5380\,
            in2 => \_gnd_net_\,
            in3 => \N__5179\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5419\,
            in2 => \_gnd_net_\,
            in3 => \N__5176\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5407\,
            in2 => \_gnd_net_\,
            in3 => \N__5173\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5394\,
            in2 => \_gnd_net_\,
            in3 => \N__5170\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5533\,
            in2 => \_gnd_net_\,
            in3 => \N__5221\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5560\,
            in2 => \_gnd_net_\,
            in3 => \N__5218\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5572\,
            in2 => \_gnd_net_\,
            in3 => \N__5215\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5547\,
            in2 => \_gnd_net_\,
            in3 => \N__5212\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5482\,
            in2 => \_gnd_net_\,
            in3 => \N__5209\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5509\,
            in2 => \_gnd_net_\,
            in3 => \N__5206\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5521\,
            in2 => \_gnd_net_\,
            in3 => \N__5203\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5496\,
            in2 => \_gnd_net_\,
            in3 => \N__5200\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5809\,
            in2 => \_gnd_net_\,
            in3 => \N__5197\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__8683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5836\,
            in2 => \_gnd_net_\,
            in3 => \N__5245\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5848\,
            in2 => \_gnd_net_\,
            in3 => \N__5242\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5823\,
            in2 => \_gnd_net_\,
            in3 => \N__5239\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5860\,
            in2 => \_gnd_net_\,
            in3 => \N__5236\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5887\,
            in2 => \_gnd_net_\,
            in3 => \N__5233\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5899\,
            in2 => \_gnd_net_\,
            in3 => \N__5230\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5874\,
            in2 => \_gnd_net_\,
            in3 => \N__5227\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI25V3_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6722\,
            in1 => \N__6767\,
            in2 => \N__6747\,
            in3 => \N__6702\,
            lcout => \VPP_VDDQ.count_2_RNI25V3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIMO1Q2_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5748\,
            in1 => \N__5683\,
            in2 => \N__6202\,
            in3 => \N__5710\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.g0_3_a3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI98JR5_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__5964\,
            in1 => \N__5263\,
            in2 => \N__5224\,
            in3 => \N__6049\,
            lcout => \VPP_VDDQ.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIJCTQ_0_1_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__8393\,
            in1 => \N__5682\,
            in2 => \N__6201\,
            in3 => \N__8237\,
            lcout => \VPP_VDDQ.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVF931_0_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8390\,
            in1 => \N__5965\,
            in2 => \_gnd_net_\,
            in3 => \N__8234\,
            lcout => \VPP_VDDQ.count_2_1_6\,
            ltout => \VPP_VDDQ.count_2_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNID7TR_6_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6768\,
            in2 => \N__5257\,
            in3 => \N__7683\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8391\,
            in1 => \N__5963\,
            in2 => \_gnd_net_\,
            in3 => \N__8236\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8754\,
            ce => \N__7684\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8235\,
            in1 => \N__5747\,
            in2 => \_gnd_net_\,
            in3 => \N__8392\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8754\,
            ce => \N__7684\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8238\,
            in1 => \N__8423\,
            in2 => \N__5929\,
            in3 => \N__7398\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8733\,
            ce => \N__7719\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8421\,
            in1 => \N__8240\,
            in2 => \_gnd_net_\,
            in3 => \N__6048\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8733\,
            ce => \N__7719\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIPT891_12_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5251\,
            in1 => \N__7706\,
            in2 => \_gnd_net_\,
            in3 => \N__6004\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => \VPP_VDDQ.count_2Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8239\,
            in1 => \N__8422\,
            in2 => \N__5254\,
            in3 => \N__6016\,
            lcout => \VPP_VDDQ.count_2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8733\,
            ce => \N__7719\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIE8TR_7_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6698\,
            in1 => \N__7705\,
            in2 => \_gnd_net_\,
            in3 => \N__6027\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_15_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6829\,
            in1 => \N__6914\,
            in2 => \N__6961\,
            in3 => \N__6889\,
            lcout => \VPP_VDDQ.N_1_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8227\,
            in1 => \N__8420\,
            in2 => \N__7409\,
            in3 => \N__5925\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINQ791_11_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__7707\,
            in1 => \_gnd_net_\,
            in2 => \N__5368\,
            in3 => \N__5365\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6174\,
            in2 => \N__5650\,
            in3 => \N__5359\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5353\,
            in1 => \N__5346\,
            in2 => \_gnd_net_\,
            in3 => \N__6175\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5345\,
            in1 => \N__5330\,
            in2 => \N__5283\,
            in3 => \N__5311\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__5312\,
            in1 => \_gnd_net_\,
            in2 => \N__5616\,
            in3 => \N__6177\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6173\,
            in2 => \N__5284\,
            in3 => \N__5293\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__5645\,
            in1 => \N__5585\,
            in2 => \N__5632\,
            in3 => \N__5609\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__5596\,
            in1 => \_gnd_net_\,
            in2 => \N__5590\,
            in3 => \N__6176\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5571\,
            in1 => \N__5559\,
            in2 => \N__5548\,
            in3 => \N__5532\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5520\,
            in1 => \N__5508\,
            in2 => \N__5497\,
            in3 => \N__5481\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5469\,
            in1 => \N__5457\,
            in2 => \N__5446\,
            in3 => \N__5430\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5418\,
            in1 => \N__5406\,
            in2 => \N__5395\,
            in3 => \N__5379\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNINUSC_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__6476\,
            in1 => \N__6417\,
            in2 => \N__6379\,
            in3 => \N__6555\,
            lcout => \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI82TR_0_1_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__5775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7505\,
            lcout => \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5731\,
            in1 => \N__5659\,
            in2 => \N__5692\,
            in3 => \N__6031\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNILHSU_0_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111111111"
        )
    port map (
            in0 => \N__5722\,
            in1 => \N__7639\,
            in2 => \N__5716\,
            in3 => \N__6844\,
            lcout => \VPP_VDDQ.m4_1\,
            ltout => \VPP_VDDQ.m4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5713\,
            in3 => \N__8108\,
            lcout => \VPP_VDDQ.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__8110\,
            in1 => \_gnd_net_\,
            in2 => \N__8394\,
            in3 => \N__5705\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8774\,
            ce => \N__7640\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI82TR_1_1_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5706\,
            in1 => \N__8336\,
            in2 => \_gnd_net_\,
            in3 => \N__8109\,
            lcout => \VPP_VDDQ.count_2_1_1\,
            ltout => \VPP_VDDQ.count_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI82TR_1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__5673\,
            in1 => \N__6172\,
            in2 => \N__5662\,
            in3 => \N__6723\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIR9731_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5752\,
            in1 => \N__8335\,
            in2 => \_gnd_net_\,
            in3 => \N__8152\,
            lcout => \VPP_VDDQ.count_2_1_4\,
            ltout => \VPP_VDDQ.count_2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIB5TR_4_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6743\,
            in2 => \N__5653\,
            in3 => \N__7682\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6550\,
            in2 => \_gnd_net_\,
            in3 => \N__6415\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_en_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIJCTQ_1_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__6486\,
            in1 => \N__6181\,
            in2 => \N__5905\,
            in3 => \N__6374\,
            lcout => \VPP_VDDQ.count_2_en\,
            ltout => \VPP_VDDQ.count_2_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIN3531_2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6100\,
            in2 => \N__5902\,
            in3 => \N__8056\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5898\,
            in1 => \N__5886\,
            in2 => \N__5875\,
            in3 => \N__5859\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5847\,
            in1 => \N__5835\,
            in2 => \N__5824\,
            in3 => \N__5808\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNI8PF7_1_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__6416\,
            in1 => \_gnd_net_\,
            in2 => \N__6567\,
            in3 => \N__8222\,
            lcout => \VPP_VDDQ.un1_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5779\,
            in2 => \N__7507\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8478\,
            in2 => \_gnd_net_\,
            in3 => \N__5764\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7579\,
            in2 => \_gnd_net_\,
            in3 => \N__5761\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIR9731_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5758\,
            in2 => \_gnd_net_\,
            in3 => \N__5734\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIRZ0Z9731\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7320\,
            in2 => \_gnd_net_\,
            in3 => \N__5974\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVF931_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5971\,
            in2 => \_gnd_net_\,
            in3 => \N__5953\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVFZ0Z931\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JA31_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5950\,
            in3 => \N__5941\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7365\,
            in3 => \N__5938\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_THRU_LUT4_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7450\,
            in3 => \N__5935\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_THRU_LUT4_0_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7538\,
            in3 => \N__5932\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_THRU_LUT4_0_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7408\,
            in3 => \N__5914\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_THRU_LUT4_0_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6913\,
            in2 => \_gnd_net_\,
            in3 => \N__5911\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_THRU_LUT4_0_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6891\,
            in3 => \N__5908\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_THRU_LUT4_0_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6959\,
            in3 => \N__6055\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_THRU_LUT4_0_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6052\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JA31_0_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8226\,
            in1 => \N__8424\,
            in2 => \_gnd_net_\,
            in3 => \N__6047\,
            lcout => \VPP_VDDQ.count_2_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8412\,
            in1 => \N__8228\,
            in2 => \N__6924\,
            in3 => \N__6015\,
            lcout => \VPP_VDDQ.count_2_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8229\,
            in1 => \N__8413\,
            in2 => \N__6892\,
            in3 => \N__5991\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIR0A91_13_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__7708\,
            in1 => \_gnd_net_\,
            in2 => \N__5998\,
            in3 => \N__5983\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => \VPP_VDDQ.count_2Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8231\,
            in1 => \N__8416\,
            in2 => \N__5995\,
            in3 => \N__5992\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8776\,
            ce => \N__7710\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8414\,
            in1 => \N__8230\,
            in2 => \N__6960\,
            in3 => \N__6114\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIT3B91_14_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6106\,
            in2 => \N__5977\,
            in3 => \N__7709\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => \VPP_VDDQ.count_2Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8415\,
            in1 => \N__8233\,
            in2 => \N__6118\,
            in3 => \N__6115\,
            lcout => \VPP_VDDQ.count_2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8776\,
            ce => \N__7710\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8232\,
            in1 => \N__8417\,
            in2 => \N__8449\,
            in3 => \N__8489\,
            lcout => \VPP_VDDQ.count_2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8776\,
            ce => \N__7710\,
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6091\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6085\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6079\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6073\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6067\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6061\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6343\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6331\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6322\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6319\,
            in1 => \N__6279\,
            in2 => \N__6252\,
            in3 => \N__6225\,
            lcout => rsmrst_pwrgd_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.G_76_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__6474\,
            in1 => \_gnd_net_\,
            in2 => \N__6187\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.GZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.G_10_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6167\,
            in2 => \_gnd_net_\,
            in3 => \N__6473\,
            lcout => \G_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6171\,
            in2 => \_gnd_net_\,
            in3 => \N__6475\,
            lcout => \clk_100Khz_signalkeep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010100000"
        )
    port map (
            in0 => \N__7255\,
            in1 => \N__6547\,
            in2 => \N__6378\,
            in3 => \N__6621\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8748\,
            ce => \N__6591\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000100000"
        )
    port map (
            in0 => \N__6548\,
            in1 => \N__6369\,
            in2 => \N__6625\,
            in3 => \N__7254\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.m4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNISBBC7_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__6469\,
            in1 => \_gnd_net_\,
            in2 => \N__6634\,
            in3 => \N__6631\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6613\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__6373\,
            in1 => \N__8354\,
            in2 => \N__6610\,
            in3 => \N__6549\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.m6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIIOCG_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6601\,
            in2 => \N__6607\,
            in3 => \N__6468\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__6554\,
            in1 => \N__8353\,
            in2 => \N__6604\,
            in3 => \N__6422\,
            lcout => \VPP_VDDQ.curr_state_2_e_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8748\,
            ce => \N__6591\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__6978\,
            in1 => \N__8340\,
            in2 => \N__7580\,
            in3 => \N__8201\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIP6631_3_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6967\,
            in2 => \N__6577\,
            in3 => \N__7700\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNO_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__6418\,
            in1 => \N__6546\,
            in2 => \N__6487\,
            in3 => \N__8200\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNI_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6423\,
            in3 => \N__6368\,
            lcout => \VPP_VDDQ.un5_clk_100khz\,
            ltout => \VPP_VDDQ.un5_clk_100khz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__6654\,
            in1 => \N__8341\,
            in2 => \N__6781\,
            in3 => \N__7322\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNITC831_5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__6640\,
            in1 => \_gnd_net_\,
            in2 => \N__6778\,
            in3 => \N__7702\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIIJV1_4_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6775\,
            in2 => \_gnd_net_\,
            in3 => \N__6751\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNILHSU_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6724\,
            in1 => \N__6706\,
            in2 => \N__6679\,
            in3 => \N__7701\,
            lcout => \VPP_VDDQ.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8384\,
            in1 => \N__8217\,
            in2 => \N__6825\,
            in3 => \N__6798\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__7360\,
            in1 => \N__8205\,
            in2 => \N__8409\,
            in3 => \N__6672\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI3MB31_8_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__6661\,
            in1 => \_gnd_net_\,
            in2 => \N__6676\,
            in3 => \N__7681\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => \VPP_VDDQ.count_2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__8218\,
            in1 => \N__6673\,
            in2 => \N__6664\,
            in3 => \N__8385\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => \N__7704\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8358\,
            in1 => \N__8207\,
            in2 => \N__6655\,
            in3 => \N__7321\,
            lcout => \VPP_VDDQ.count_2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => \N__7704\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__8206\,
            in1 => \N__7569\,
            in2 => \N__6982\,
            in3 => \N__8359\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => \N__7704\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__7451\,
            in1 => \N__7036\,
            in2 => \N__8245\,
            in3 => \N__8386\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => \N__7704\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_15_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6958\,
            in1 => \N__6818\,
            in2 => \N__6928\,
            in3 => \N__6890\,
            lcout => \VPP_VDDQ.g0_2_a2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_10_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7416\,
            in1 => \N__6862\,
            in2 => \N__7539\,
            in3 => \N__7452\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_14_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7361\,
            in1 => \N__7582\,
            in2 => \N__6850\,
            in3 => \N__7327\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_RNIZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_2_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8488\,
            in2 => \N__6847\,
            in3 => \N__7506\,
            lcout => \VPP_VDDQ.count_2_RNI_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIV6C91_15_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6787\,
            in1 => \N__7703\,
            in2 => \_gnd_net_\,
            in3 => \N__6835\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => \VPP_VDDQ.count_2Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__8224\,
            in1 => \N__8419\,
            in2 => \N__6802\,
            in3 => \N__6799\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8773\,
            ce => \N__7720\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__7449\,
            in1 => \N__8410\,
            in2 => \N__8242\,
            in3 => \N__7035\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI5PC31_9_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7024\,
            in2 => \N__7015\,
            in3 => \N__7697\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__7531\,
            in1 => \N__8411\,
            in2 => \N__8243\,
            in3 => \N__7008\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIES131_10_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6997\,
            in2 => \N__7012\,
            in3 => \N__7698\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => \VPP_VDDQ.count_2Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__8418\,
            in1 => \N__7009\,
            in2 => \N__7000\,
            in3 => \N__8223\,
            lcout => \VPP_VDDQ.count_2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => \N__7699\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9098\,
            in1 => \N__7852\,
            in2 => \N__7168\,
            in3 => \N__7167\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9052\,
            in1 => \N__7903\,
            in2 => \_gnd_net_\,
            in3 => \N__6991\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9099\,
            in1 => \N__7930\,
            in2 => \_gnd_net_\,
            in3 => \N__6988\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_3_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9053\,
            in1 => \N__8005\,
            in2 => \_gnd_net_\,
            in3 => \N__6985\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_4_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9100\,
            in1 => \N__7942\,
            in2 => \_gnd_net_\,
            in3 => \N__7063\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_5_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9054\,
            in1 => \N__8032\,
            in2 => \_gnd_net_\,
            in3 => \N__7060\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_6_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9101\,
            in1 => \N__8044\,
            in2 => \_gnd_net_\,
            in3 => \N__7057\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_7_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9055\,
            in1 => \N__8019\,
            in2 => \_gnd_net_\,
            in3 => \N__7054\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__8758\,
            ce => 'H',
            sr => \N__7144\
        );

    \RSMRST_PWRGD.count_8_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9051\,
            in1 => \N__7954\,
            in2 => \_gnd_net_\,
            in3 => \N__7051\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__8619\,
            ce => 'H',
            sr => \N__7139\
        );

    \RSMRST_PWRGD.count_9_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9047\,
            in1 => \N__7917\,
            in2 => \_gnd_net_\,
            in3 => \N__7048\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__8619\,
            ce => 'H',
            sr => \N__7139\
        );

    \RSMRST_PWRGD.count_10_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9048\,
            in1 => \N__7981\,
            in2 => \_gnd_net_\,
            in3 => \N__7045\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__8619\,
            ce => 'H',
            sr => \N__7139\
        );

    \RSMRST_PWRGD.count_11_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9045\,
            in1 => \N__7993\,
            in2 => \_gnd_net_\,
            in3 => \N__7042\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__8619\,
            ce => 'H',
            sr => \N__7139\
        );

    \RSMRST_PWRGD.count_12_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9049\,
            in1 => \N__7968\,
            in2 => \_gnd_net_\,
            in3 => \N__7039\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__8619\,
            ce => 'H',
            sr => \N__7139\
        );

    \RSMRST_PWRGD.count_13_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9046\,
            in1 => \N__7879\,
            in2 => \_gnd_net_\,
            in3 => \N__7240\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__8619\,
            ce => 'H',
            sr => \N__7139\
        );

    \RSMRST_PWRGD.count_14_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9050\,
            in1 => \N__7891\,
            in2 => \_gnd_net_\,
            in3 => \N__7237\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__8619\,
            ce => 'H',
            sr => \N__7139\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7220\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7866\,
            in2 => \_gnd_net_\,
            in3 => \N__7171\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8759\,
            ce => \N__7111\,
            sr => \N__7143\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__9131\,
            in1 => \N__9184\,
            in2 => \_gnd_net_\,
            in3 => \N__8807\,
            lcout => \RSMRST_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNINN7M6_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__9152\,
            in1 => \N__9183\,
            in2 => \N__8815\,
            in3 => \N__9132\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.G_29_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7147\,
            in3 => \N__8905\,
            lcout => \G_29\,
            ltout => \G_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__8906\,
            in1 => \_gnd_net_\,
            in2 => \N__7114\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.N_15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_1_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7077\,
            in1 => \N__9185\,
            in2 => \_gnd_net_\,
            in3 => \N__7768\,
            lcout => \VCCIN_PWRGD.un10_outputZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_RNO_0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9133\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.curr_state10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__9182\,
            in1 => \N__7767\,
            in2 => \N__7816\,
            in3 => \N__8907\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI71TR_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__7717\,
            in1 => \N__7491\,
            in2 => \N__7729\,
            in3 => \N__7741\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8405\,
            in2 => \N__7732\,
            in3 => \N__8241\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8779\,
            ce => \N__7718\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_2_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7581\,
            in2 => \_gnd_net_\,
            in3 => \N__8490\,
            lcout => \VPP_VDDQ.g0_2_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_10_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7543\,
            in1 => \N__7498\,
            in2 => \N__7459\,
            in3 => \N__7417\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.g0_2_a2_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_5_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7369\,
            in1 => \N__7336\,
            in2 => \N__7330\,
            in3 => \N__7326\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.g0_2_a2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIUPFQ6_1_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__7291\,
            in1 => \N__7279\,
            in2 => \N__7267\,
            in3 => \N__7264\,
            lcout => \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__8494\,
            in1 => \N__8448\,
            in2 => \N__8428\,
            in3 => \N__8225\,
            lcout => \VPP_VDDQ.count_2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI9RLK1_3_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8043\,
            in1 => \N__8031\,
            in2 => \N__8020\,
            in3 => \N__8004\,
            lcout => \RSMRST_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIIRGK_10_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7992\,
            in1 => \N__7980\,
            in2 => \N__7969\,
            in3 => \N__7953\,
            lcout => \RSMRST_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI4MLK1_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7941\,
            in1 => \N__7929\,
            in2 => \N__7918\,
            in3 => \N__7902\,
            lcout => \RSMRST_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7890\,
            in1 => \N__7878\,
            in2 => \N__7867\,
            in3 => \N__7851\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un4_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIR8OP4_10_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7840\,
            in1 => \N__7834\,
            in2 => \N__7828\,
            in3 => \N__7825\,
            lcout => \RSMRST_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m3_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9186\,
            in1 => \N__9134\,
            in2 => \_gnd_net_\,
            in3 => \N__9153\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.i3_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000011001100"
        )
    port map (
            in0 => \N__8813\,
            in1 => \N__9135\,
            in2 => \N__7819\,
            in3 => \N__8979\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9253\,
            in1 => \N__9241\,
            in2 => \N__9226\,
            in3 => \N__9208\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m5_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__9187\,
            in1 => \N__8812\,
            in2 => \_gnd_net_\,
            in3 => \N__9154\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__8814\,
            in1 => \N__9136\,
            in2 => \N__9109\,
            in3 => \N__8980\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8788\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
