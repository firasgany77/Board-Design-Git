-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 13 2022 11:36:22

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : in std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__33702\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \VCCG0\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9\ : std_logic;
signal \PCH_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_5\ : std_logic;
signal \PCH_PWRGD.count_rst_11_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_4_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.count_rst_10\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \PCH_PWRGD.count_rst_10_cascade_\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \PCH_PWRGD.count_rst_12\ : std_logic;
signal \PCH_PWRGD.count_0_2\ : std_logic;
signal \PCH_PWRGD.count_0_14\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.count_0_6\ : std_logic;
signal \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1_cascade_\ : std_logic;
signal \PCH_PWRGD.N_2284_i_cascade_\ : std_logic;
signal \PCH_PWRGD.N_655_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1\ : std_logic;
signal \PCH_PWRGD.count_0_1\ : std_logic;
signal \PCH_PWRGD.count_rst_13\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.N_2284_i\ : std_logic;
signal \POWERLED.count_0_2\ : std_logic;
signal \G_12\ : std_logic;
signal \POWERLED.count_0_11\ : std_logic;
signal \POWERLED.count_0_3\ : std_logic;
signal \POWERLED.count_0_0\ : std_logic;
signal \POWERLED.count_1_0_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_1_1_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_0_1\ : std_logic;
signal \POWERLED.count_0_4\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \POWERLED.count_1_2\ : std_logic;
signal \POWERLED.un1_count_cry_1\ : std_logic;
signal \POWERLED.count_1_3\ : std_logic;
signal \POWERLED.un1_count_cry_2_cZ0\ : std_logic;
signal \POWERLED.count_1_4\ : std_logic;
signal \POWERLED.un1_count_cry_3_cZ0\ : std_logic;
signal \POWERLED.un1_count_cry_4_cZ0\ : std_logic;
signal \POWERLED.un1_count_cry_5\ : std_logic;
signal \POWERLED.un1_count_cry_6\ : std_logic;
signal \POWERLED.un1_count_cry_7\ : std_logic;
signal \POWERLED.un1_count_cry_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \POWERLED.un1_count_cry_9\ : std_logic;
signal \POWERLED.count_1_11\ : std_logic;
signal \POWERLED.un1_count_cry_10\ : std_logic;
signal \POWERLED.un1_count_cry_11\ : std_logic;
signal \POWERLED.un1_count_cry_12\ : std_logic;
signal \POWERLED.un1_count_cry_13\ : std_logic;
signal \POWERLED.un1_count_cry_14\ : std_logic;
signal \POWERLED.count_1_12\ : std_logic;
signal \POWERLED.count_0_12\ : std_logic;
signal \POWERLED.N_437_cascade_\ : std_logic;
signal \POWERLED.N_2305_i_cascade_\ : std_logic;
signal \POWERLED.N_660_cascade_\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i\ : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa_0\ : std_logic;
signal \POWERLED.pwm_out_en_cascade_\ : std_logic;
signal \POWERLED.pwm_outZ0\ : std_logic;
signal pwrbtn_led : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_2_1_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.count_0_12\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \PCH_PWRGD.N_386_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \PCH_PWRGD.count_rst_3_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_7_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_14_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_7\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_6_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_4_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_5_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_3_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_12_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_12_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_1_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_0_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_2_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_11_0\ : std_logic;
signal \PCH_PWRGD.count_rst\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \PCH_PWRGD.count_rst_1\ : std_logic;
signal \PCH_PWRGD.count_0_13\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.count_0_10\ : std_logic;
signal \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \PCH_PWRGD.N_2266_i_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1\ : std_logic;
signal \PCH_PWRGD.m6_i_i_a2_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_7_0\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_655\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.N_386\ : std_logic;
signal \PCH_PWRGD.curr_state_0_sqmuxa_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_0_0\ : std_logic;
signal \VPP_VDDQ.N_53_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.m4_0_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_60_cascade_\ : std_logic;
signal \VPP_VDDQ.N_60_i\ : std_logic;
signal \VPP_VDDQ.N_60\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_ok_cascade_\ : std_logic;
signal vccst_pwrgd : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_\ : std_logic;
signal pch_pwrok : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa\ : std_logic;
signal \POWERLED.un79_clk_100khzlt6\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_4\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khz\ : std_logic;
signal \POWERLED.un79_clk_100khz_cascade_\ : std_logic;
signal \POWERLED.g0_2_1\ : std_logic;
signal \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0\ : std_logic;
signal \POWERLED.count_0_15\ : std_logic;
signal \POWERLED.count_1_7\ : std_logic;
signal \POWERLED.count_0_7\ : std_logic;
signal \POWERLED.count_1_8\ : std_logic;
signal \POWERLED.count_0_8\ : std_logic;
signal \POWERLED.count_1_9\ : std_logic;
signal \POWERLED.count_0_9\ : std_logic;
signal \POWERLED.count_1_13\ : std_logic;
signal \POWERLED.count_0_13\ : std_logic;
signal \POWERLED.count_1_5\ : std_logic;
signal \POWERLED.count_0_5\ : std_logic;
signal \POWERLED.count_1_14\ : std_logic;
signal \POWERLED.count_0_14\ : std_logic;
signal \POWERLED.count_1_6\ : std_logic;
signal \POWERLED.count_0_6\ : std_logic;
signal \POWERLED.count_1_10\ : std_logic;
signal \POWERLED.count_0_10\ : std_logic;
signal v33a_enn : std_logic;
signal \HDA_STRAP.N_16_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_okZ0_cascade_\ : std_logic;
signal \N_428_cascade_\ : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \HDA_STRAP.m14_i_0_cascade_\ : std_logic;
signal \N_428\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal \HDA_STRAP.HDA_SDO_ATP_3_0\ : std_logic;
signal \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \PCH_PWRGD.N_670\ : std_logic;
signal \PCH_PWRGD.N_2266_i\ : std_logic;
signal \PCH_PWRGD.N_38_f0\ : std_logic;
signal \PCH_PWRGD.curr_state_0_sqmuxa\ : std_logic;
signal \PCH_PWRGD.N_38_f0_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_sqmuxa_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \VPP_VDDQ.count_2_1_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_1_cascade_\ : std_logic;
signal slp_susn : std_logic;
signal v5a_ok : std_logic;
signal v33a_ok : std_logic;
signal v1p8a_ok : std_logic;
signal \rsmrst_pwrgd_signal_cascade_\ : std_logic;
signal \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_264_i\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_1\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_13_cascade_\ : std_logic;
signal \VPP_VDDQ.N_1_i\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.N_1_i_cascade_\ : std_logic;
signal \VPP_VDDQ.N_664\ : std_logic;
signal \N_639\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_7\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_10\ : std_logic;
signal \VPP_VDDQ.count_2_0_12\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.count_2_0_14\ : std_logic;
signal \POWERLED.N_2305_i\ : std_logic;
signal \POWERLED.N_660\ : std_logic;
signal \POWERLED.curr_state_1_0\ : std_logic;
signal \N_557_g\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_4_l_fx\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_7_l_fx\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.un1_count_cry_0_i\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.N_5036_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_0\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.N_5037_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.N_5038_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.N_5039_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_3\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.N_5040_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_4\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.N_5041_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_8\ : std_logic;
signal \POWERLED.N_5042_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_8\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.N_5043_i\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \POWERLED.N_5044_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_8\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_8\ : std_logic;
signal \POWERLED.N_5045_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.N_5046_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.N_5047_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_11\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.N_5048_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.N_5049_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_13\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.N_5050_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_14\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_8\ : std_logic;
signal \bfn_5_1_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_0\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7_THRU_CO\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_8\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_16\ : std_logic;
signal \RSMRST_PWRGD.N_92_1\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \VPP_VDDQ.count_2_0_5\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.count_2_0_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.count_2_1_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.count_2_1_9\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.count_2_1_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.count_2_1_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.count_2_1_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.count_2_1_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.count_2_1_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.count_2_1_sqmuxa\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2_c\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_c\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_c\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_c\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_c\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8_cascade_\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2150\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_0\ : std_logic;
signal \POWERLED.un85_clk_100khz_2\ : std_logic;
signal \POWERLED.un85_clk_100khz_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_1\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_8\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_8\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_8\ : std_logic;
signal \HDA_STRAP.countZ0Z_8\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \HDA_STRAP.countZ0Z_15\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.countZ0Z_3\ : std_logic;
signal \HDA_STRAP.countZ0Z_5\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.un4_count_12\ : std_logic;
signal \HDA_STRAP.un4_count_13_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_10\ : std_logic;
signal \HDA_STRAP.countZ0Z_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.countZ0Z_13\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.un4_count_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_1\ : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \HDA_STRAP.un4_count_9\ : std_logic;
signal \HDA_STRAP.un4_count\ : std_logic;
signal \HDA_STRAP.curr_state_RNIH91AZ0Z_0\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15_THRU_CO\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_6\ : std_logic;
signal \VPP_VDDQ.count_2_0_4\ : std_logic;
signal \VPP_VDDQ.count_2_1_4\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_6\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_0\ : std_logic;
signal \VPP_VDDQ.count_2_0_2\ : std_logic;
signal \VPP_VDDQ.count_2_1_2\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_9\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_8\ : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8_cascade_\ : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \bfn_6_16_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.count_off_0_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.count_off_0_10\ : std_logic;
signal \POWERLED.count_off_0_11\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1_cZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_off_1_9\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_off_1_10\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_off_1_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14\ : std_logic;
signal \POWERLED.count_off_1_12\ : std_logic;
signal \POWERLED.count_off_0_12\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \N_555\ : std_logic;
signal \G_14\ : std_logic;
signal \N_662\ : std_logic;
signal \RSMRST_PWRGD_curr_state_0\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \VCCST_EN_i_1_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_5_cascade_\ : std_logic;
signal \POWERLED.N_432\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_7_2\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_0_1_1_cascade_\ : std_logic;
signal \POWERLED.N_423\ : std_logic;
signal \POWERLED.N_671\ : std_logic;
signal \POWERLED.func_state_enZ0\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.N_512_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_39_and_i_1_cascade_\ : std_logic;
signal \POWERLED.N_514\ : std_logic;
signal \POWERLED.N_508\ : std_logic;
signal \POWERLED.un1_clk_100khz_33_and_i_1_cascade_\ : std_logic;
signal \POWERLED.count_off_1_7\ : std_logic;
signal \POWERLED.count_off_0_7\ : std_logic;
signal \POWERLED.count_off_1_8\ : std_logic;
signal \POWERLED.count_off_0_8\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_28\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_0\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_1\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_11\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_14\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_15\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.N_598_cascade_\ : std_logic;
signal \POWERLED.N_450_cascade_\ : std_logic;
signal \POWERLED.N_599\ : std_logic;
signal \POWERLED.N_449_cascade_\ : std_logic;
signal \POWERLED.N_2376_i\ : std_logic;
signal \POWERLED.N_2376_i_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_0_5\ : std_logic;
signal \POWERLED.count_off_1_5\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.count_offZ0Z_5_cascade_\ : std_logic;
signal \POWERLED.count_off_0_0\ : std_logic;
signal \POWERLED.count_off_1_0\ : std_logic;
signal \POWERLED.count_off_0_2\ : std_logic;
signal \POWERLED.count_off_1_2\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.count_off_1_13\ : std_logic;
signal \POWERLED.count_off_0_13\ : std_logic;
signal \POWERLED.count_off_1_14\ : std_logic;
signal \POWERLED.count_off_0_14\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14_c_RNIPGZ0Z497\ : std_logic;
signal \POWERLED.count_off_0_15\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_offZ0Z_15_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.count_off_0_6\ : std_logic;
signal \POWERLED.count_off_1_6\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \POWERLED.N_673_0_cascade_\ : std_logic;
signal \POWERLED.N_423_0\ : std_logic;
signal \v5s_enn_cascade_\ : std_logic;
signal \POWERLED.func_state_en_0_0\ : std_logic;
signal \POWERLED.func_stateZ1Z_0\ : std_logic;
signal \POWERLED.func_state_en_0_0_cascade_\ : std_logic;
signal \RSMRSTn_fast\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_0_2\ : std_logic;
signal \POWERLED.func_state_RNI5SKJ1Z0Z_1\ : std_logic;
signal vddq_ok : std_logic;
signal \func_state_RNI_2_0_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m0_1_1\ : std_logic;
signal \POWERLED.N_540_1\ : std_logic;
signal \POWERLED.N_542\ : std_logic;
signal \POWERLED.N_673\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_0_1_cascade_\ : std_logic;
signal \POWERLED.N_6_1\ : std_logic;
signal \POWERLED.N_74_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_ns_1_1\ : std_logic;
signal \POWERLED.func_state_1_m2_1\ : std_logic;
signal \POWERLED.func_state_RNIBVNSZ0Z_0\ : std_logic;
signal \POWERLED.N_6_2\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_a2_0_1_2\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_0_2_cascade_\ : std_logic;
signal \POWERLED.N_71_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.N_426_i_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_1\ : std_logic;
signal \POWERLED.N_71\ : std_logic;
signal \POWERLED.dutycycle_eena_1_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_2\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_29\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\ : std_logic;
signal \POWERLED.mult1_un47_sum_axb_4\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.dutycycle_en_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_41_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_40_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_a4_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_a5_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_a0_2\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_12\ : std_logic;
signal \POWERLED.dutycycleZ1Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNI_12Z0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_15\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14_cascade_\ : std_logic;
signal \POWERLED.N_2381_i_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_0_a2_0_5\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ1Z_11\ : std_logic;
signal \POWERLED.dutycycle_en_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_13\ : std_logic;
signal \VPP_VDDQ.un6_count_8_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \VPP_VDDQ.un6_count_9\ : std_logic;
signal \POWERLED.G_30Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ_un6_count\ : std_logic;
signal \G_30_cascade_\ : std_logic;
signal \N_626\ : std_logic;
signal \VPP_VDDQ_curr_state_1\ : std_logic;
signal \VPP_VDDQ_curr_state_0\ : std_logic;
signal \POWERLED.count_off_0_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_offZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.un34_clk_100khz_10\ : std_logic;
signal \POWERLED.un34_clk_100khz_11\ : std_logic;
signal \POWERLED.un34_clk_100khz_8_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_9\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\ : std_logic;
signal \POWERLED.count_off_0_4\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1\ : std_logic;
signal \POWERLED.count_off_0_1\ : std_logic;
signal \POWERLED.func_state_RNI7LSV8Z0Z_0\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \N_7_cascade_\ : std_logic;
signal \N_8_0_cascade_\ : std_logic;
signal \POWERLED.g0_5Z0Z_1_cascade_\ : std_logic;
signal \POWERLED_g2_1_0_0\ : std_logic;
signal \POWERLED.N_74\ : std_logic;
signal \POWERLED.N_4_0_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_0_0_0\ : std_logic;
signal \POWERLED.g1_0_0\ : std_logic;
signal \POWERLED.func_state_1_m2_N_3_7_1\ : std_logic;
signal \clk_100Khz_signalkeep_3_fast\ : std_logic;
signal \POWERLED.N_671_0\ : std_logic;
signal \G_7_i_a4_1_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.G_7_i_0\ : std_logic;
signal \POWERLED.N_533_cascade_\ : std_logic;
signal \POWERLED.N_533\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_3_0_sx\ : std_logic;
signal \POWERLED.un1_dutycycle_164_0_a3_0_a2_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_4\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_9_0\ : std_logic;
signal \POWERLED.count_clk_0_7\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m3\ : std_logic;
signal \POWERLED.un1_clk_100khz_52_and_i_0_m2_ns_1_cascade_\ : std_logic;
signal \POWERLED.N_448_cascade_\ : std_logic;
signal \POWERLED.N_656_0\ : std_logic;
signal \POWERLED.N_133_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m4\ : std_logic;
signal \POWERLED.dutycycle_eena_14_c\ : std_logic;
signal \POWERLED.N_488_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m2\ : std_logic;
signal \POWERLED.un1_clk_100khz_30_and_i_0_0_sx_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_0_a2_1_0\ : std_logic;
signal \POWERLED.un1_dutycycle_96_0_a3_0_a2_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_3\ : std_logic;
signal \POWERLED.N_251_cascade_\ : std_logic;
signal \POWERLED.N_506\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_cZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12\ : std_logic;
signal \POWERLED.N_435_i\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\ : std_logic;
signal vccst_en : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\ : std_logic;
signal \POWERLED.dutycycle_RNIP1UTZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIF86R3Z0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNIP1UTZ0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNIF86R3Z0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_4\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_0_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_11\ : std_logic;
signal \POWERLED.dutycycleZ1Z_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\ : std_logic;
signal \POWERLED.dutycycle_RNIRT5H5Z0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_10_8_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_4\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_4_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_4_1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_a0_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_4\ : std_logic;
signal \POWERLED.un1_dutycycle_53_40_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_11_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_11_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_45_0\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_4\ : std_logic;
signal \POWERLED.un1_dutycycle_53_35_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_22\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_10_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_35_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_a0_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_a0_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_a0_0_0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\ : std_logic;
signal \POWERLED.dutycycle_en_4\ : std_logic;
signal \POWERLED.dutycycleZ1Z_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_0_a2_0_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_0_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_2_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_a1_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_3_0\ : std_logic;
signal \VPP_VDDQ.N_64_i\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \N_92_g\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.N_92_0\ : std_logic;
signal \G_30\ : std_logic;
signal \POWERLED.count_clk_0_4\ : std_logic;
signal \POWERLED.count_clk_0_5\ : std_logic;
signal \POWERLED.count_clk_0_6\ : std_logic;
signal \clk_100Khz_signalkeep_3\ : std_logic;
signal \clk_100Khz_signalkeep_3_rep1\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_1\ : std_logic;
signal \POWERLED.count_clk_0_11\ : std_logic;
signal \POWERLED.count_off_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3_cascade_\ : std_logic;
signal \POWERLED.N_668_cascade_\ : std_logic;
signal \POWERLED.N_490\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_\ : std_logic;
signal \POWERLED.N_123\ : std_logic;
signal \POWERLED.N_443\ : std_logic;
signal \POWERLED.count_off_RNIH9TEZ0Z_10\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_0_2_1\ : std_logic;
signal \POWERLED.N_668\ : std_logic;
signal \POWERLED.count_off_1_sqmuxa\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m0\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1\ : std_logic;
signal \POWERLED.func_state_RNI_3Z0Z_1\ : std_logic;
signal \N_247\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_2\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_1_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_4\ : std_logic;
signal \POWERLED.func_state_RNI_0Z0Z_1\ : std_logic;
signal \func_state_RNI_4_1\ : std_logic;
signal \func_state_RNI_0_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_N_3_mux_0\ : std_logic;
signal \POWERLED.N_546_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_0\ : std_logic;
signal \POWERLED.N_482\ : std_logic;
signal \POWERLED.g0_i_m2_rn_1_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_0_0\ : std_logic;
signal \POWERLED.g0_1\ : std_logic;
signal \POWERLED.dutycycle_eena_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_cascade_\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \POWERLED.g0_i_m2_sn\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.g0_i_m2_rn_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_1\ : std_logic;
signal \POWERLED.dutycycle_1_0_0\ : std_logic;
signal \POWERLED.dutycycle_eena\ : std_logic;
signal \POWERLED.dutycycleZ1Z_0\ : std_logic;
signal \POWERLED.N_510\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_a2_c_cascade_\ : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_a2_d\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_0_2\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_5\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.N_249_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_0_3_1\ : std_logic;
signal \POWERLED.N_203_cascade_\ : std_logic;
signal \POWERLED.N_521_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_43_and_i_1_cascade_\ : std_logic;
signal \POWERLED.N_523\ : std_logic;
signal \POWERLED.N_503_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.un1_clk_100khz_30_and_i_0_a2_5_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_2_0_0_tz_1\ : std_logic;
signal \POWERLED.dutycycle_eena_2_d_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIRUFD6Z0Z_9\ : std_logic;
signal \POWERLED.func_state_RNI2MQDZ0Z_1\ : std_logic;
signal \RSMRSTn_rep1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6\ : std_logic;
signal \POWERLED.N_520_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIRUFD6Z0Z_12\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.N_518_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_42_and_i_1\ : std_logic;
signal \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_d\ : std_logic;
signal \POWERLED.N_526_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI36306Z0Z_14\ : std_logic;
signal \POWERLED.func_state_RNI_8Z0Z_1\ : std_logic;
signal \POWERLED.N_203\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.N_524_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_47_and_i_1\ : std_logic;
signal rsmrstn : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.N_2381_i\ : std_logic;
signal \POWERLED.N_91_1_N\ : std_logic;
signal \POWERLED.N_527_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_48_and_i_1_cascade_\ : std_logic;
signal \POWERLED.N_529\ : std_logic;
signal \POWERLED.dutycycle_en_12\ : std_logic;
signal \POWERLED.count_clk_0_8\ : std_logic;
signal \POWERLED.count_clk_0_9\ : std_logic;
signal \POWERLED.count_clk_0_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_3\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_\ : std_logic;
signal \POWERLED.N_625\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_1\ : std_logic;
signal \POWERLED.N_625_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNIPGQN2_5Z0Z_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13_cZ0\ : std_logic;
signal \POWERLED.func_state_RNI2VV9A_0_0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14\ : std_logic;
signal \POWERLED.count_clk_0_15\ : std_logic;
signal \POWERLED.count_clk_1_15\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_axb_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_axb_14\ : std_logic;
signal \POWERLED.count_clk_0_0\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.count_clk_1_14\ : std_logic;
signal \POWERLED.count_clkZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_1_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_2\ : std_logic;
signal \POWERLED.count_clk_RNISLCE7Z0Z_10\ : std_logic;
signal \POWERLED.count_clk_en_917_0\ : std_logic;
signal \POWERLED.func_state_RNIBVNS_2Z0Z_0\ : std_logic;
signal \POWERLED.count_clk_en_1_cascade_\ : std_logic;
signal \POWERLED.N_617\ : std_logic;
signal \POWERLED.count_clk_en_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_axb_12\ : std_logic;
signal \POWERLED.count_clk_1_13\ : std_logic;
signal \POWERLED.count_clk_0_13\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\ : std_logic;
signal \POWERLED.count_clk_en\ : std_logic;
signal \POWERLED.count_clkZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_0\ : std_logic;
signal \POWERLED.N_676\ : std_logic;
signal \POWERLED.N_492\ : std_logic;
signal \POWERLED.dutycycle_0_5\ : std_logic;
signal \POWERLED.func_state_RNIS28SBZ0Z_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_a2_0_cascade_\ : std_logic;
signal \func_state_RNI_2_0\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_ns_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.N_251\ : std_logic;
signal \POWERLED.N_633\ : std_logic;
signal \POWERLED.func_state_RNIOGRSZ0Z_1_cascade_\ : std_logic;
signal v5s_enn : std_logic;
signal \POWERLED.N_413_N\ : std_logic;
signal \POWERLED.dutycycle_0_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.N_612\ : std_logic;
signal \POWERLED.N_672\ : std_logic;
signal \POWERLED.N_672_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_168_0\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_0\ : std_logic;
signal \POWERLED.N_412_i_cascade_\ : std_logic;
signal \POWERLED.N_604\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_3\ : std_logic;
signal \POWERLED.N_435\ : std_logic;
signal \POWERLED.N_412_i\ : std_logic;
signal \POWERLED.func_state_RNI_5Z0Z_1\ : std_logic;
signal \POWERLED.func_state_RNI_5Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_23_i\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\ : std_logic;
signal \POWERLED.N_85\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_5\ : std_logic;
signal \POWERLED.func_state_RNI12ASZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_613\ : std_logic;
signal slp_s4n : std_logic;
signal \POWERLED.func_state_RNI8AQHZ0Z_0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\ : std_logic;
signal \POWERLED.func_state_RNI12ASZ0Z_1\ : std_logic;
signal \POWERLED.N_83\ : std_logic;
signal slp_s3n : std_logic;
signal \func_state_RNIMJ6IF_0_1\ : std_logic;
signal \RSMRSTn_rep2\ : std_logic;
signal \POWERLED.N_531\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_3_0\ : std_logic;
signal \POWERLED.N_532_cascade_\ : std_logic;
signal \POWERLED.N_530\ : std_logic;
signal \POWERLED.dutycycle_eena_13_c_1\ : std_logic;
signal \POWERLED.N_430\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_3_cascade_\ : std_logic;
signal \G_141\ : std_logic;
signal \POWERLED.dutycycle_RNI0DF58Z0Z_5\ : std_logic;
signal fpga_osc : std_logic;
signal \POWERLED.N_430_iZ0\ : std_logic;
signal \POWERLED.dutycycle_en_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\ : std_logic;
signal \POWERLED.dutycycleZ1Z_3\ : std_logic;
signal \POWERLED.N_421\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_3_1_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5\ : std_logic;
signal \POWERLED.un1_i3_mux_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.d_i3_mux\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VCCST_EN_i_1\ : std_logic;
signal vpp_en : std_logic;
signal vccst_cpu_ok : std_logic;
signal v5s_ok : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_1\ : std_logic;
signal v33s_ok : std_logic;
signal vccin_en : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_2\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    \SUSWARN_N_wire\ <= SUSWARN_N;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33702\,
            DIN => \N__33701\,
            DOUT => \N__33700\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33702\,
            PADOUT => \N__33701\,
            PADIN => \N__33700\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33693\,
            DIN => \N__33692\,
            DOUT => \N__33691\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33693\,
            PADOUT => \N__33692\,
            PADIN => \N__33691\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15680\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33684\,
            DIN => \N__33683\,
            DOUT => \N__33682\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33684\,
            PADOUT => \N__33683\,
            PADIN => \N__33682\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16225\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33675\,
            DIN => \N__33674\,
            DOUT => \N__33673\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33675\,
            PADOUT => \N__33674\,
            PADIN => \N__33673\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14081\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33666\,
            DIN => \N__33665\,
            DOUT => \N__33664\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33666\,
            PADOUT => \N__33665\,
            PADIN => \N__33664\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33657\,
            DIN => \N__33656\,
            DOUT => \N__33655\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33657\,
            PADOUT => \N__33656\,
            PADIN => \N__33655\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33648\,
            DIN => \N__33647\,
            DOUT => \N__33646\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33648\,
            PADOUT => \N__33647\,
            PADIN => \N__33646\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33639\,
            DIN => \N__33638\,
            DOUT => \N__33637\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33639\,
            PADOUT => \N__33638\,
            PADIN => \N__33637\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33630\,
            DIN => \N__33629\,
            DOUT => \N__33628\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33630\,
            PADOUT => \N__33629\,
            PADIN => \N__33628\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29626\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33621\,
            DIN => \N__33620\,
            DOUT => \N__33619\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33621\,
            PADOUT => \N__33620\,
            PADIN => \N__33619\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33612\,
            DIN => \N__33611\,
            DOUT => \N__33610\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33612\,
            PADOUT => \N__33611\,
            PADIN => \N__33610\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33603\,
            DIN => \N__33602\,
            DOUT => \N__33601\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33603\,
            PADOUT => \N__33602\,
            PADIN => \N__33601\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14102\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33594\,
            DIN => \N__33593\,
            DOUT => \N__33592\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33594\,
            PADOUT => \N__33593\,
            PADIN => \N__33592\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33585\,
            DIN => \N__33584\,
            DOUT => \N__33583\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33585\,
            PADOUT => \N__33584\,
            PADIN => \N__33583\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33576\,
            DIN => \N__33575\,
            DOUT => \N__33574\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33576\,
            PADOUT => \N__33575\,
            PADIN => \N__33574\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33567\,
            DIN => \N__33566\,
            DOUT => \N__33565\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33567\,
            PADOUT => \N__33566\,
            PADIN => \N__33565\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33558\,
            DIN => \N__33557\,
            DOUT => \N__33556\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33558\,
            PADOUT => \N__33557\,
            PADIN => \N__33556\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23918\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33549\,
            DIN => \N__33548\,
            DOUT => \N__33547\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33549\,
            PADOUT => \N__33548\,
            PADIN => \N__33547\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33540\,
            DIN => \N__33539\,
            DOUT => \N__33538\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33540\,
            PADOUT => \N__33539\,
            PADIN => \N__33538\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33531\,
            DIN => \N__33530\,
            DOUT => \N__33529\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33531\,
            PADOUT => \N__33530\,
            PADIN => \N__33529\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33522\,
            DIN => \N__33521\,
            DOUT => \N__33520\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33522\,
            PADOUT => \N__33521\,
            PADIN => \N__33520\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33513\,
            DIN => \N__33512\,
            DOUT => \N__33511\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33513\,
            PADOUT => \N__33512\,
            PADIN => \N__33511\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33504\,
            DIN => \N__33503\,
            DOUT => \N__33502\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33504\,
            PADOUT => \N__33503\,
            PADIN => \N__33502\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33495\,
            DIN => \N__33494\,
            DOUT => \N__33493\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33495\,
            PADOUT => \N__33494\,
            PADIN => \N__33493\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33486\,
            DIN => \N__33485\,
            DOUT => \N__33484\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33486\,
            PADOUT => \N__33485\,
            PADIN => \N__33484\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27692\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33477\,
            DIN => \N__33476\,
            DOUT => \N__33475\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33477\,
            PADOUT => \N__33476\,
            PADIN => \N__33475\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33468\,
            DIN => \N__33467\,
            DOUT => \N__33466\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33468\,
            PADOUT => \N__33467\,
            PADIN => \N__33466\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15461\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33459\,
            DIN => \N__33458\,
            DOUT => \N__33457\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33459\,
            PADOUT => \N__33458\,
            PADIN => \N__33457\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15439\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33450\,
            DIN => \N__33449\,
            DOUT => \N__33448\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33450\,
            PADOUT => \N__33449\,
            PADIN => \N__33448\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33441\,
            DIN => \N__33440\,
            DOUT => \N__33439\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33441\,
            PADOUT => \N__33440\,
            PADIN => \N__33439\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33432\,
            DIN => \N__33431\,
            DOUT => \N__33430\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33432\,
            PADOUT => \N__33431\,
            PADIN => \N__33430\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33423\,
            DIN => \N__33422\,
            DOUT => \N__33421\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33423\,
            PADOUT => \N__33422\,
            PADIN => \N__33421\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33414\,
            DIN => \N__33413\,
            DOUT => \N__33412\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33414\,
            PADOUT => \N__33413\,
            PADIN => \N__33412\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33405\,
            DIN => \N__33404\,
            DOUT => \N__33403\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33405\,
            PADOUT => \N__33404\,
            PADIN => \N__33403\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15884\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33396\,
            DIN => \N__33395\,
            DOUT => \N__33394\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33396\,
            PADOUT => \N__33395\,
            PADIN => \N__33394\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33387\,
            DIN => \N__33386\,
            DOUT => \N__33385\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33387\,
            PADOUT => \N__33386\,
            PADIN => \N__33385\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__33026\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33378\,
            DIN => \N__33377\,
            DOUT => \N__33376\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33378\,
            PADOUT => \N__33377\,
            PADIN => \N__33376\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33369\,
            DIN => \N__33368\,
            DOUT => \N__33367\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33369\,
            PADOUT => \N__33368\,
            PADIN => \N__33367\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33360\,
            DIN => \N__33359\,
            DOUT => \N__33358\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33360\,
            PADOUT => \N__33359\,
            PADIN => \N__33358\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33351\,
            DIN => \N__33350\,
            DOUT => \N__33349\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33351\,
            PADOUT => \N__33350\,
            PADIN => \N__33349\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33342\,
            DIN => \N__33341\,
            DOUT => \N__33340\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33342\,
            PADOUT => \N__33341\,
            PADIN => \N__33340\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16181\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33333\,
            DIN => \N__33332\,
            DOUT => \N__33331\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33333\,
            PADOUT => \N__33332\,
            PADIN => \N__33331\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33324\,
            DIN => \N__33323\,
            DOUT => \N__33322\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33324\,
            PADOUT => \N__33323\,
            PADIN => \N__33322\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29630\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33315\,
            DIN => \N__33314\,
            DOUT => \N__33313\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33315\,
            PADOUT => \N__33314\,
            PADIN => \N__33313\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33306\,
            DIN => \N__33305\,
            DOUT => \N__33304\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33306\,
            PADOUT => \N__33305\,
            PADIN => \N__33304\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25181\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33297\,
            DIN => \N__33296\,
            DOUT => \N__33295\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33297\,
            PADOUT => \N__33296\,
            PADIN => \N__33295\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16226\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33288\,
            DIN => \N__33287\,
            DOUT => \N__33286\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33288\,
            PADOUT => \N__33287\,
            PADIN => \N__33286\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33279\,
            DIN => \N__33278\,
            DOUT => \N__33277\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33279\,
            PADOUT => \N__33278\,
            PADIN => \N__33277\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33270\,
            DIN => \N__33269\,
            DOUT => \N__33268\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33270\,
            PADOUT => \N__33269\,
            PADIN => \N__33268\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33261\,
            DIN => \N__33260\,
            DOUT => \N__33259\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33261\,
            PADOUT => \N__33260\,
            PADIN => \N__33259\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25202\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33252\,
            DIN => \N__33251\,
            DOUT => \N__33250\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33252\,
            PADOUT => \N__33251\,
            PADIN => \N__33250\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32969\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33243\,
            DIN => \N__33242\,
            DOUT => \N__33241\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33243\,
            PADOUT => \N__33242\,
            PADIN => \N__33241\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33234\,
            DIN => \N__33233\,
            DOUT => \N__33232\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33234\,
            PADOUT => \N__33233\,
            PADIN => \N__33232\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33225\,
            DIN => \N__33224\,
            DOUT => \N__33223\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33225\,
            PADOUT => \N__33224\,
            PADIN => \N__33223\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33216\,
            DIN => \N__33215\,
            DOUT => \N__33214\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33216\,
            PADOUT => \N__33215\,
            PADIN => \N__33214\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33207\,
            DIN => \N__33206\,
            DOUT => \N__33205\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33207\,
            PADOUT => \N__33206\,
            PADIN => \N__33205\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33198\,
            DIN => \N__33197\,
            DOUT => \N__33196\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33198\,
            PADOUT => \N__33197\,
            PADIN => \N__33196\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33189\,
            DIN => \N__33188\,
            DOUT => \N__33187\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33189\,
            PADOUT => \N__33188\,
            PADIN => \N__33187\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15440\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33180\,
            DIN => \N__33179\,
            DOUT => \N__33178\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33180\,
            PADOUT => \N__33179\,
            PADIN => \N__33178\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__7709\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33158\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__33158\,
            I => \N__33155\
        );

    \I__7707\ : Span4Mux_v
    port map (
            O => \N__33155\,
            I => \N__33152\
        );

    \I__7706\ : Span4Mux_h
    port map (
            O => \N__33152\,
            I => \N__33149\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__33149\,
            I => \N__33146\
        );

    \I__7704\ : Span4Mux_v
    port map (
            O => \N__33146\,
            I => \N__33141\
        );

    \I__7703\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33136\
        );

    \I__7702\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33136\
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__33141\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__33136\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__7699\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33124\
        );

    \I__7698\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33120\
        );

    \I__7697\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33117\
        );

    \I__7696\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33112\
        );

    \I__7695\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33112\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__33124\,
            I => \N__33109\
        );

    \I__7693\ : InMux
    port map (
            O => \N__33123\,
            I => \N__33106\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__33120\,
            I => \N__33101\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33101\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__33098\
        );

    \I__7689\ : Span4Mux_v
    port map (
            O => \N__33109\,
            I => \N__33095\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__33106\,
            I => \N__33092\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__33101\,
            I => \N__33087\
        );

    \I__7686\ : Span4Mux_s2_v
    port map (
            O => \N__33098\,
            I => \N__33087\
        );

    \I__7685\ : Span4Mux_h
    port map (
            O => \N__33095\,
            I => \N__33081\
        );

    \I__7684\ : Span4Mux_v
    port map (
            O => \N__33092\,
            I => \N__33078\
        );

    \I__7683\ : Span4Mux_h
    port map (
            O => \N__33087\,
            I => \N__33074\
        );

    \I__7682\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33069\
        );

    \I__7681\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33069\
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__33084\,
            I => \N__33064\
        );

    \I__7679\ : Span4Mux_v
    port map (
            O => \N__33081\,
            I => \N__33060\
        );

    \I__7678\ : Span4Mux_h
    port map (
            O => \N__33078\,
            I => \N__33057\
        );

    \I__7677\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33054\
        );

    \I__7676\ : Span4Mux_v
    port map (
            O => \N__33074\,
            I => \N__33049\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__33069\,
            I => \N__33049\
        );

    \I__7674\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33044\
        );

    \I__7673\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33044\
        );

    \I__7672\ : InMux
    port map (
            O => \N__33064\,
            I => \N__33039\
        );

    \I__7671\ : InMux
    port map (
            O => \N__33063\,
            I => \N__33039\
        );

    \I__7670\ : Odrv4
    port map (
            O => \N__33060\,
            I => \VCCST_EN_i_1\
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__33057\,
            I => \VCCST_EN_i_1\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__33054\,
            I => \VCCST_EN_i_1\
        );

    \I__7667\ : Odrv4
    port map (
            O => \N__33049\,
            I => \VCCST_EN_i_1\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__33044\,
            I => \VCCST_EN_i_1\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__33039\,
            I => \VCCST_EN_i_1\
        );

    \I__7664\ : IoInMux
    port map (
            O => \N__33026\,
            I => \N__33023\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__33023\,
            I => vpp_en
        );

    \I__7662\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33017\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__33017\,
            I => \N__33014\
        );

    \I__7660\ : Span4Mux_s2_h
    port map (
            O => \N__33014\,
            I => \N__33011\
        );

    \I__7659\ : Sp12to4
    port map (
            O => \N__33011\,
            I => \N__33008\
        );

    \I__7658\ : Span12Mux_v
    port map (
            O => \N__33008\,
            I => \N__33005\
        );

    \I__7657\ : Odrv12
    port map (
            O => \N__33005\,
            I => vccst_cpu_ok
        );

    \I__7656\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32999\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__32999\,
            I => \N__32996\
        );

    \I__7654\ : IoSpan4Mux
    port map (
            O => \N__32996\,
            I => \N__32993\
        );

    \I__7653\ : IoSpan4Mux
    port map (
            O => \N__32993\,
            I => \N__32990\
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__32990\,
            I => v5s_ok
        );

    \I__7651\ : CascadeMux
    port map (
            O => \N__32987\,
            I => \N__32984\
        );

    \I__7650\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32981\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__32981\,
            I => \N__32978\
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__32978\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_1\
        );

    \I__7647\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32972\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__32972\,
            I => v33s_ok
        );

    \I__7645\ : IoInMux
    port map (
            O => \N__32969\,
            I => \N__32966\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__32966\,
            I => \N__32963\
        );

    \I__7643\ : Span4Mux_s3_v
    port map (
            O => \N__32963\,
            I => \N__32960\
        );

    \I__7642\ : Odrv4
    port map (
            O => \N__32960\,
            I => vccin_en
        );

    \I__7641\ : CascadeMux
    port map (
            O => \N__32957\,
            I => \N__32950\
        );

    \I__7640\ : CascadeMux
    port map (
            O => \N__32956\,
            I => \N__32945\
        );

    \I__7639\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32941\
        );

    \I__7638\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32937\
        );

    \I__7637\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32934\
        );

    \I__7636\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32929\
        );

    \I__7635\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32929\
        );

    \I__7634\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32926\
        );

    \I__7633\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32923\
        );

    \I__7632\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32920\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__32941\,
            I => \N__32917\
        );

    \I__7630\ : CascadeMux
    port map (
            O => \N__32940\,
            I => \N__32914\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__32937\,
            I => \N__32910\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__32934\,
            I => \N__32905\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__32929\,
            I => \N__32905\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__32926\,
            I => \N__32902\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__32923\,
            I => \N__32899\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32896\
        );

    \I__7623\ : Span12Mux_s7_h
    port map (
            O => \N__32917\,
            I => \N__32893\
        );

    \I__7622\ : InMux
    port map (
            O => \N__32914\,
            I => \N__32890\
        );

    \I__7621\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32887\
        );

    \I__7620\ : Span4Mux_v
    port map (
            O => \N__32910\,
            I => \N__32880\
        );

    \I__7619\ : Span4Mux_v
    port map (
            O => \N__32905\,
            I => \N__32880\
        );

    \I__7618\ : Span4Mux_v
    port map (
            O => \N__32902\,
            I => \N__32880\
        );

    \I__7617\ : Span4Mux_s3_h
    port map (
            O => \N__32899\,
            I => \N__32875\
        );

    \I__7616\ : Span4Mux_s3_h
    port map (
            O => \N__32896\,
            I => \N__32875\
        );

    \I__7615\ : Odrv12
    port map (
            O => \N__32893\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__32890\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__32887\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7612\ : Odrv4
    port map (
            O => \N__32880\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__32875\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7610\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32861\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__32861\,
            I => \POWERLED.un1_dutycycle_53_axb_3\
        );

    \I__7608\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32855\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__32855\,
            I => \N__32852\
        );

    \I__7606\ : Odrv12
    port map (
            O => \N__32852\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_2\
        );

    \I__7605\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__32846\,
            I => \POWERLED.dutycycle_eena_13_c_1\
        );

    \I__7603\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32837\
        );

    \I__7602\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32837\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32828\
        );

    \I__7600\ : CascadeMux
    port map (
            O => \N__32836\,
            I => \N__32822\
        );

    \I__7599\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32816\
        );

    \I__7598\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32816\
        );

    \I__7597\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32806\
        );

    \I__7596\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32806\
        );

    \I__7595\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32803\
        );

    \I__7594\ : Span4Mux_s1_v
    port map (
            O => \N__32828\,
            I => \N__32800\
        );

    \I__7593\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32797\
        );

    \I__7592\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32794\
        );

    \I__7591\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32789\
        );

    \I__7590\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32784\
        );

    \I__7589\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32784\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32780\
        );

    \I__7587\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32775\
        );

    \I__7586\ : InMux
    port map (
            O => \N__32814\,
            I => \N__32775\
        );

    \I__7585\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32772\
        );

    \I__7584\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32769\
        );

    \I__7583\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32765\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__32806\,
            I => \N__32754\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__32803\,
            I => \N__32754\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__32800\,
            I => \N__32754\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__32797\,
            I => \N__32754\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__32794\,
            I => \N__32754\
        );

    \I__7577\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32749\
        );

    \I__7576\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32749\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__32789\,
            I => \N__32746\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__32784\,
            I => \N__32741\
        );

    \I__7573\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32737\
        );

    \I__7572\ : Span4Mux_v
    port map (
            O => \N__32780\,
            I => \N__32732\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__32775\,
            I => \N__32732\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32727\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__32769\,
            I => \N__32727\
        );

    \I__7568\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32724\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__32765\,
            I => \N__32715\
        );

    \I__7566\ : Span4Mux_v
    port map (
            O => \N__32754\,
            I => \N__32715\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__32749\,
            I => \N__32715\
        );

    \I__7564\ : Span4Mux_s1_h
    port map (
            O => \N__32746\,
            I => \N__32715\
        );

    \I__7563\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32712\
        );

    \I__7562\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32709\
        );

    \I__7561\ : Span4Mux_s3_h
    port map (
            O => \N__32741\,
            I => \N__32706\
        );

    \I__7560\ : InMux
    port map (
            O => \N__32740\,
            I => \N__32703\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__32737\,
            I => \N__32698\
        );

    \I__7558\ : Span4Mux_s3_h
    port map (
            O => \N__32732\,
            I => \N__32698\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__32727\,
            I => \N__32691\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32691\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__32715\,
            I => \N__32691\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__32712\,
            I => \POWERLED.N_430\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__32709\,
            I => \POWERLED.N_430\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__32706\,
            I => \POWERLED.N_430\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__32703\,
            I => \POWERLED.N_430\
        );

    \I__7550\ : Odrv4
    port map (
            O => \N__32698\,
            I => \POWERLED.N_430\
        );

    \I__7549\ : Odrv4
    port map (
            O => \N__32691\,
            I => \POWERLED.N_430\
        );

    \I__7548\ : CascadeMux
    port map (
            O => \N__32678\,
            I => \POWERLED.un1_clk_100khz_51_and_i_3_cascade_\
        );

    \I__7547\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32664\
        );

    \I__7546\ : IoInMux
    port map (
            O => \N__32674\,
            I => \N__32661\
        );

    \I__7545\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32656\
        );

    \I__7544\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32656\
        );

    \I__7543\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32653\
        );

    \I__7542\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32650\
        );

    \I__7541\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32647\
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__32668\,
            I => \N__32641\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__32667\,
            I => \N__32634\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__32664\,
            I => \N__32631\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32621\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__32656\,
            I => \N__32621\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32614\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__32650\,
            I => \N__32614\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32614\
        );

    \I__7532\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32611\
        );

    \I__7531\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32608\
        );

    \I__7530\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32604\
        );

    \I__7529\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32601\
        );

    \I__7528\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32594\
        );

    \I__7527\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32594\
        );

    \I__7526\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32594\
        );

    \I__7525\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32590\
        );

    \I__7524\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32587\
        );

    \I__7523\ : Span4Mux_v
    port map (
            O => \N__32631\,
            I => \N__32584\
        );

    \I__7522\ : InMux
    port map (
            O => \N__32630\,
            I => \N__32579\
        );

    \I__7521\ : InMux
    port map (
            O => \N__32629\,
            I => \N__32579\
        );

    \I__7520\ : CascadeMux
    port map (
            O => \N__32628\,
            I => \N__32576\
        );

    \I__7519\ : InMux
    port map (
            O => \N__32627\,
            I => \N__32570\
        );

    \I__7518\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32570\
        );

    \I__7517\ : Span4Mux_s3_v
    port map (
            O => \N__32621\,
            I => \N__32567\
        );

    \I__7516\ : Span4Mux_s3_v
    port map (
            O => \N__32614\,
            I => \N__32562\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__32611\,
            I => \N__32562\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__32608\,
            I => \N__32559\
        );

    \I__7513\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32556\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__32604\,
            I => \N__32553\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__32601\,
            I => \N__32548\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__32594\,
            I => \N__32548\
        );

    \I__7509\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32545\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__32590\,
            I => \N__32542\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__32587\,
            I => \N__32539\
        );

    \I__7506\ : Span4Mux_h
    port map (
            O => \N__32584\,
            I => \N__32534\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__32579\,
            I => \N__32534\
        );

    \I__7504\ : InMux
    port map (
            O => \N__32576\,
            I => \N__32529\
        );

    \I__7503\ : InMux
    port map (
            O => \N__32575\,
            I => \N__32529\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32522\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__32567\,
            I => \N__32522\
        );

    \I__7500\ : Span4Mux_v
    port map (
            O => \N__32562\,
            I => \N__32522\
        );

    \I__7499\ : Span4Mux_s3_h
    port map (
            O => \N__32559\,
            I => \N__32515\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__32556\,
            I => \N__32515\
        );

    \I__7497\ : Span4Mux_s3_h
    port map (
            O => \N__32553\,
            I => \N__32515\
        );

    \I__7496\ : Span4Mux_s3_h
    port map (
            O => \N__32548\,
            I => \N__32510\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32510\
        );

    \I__7494\ : Span4Mux_s3_h
    port map (
            O => \N__32542\,
            I => \N__32507\
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__32539\,
            I => \G_141\
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__32534\,
            I => \G_141\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__32529\,
            I => \G_141\
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__32522\,
            I => \G_141\
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__32515\,
            I => \G_141\
        );

    \I__7488\ : Odrv4
    port map (
            O => \N__32510\,
            I => \G_141\
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__32507\,
            I => \G_141\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__32492\,
            I => \N__32489\
        );

    \I__7485\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32483\
        );

    \I__7484\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32483\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__32483\,
            I => \POWERLED.dutycycle_RNI0DF58Z0Z_5\
        );

    \I__7482\ : ClkMux
    port map (
            O => \N__32480\,
            I => \N__32476\
        );

    \I__7481\ : ClkMux
    port map (
            O => \N__32479\,
            I => \N__32473\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__32476\,
            I => \N__32454\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32454\
        );

    \I__7478\ : ClkMux
    port map (
            O => \N__32472\,
            I => \N__32451\
        );

    \I__7477\ : ClkMux
    port map (
            O => \N__32471\,
            I => \N__32446\
        );

    \I__7476\ : ClkMux
    port map (
            O => \N__32470\,
            I => \N__32443\
        );

    \I__7475\ : ClkMux
    port map (
            O => \N__32469\,
            I => \N__32440\
        );

    \I__7474\ : ClkMux
    port map (
            O => \N__32468\,
            I => \N__32437\
        );

    \I__7473\ : ClkMux
    port map (
            O => \N__32467\,
            I => \N__32432\
        );

    \I__7472\ : ClkMux
    port map (
            O => \N__32466\,
            I => \N__32427\
        );

    \I__7471\ : ClkMux
    port map (
            O => \N__32465\,
            I => \N__32424\
        );

    \I__7470\ : ClkMux
    port map (
            O => \N__32464\,
            I => \N__32420\
        );

    \I__7469\ : ClkMux
    port map (
            O => \N__32463\,
            I => \N__32416\
        );

    \I__7468\ : ClkMux
    port map (
            O => \N__32462\,
            I => \N__32413\
        );

    \I__7467\ : ClkMux
    port map (
            O => \N__32461\,
            I => \N__32408\
        );

    \I__7466\ : ClkMux
    port map (
            O => \N__32460\,
            I => \N__32403\
        );

    \I__7465\ : ClkMux
    port map (
            O => \N__32459\,
            I => \N__32398\
        );

    \I__7464\ : Span4Mux_s1_v
    port map (
            O => \N__32454\,
            I => \N__32392\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__32451\,
            I => \N__32392\
        );

    \I__7462\ : ClkMux
    port map (
            O => \N__32450\,
            I => \N__32389\
        );

    \I__7461\ : ClkMux
    port map (
            O => \N__32449\,
            I => \N__32386\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__32446\,
            I => \N__32381\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__32443\,
            I => \N__32377\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__32440\,
            I => \N__32372\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__32437\,
            I => \N__32372\
        );

    \I__7456\ : ClkMux
    port map (
            O => \N__32436\,
            I => \N__32369\
        );

    \I__7455\ : ClkMux
    port map (
            O => \N__32435\,
            I => \N__32366\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__32432\,
            I => \N__32363\
        );

    \I__7453\ : ClkMux
    port map (
            O => \N__32431\,
            I => \N__32360\
        );

    \I__7452\ : ClkMux
    port map (
            O => \N__32430\,
            I => \N__32357\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__32427\,
            I => \N__32351\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__32424\,
            I => \N__32346\
        );

    \I__7449\ : ClkMux
    port map (
            O => \N__32423\,
            I => \N__32343\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__32420\,
            I => \N__32339\
        );

    \I__7447\ : ClkMux
    port map (
            O => \N__32419\,
            I => \N__32336\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__32416\,
            I => \N__32329\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__32413\,
            I => \N__32326\
        );

    \I__7444\ : ClkMux
    port map (
            O => \N__32412\,
            I => \N__32323\
        );

    \I__7443\ : ClkMux
    port map (
            O => \N__32411\,
            I => \N__32319\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__32408\,
            I => \N__32313\
        );

    \I__7441\ : ClkMux
    port map (
            O => \N__32407\,
            I => \N__32310\
        );

    \I__7440\ : ClkMux
    port map (
            O => \N__32406\,
            I => \N__32306\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__32403\,
            I => \N__32303\
        );

    \I__7438\ : ClkMux
    port map (
            O => \N__32402\,
            I => \N__32300\
        );

    \I__7437\ : ClkMux
    port map (
            O => \N__32401\,
            I => \N__32296\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__32398\,
            I => \N__32293\
        );

    \I__7435\ : ClkMux
    port map (
            O => \N__32397\,
            I => \N__32290\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__32392\,
            I => \N__32285\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__32389\,
            I => \N__32285\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__32386\,
            I => \N__32276\
        );

    \I__7431\ : ClkMux
    port map (
            O => \N__32385\,
            I => \N__32273\
        );

    \I__7430\ : ClkMux
    port map (
            O => \N__32384\,
            I => \N__32270\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__32381\,
            I => \N__32266\
        );

    \I__7428\ : ClkMux
    port map (
            O => \N__32380\,
            I => \N__32262\
        );

    \I__7427\ : Span4Mux_v
    port map (
            O => \N__32377\,
            I => \N__32252\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__32372\,
            I => \N__32252\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32252\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__32366\,
            I => \N__32252\
        );

    \I__7423\ : Span4Mux_v
    port map (
            O => \N__32363\,
            I => \N__32245\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__32360\,
            I => \N__32245\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__32357\,
            I => \N__32245\
        );

    \I__7420\ : ClkMux
    port map (
            O => \N__32356\,
            I => \N__32242\
        );

    \I__7419\ : ClkMux
    port map (
            O => \N__32355\,
            I => \N__32239\
        );

    \I__7418\ : ClkMux
    port map (
            O => \N__32354\,
            I => \N__32236\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__32351\,
            I => \N__32232\
        );

    \I__7416\ : ClkMux
    port map (
            O => \N__32350\,
            I => \N__32229\
        );

    \I__7415\ : ClkMux
    port map (
            O => \N__32349\,
            I => \N__32221\
        );

    \I__7414\ : Span4Mux_s1_h
    port map (
            O => \N__32346\,
            I => \N__32215\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32215\
        );

    \I__7412\ : ClkMux
    port map (
            O => \N__32342\,
            I => \N__32212\
        );

    \I__7411\ : Span4Mux_s1_h
    port map (
            O => \N__32339\,
            I => \N__32207\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__32336\,
            I => \N__32207\
        );

    \I__7409\ : ClkMux
    port map (
            O => \N__32335\,
            I => \N__32202\
        );

    \I__7408\ : ClkMux
    port map (
            O => \N__32334\,
            I => \N__32198\
        );

    \I__7407\ : ClkMux
    port map (
            O => \N__32333\,
            I => \N__32195\
        );

    \I__7406\ : ClkMux
    port map (
            O => \N__32332\,
            I => \N__32192\
        );

    \I__7405\ : Span4Mux_h
    port map (
            O => \N__32329\,
            I => \N__32189\
        );

    \I__7404\ : Span4Mux_s1_h
    port map (
            O => \N__32326\,
            I => \N__32184\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__32323\,
            I => \N__32184\
        );

    \I__7402\ : ClkMux
    port map (
            O => \N__32322\,
            I => \N__32181\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__32319\,
            I => \N__32176\
        );

    \I__7400\ : ClkMux
    port map (
            O => \N__32318\,
            I => \N__32173\
        );

    \I__7399\ : ClkMux
    port map (
            O => \N__32317\,
            I => \N__32170\
        );

    \I__7398\ : ClkMux
    port map (
            O => \N__32316\,
            I => \N__32167\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__32313\,
            I => \N__32161\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__32310\,
            I => \N__32161\
        );

    \I__7395\ : ClkMux
    port map (
            O => \N__32309\,
            I => \N__32158\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32155\
        );

    \I__7393\ : Span4Mux_v
    port map (
            O => \N__32303\,
            I => \N__32150\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__32300\,
            I => \N__32150\
        );

    \I__7391\ : ClkMux
    port map (
            O => \N__32299\,
            I => \N__32147\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32144\
        );

    \I__7389\ : Span4Mux_h
    port map (
            O => \N__32293\,
            I => \N__32139\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__32290\,
            I => \N__32139\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__32285\,
            I => \N__32136\
        );

    \I__7386\ : ClkMux
    port map (
            O => \N__32284\,
            I => \N__32133\
        );

    \I__7385\ : ClkMux
    port map (
            O => \N__32283\,
            I => \N__32130\
        );

    \I__7384\ : ClkMux
    port map (
            O => \N__32282\,
            I => \N__32127\
        );

    \I__7383\ : ClkMux
    port map (
            O => \N__32281\,
            I => \N__32123\
        );

    \I__7382\ : ClkMux
    port map (
            O => \N__32280\,
            I => \N__32120\
        );

    \I__7381\ : ClkMux
    port map (
            O => \N__32279\,
            I => \N__32117\
        );

    \I__7380\ : Span4Mux_v
    port map (
            O => \N__32276\,
            I => \N__32112\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__32273\,
            I => \N__32112\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__32270\,
            I => \N__32109\
        );

    \I__7377\ : ClkMux
    port map (
            O => \N__32269\,
            I => \N__32106\
        );

    \I__7376\ : Span4Mux_s0_v
    port map (
            O => \N__32266\,
            I => \N__32103\
        );

    \I__7375\ : ClkMux
    port map (
            O => \N__32265\,
            I => \N__32100\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32097\
        );

    \I__7373\ : ClkMux
    port map (
            O => \N__32261\,
            I => \N__32094\
        );

    \I__7372\ : Span4Mux_v
    port map (
            O => \N__32252\,
            I => \N__32083\
        );

    \I__7371\ : Span4Mux_v
    port map (
            O => \N__32245\,
            I => \N__32083\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32083\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__32239\,
            I => \N__32083\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__32236\,
            I => \N__32083\
        );

    \I__7367\ : ClkMux
    port map (
            O => \N__32235\,
            I => \N__32080\
        );

    \I__7366\ : Span4Mux_v
    port map (
            O => \N__32232\,
            I => \N__32075\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__32229\,
            I => \N__32075\
        );

    \I__7364\ : ClkMux
    port map (
            O => \N__32228\,
            I => \N__32072\
        );

    \I__7363\ : ClkMux
    port map (
            O => \N__32227\,
            I => \N__32069\
        );

    \I__7362\ : ClkMux
    port map (
            O => \N__32226\,
            I => \N__32066\
        );

    \I__7361\ : ClkMux
    port map (
            O => \N__32225\,
            I => \N__32063\
        );

    \I__7360\ : ClkMux
    port map (
            O => \N__32224\,
            I => \N__32060\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__32221\,
            I => \N__32057\
        );

    \I__7358\ : ClkMux
    port map (
            O => \N__32220\,
            I => \N__32054\
        );

    \I__7357\ : Span4Mux_v
    port map (
            O => \N__32215\,
            I => \N__32047\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__32212\,
            I => \N__32047\
        );

    \I__7355\ : Span4Mux_h
    port map (
            O => \N__32207\,
            I => \N__32042\
        );

    \I__7354\ : ClkMux
    port map (
            O => \N__32206\,
            I => \N__32039\
        );

    \I__7353\ : ClkMux
    port map (
            O => \N__32205\,
            I => \N__32036\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__32202\,
            I => \N__32033\
        );

    \I__7351\ : ClkMux
    port map (
            O => \N__32201\,
            I => \N__32030\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32025\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__32195\,
            I => \N__32025\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__32192\,
            I => \N__32022\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__32189\,
            I => \N__32017\
        );

    \I__7346\ : Span4Mux_h
    port map (
            O => \N__32184\,
            I => \N__32017\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__32181\,
            I => \N__32014\
        );

    \I__7344\ : ClkMux
    port map (
            O => \N__32180\,
            I => \N__32011\
        );

    \I__7343\ : ClkMux
    port map (
            O => \N__32179\,
            I => \N__32008\
        );

    \I__7342\ : Span4Mux_s2_h
    port map (
            O => \N__32176\,
            I => \N__32003\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__32173\,
            I => \N__32003\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__32170\,
            I => \N__32000\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__32167\,
            I => \N__31997\
        );

    \I__7338\ : ClkMux
    port map (
            O => \N__32166\,
            I => \N__31994\
        );

    \I__7337\ : Span4Mux_v
    port map (
            O => \N__32161\,
            I => \N__31991\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__32158\,
            I => \N__31988\
        );

    \I__7335\ : Span4Mux_v
    port map (
            O => \N__32155\,
            I => \N__31981\
        );

    \I__7334\ : Span4Mux_h
    port map (
            O => \N__32150\,
            I => \N__31981\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__32147\,
            I => \N__31981\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__32144\,
            I => \N__31968\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__32139\,
            I => \N__31968\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__32136\,
            I => \N__31968\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__32133\,
            I => \N__31968\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__31968\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__32127\,
            I => \N__31968\
        );

    \I__7326\ : ClkMux
    port map (
            O => \N__32126\,
            I => \N__31965\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__32123\,
            I => \N__31958\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__31958\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__32117\,
            I => \N__31958\
        );

    \I__7322\ : Span4Mux_v
    port map (
            O => \N__32112\,
            I => \N__31947\
        );

    \I__7321\ : Span4Mux_v
    port map (
            O => \N__32109\,
            I => \N__31947\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__31947\
        );

    \I__7319\ : Span4Mux_h
    port map (
            O => \N__32103\,
            I => \N__31947\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__32100\,
            I => \N__31947\
        );

    \I__7317\ : IoSpan4Mux
    port map (
            O => \N__32097\,
            I => \N__31944\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__32094\,
            I => \N__31941\
        );

    \I__7315\ : Span4Mux_v
    port map (
            O => \N__32083\,
            I => \N__31936\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__32080\,
            I => \N__31936\
        );

    \I__7313\ : Span4Mux_v
    port map (
            O => \N__32075\,
            I => \N__31925\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__32072\,
            I => \N__31925\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__31925\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__31925\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__32063\,
            I => \N__31925\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__32060\,
            I => \N__31918\
        );

    \I__7307\ : Span4Mux_h
    port map (
            O => \N__32057\,
            I => \N__31918\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__32054\,
            I => \N__31918\
        );

    \I__7305\ : ClkMux
    port map (
            O => \N__32053\,
            I => \N__31915\
        );

    \I__7304\ : ClkMux
    port map (
            O => \N__32052\,
            I => \N__31912\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__32047\,
            I => \N__31909\
        );

    \I__7302\ : ClkMux
    port map (
            O => \N__32046\,
            I => \N__31906\
        );

    \I__7301\ : ClkMux
    port map (
            O => \N__32045\,
            I => \N__31903\
        );

    \I__7300\ : Span4Mux_v
    port map (
            O => \N__32042\,
            I => \N__31896\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__32039\,
            I => \N__31896\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__32036\,
            I => \N__31896\
        );

    \I__7297\ : Span4Mux_s2_h
    port map (
            O => \N__32033\,
            I => \N__31891\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__31891\
        );

    \I__7295\ : Span4Mux_v
    port map (
            O => \N__32025\,
            I => \N__31886\
        );

    \I__7294\ : Span4Mux_s1_h
    port map (
            O => \N__32022\,
            I => \N__31886\
        );

    \I__7293\ : Span4Mux_v
    port map (
            O => \N__32017\,
            I => \N__31877\
        );

    \I__7292\ : Span4Mux_v
    port map (
            O => \N__32014\,
            I => \N__31877\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__32011\,
            I => \N__31877\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__32008\,
            I => \N__31877\
        );

    \I__7289\ : Span4Mux_v
    port map (
            O => \N__32003\,
            I => \N__31868\
        );

    \I__7288\ : Span4Mux_s2_h
    port map (
            O => \N__32000\,
            I => \N__31868\
        );

    \I__7287\ : Span4Mux_s2_h
    port map (
            O => \N__31997\,
            I => \N__31868\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__31994\,
            I => \N__31868\
        );

    \I__7285\ : IoSpan4Mux
    port map (
            O => \N__31991\,
            I => \N__31863\
        );

    \I__7284\ : IoSpan4Mux
    port map (
            O => \N__31988\,
            I => \N__31863\
        );

    \I__7283\ : Span4Mux_v
    port map (
            O => \N__31981\,
            I => \N__31856\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__31968\,
            I => \N__31856\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__31965\,
            I => \N__31856\
        );

    \I__7280\ : Span4Mux_v
    port map (
            O => \N__31958\,
            I => \N__31851\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__31947\,
            I => \N__31851\
        );

    \I__7278\ : IoSpan4Mux
    port map (
            O => \N__31944\,
            I => \N__31846\
        );

    \I__7277\ : IoSpan4Mux
    port map (
            O => \N__31941\,
            I => \N__31846\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__31936\,
            I => \N__31837\
        );

    \I__7275\ : Span4Mux_v
    port map (
            O => \N__31925\,
            I => \N__31837\
        );

    \I__7274\ : Span4Mux_v
    port map (
            O => \N__31918\,
            I => \N__31837\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__31915\,
            I => \N__31837\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__31912\,
            I => \N__31833\
        );

    \I__7271\ : Span4Mux_h
    port map (
            O => \N__31909\,
            I => \N__31826\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__31906\,
            I => \N__31826\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__31903\,
            I => \N__31826\
        );

    \I__7268\ : Span4Mux_v
    port map (
            O => \N__31896\,
            I => \N__31821\
        );

    \I__7267\ : Span4Mux_h
    port map (
            O => \N__31891\,
            I => \N__31821\
        );

    \I__7266\ : Span4Mux_h
    port map (
            O => \N__31886\,
            I => \N__31814\
        );

    \I__7265\ : Span4Mux_v
    port map (
            O => \N__31877\,
            I => \N__31814\
        );

    \I__7264\ : Span4Mux_h
    port map (
            O => \N__31868\,
            I => \N__31814\
        );

    \I__7263\ : IoSpan4Mux
    port map (
            O => \N__31863\,
            I => \N__31807\
        );

    \I__7262\ : IoSpan4Mux
    port map (
            O => \N__31856\,
            I => \N__31807\
        );

    \I__7261\ : IoSpan4Mux
    port map (
            O => \N__31851\,
            I => \N__31807\
        );

    \I__7260\ : IoSpan4Mux
    port map (
            O => \N__31846\,
            I => \N__31802\
        );

    \I__7259\ : IoSpan4Mux
    port map (
            O => \N__31837\,
            I => \N__31802\
        );

    \I__7258\ : ClkMux
    port map (
            O => \N__31836\,
            I => \N__31799\
        );

    \I__7257\ : Sp12to4
    port map (
            O => \N__31833\,
            I => \N__31794\
        );

    \I__7256\ : Sp12to4
    port map (
            O => \N__31826\,
            I => \N__31794\
        );

    \I__7255\ : Odrv4
    port map (
            O => \N__31821\,
            I => fpga_osc
        );

    \I__7254\ : Odrv4
    port map (
            O => \N__31814\,
            I => fpga_osc
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__31807\,
            I => fpga_osc
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__31802\,
            I => fpga_osc
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__31799\,
            I => fpga_osc
        );

    \I__7250\ : Odrv12
    port map (
            O => \N__31794\,
            I => fpga_osc
        );

    \I__7249\ : SRMux
    port map (
            O => \N__31781\,
            I => \N__31777\
        );

    \I__7248\ : SRMux
    port map (
            O => \N__31780\,
            I => \N__31774\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__31777\,
            I => \N__31768\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__31774\,
            I => \N__31764\
        );

    \I__7245\ : SRMux
    port map (
            O => \N__31773\,
            I => \N__31761\
        );

    \I__7244\ : SRMux
    port map (
            O => \N__31772\,
            I => \N__31758\
        );

    \I__7243\ : SRMux
    port map (
            O => \N__31771\,
            I => \N__31751\
        );

    \I__7242\ : Span4Mux_h
    port map (
            O => \N__31768\,
            I => \N__31747\
        );

    \I__7241\ : SRMux
    port map (
            O => \N__31767\,
            I => \N__31744\
        );

    \I__7240\ : Span4Mux_h
    port map (
            O => \N__31764\,
            I => \N__31741\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__31761\,
            I => \N__31738\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__31758\,
            I => \N__31735\
        );

    \I__7237\ : SRMux
    port map (
            O => \N__31757\,
            I => \N__31732\
        );

    \I__7236\ : SRMux
    port map (
            O => \N__31756\,
            I => \N__31728\
        );

    \I__7235\ : SRMux
    port map (
            O => \N__31755\,
            I => \N__31725\
        );

    \I__7234\ : SRMux
    port map (
            O => \N__31754\,
            I => \N__31722\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__31751\,
            I => \N__31718\
        );

    \I__7232\ : SRMux
    port map (
            O => \N__31750\,
            I => \N__31715\
        );

    \I__7231\ : Span4Mux_s1_v
    port map (
            O => \N__31747\,
            I => \N__31710\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__31744\,
            I => \N__31710\
        );

    \I__7229\ : Span4Mux_s0_v
    port map (
            O => \N__31741\,
            I => \N__31707\
        );

    \I__7228\ : Span4Mux_s1_h
    port map (
            O => \N__31738\,
            I => \N__31700\
        );

    \I__7227\ : Span4Mux_v
    port map (
            O => \N__31735\,
            I => \N__31700\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__31732\,
            I => \N__31700\
        );

    \I__7225\ : SRMux
    port map (
            O => \N__31731\,
            I => \N__31697\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__31728\,
            I => \N__31694\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31691\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31688\
        );

    \I__7221\ : SRMux
    port map (
            O => \N__31721\,
            I => \N__31685\
        );

    \I__7220\ : Span4Mux_h
    port map (
            O => \N__31718\,
            I => \N__31680\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31680\
        );

    \I__7218\ : Span4Mux_v
    port map (
            O => \N__31710\,
            I => \N__31677\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__31707\,
            I => \N__31672\
        );

    \I__7216\ : Span4Mux_h
    port map (
            O => \N__31700\,
            I => \N__31672\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__31697\,
            I => \N__31669\
        );

    \I__7214\ : Span4Mux_s0_h
    port map (
            O => \N__31694\,
            I => \N__31664\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__31691\,
            I => \N__31664\
        );

    \I__7212\ : Span4Mux_v
    port map (
            O => \N__31688\,
            I => \N__31657\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__31685\,
            I => \N__31657\
        );

    \I__7210\ : Span4Mux_s3_v
    port map (
            O => \N__31680\,
            I => \N__31657\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__31677\,
            I => \N__31654\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__31672\,
            I => \N__31651\
        );

    \I__7207\ : Span4Mux_v
    port map (
            O => \N__31669\,
            I => \N__31644\
        );

    \I__7206\ : Span4Mux_h
    port map (
            O => \N__31664\,
            I => \N__31644\
        );

    \I__7205\ : Span4Mux_v
    port map (
            O => \N__31657\,
            I => \N__31644\
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__31654\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__31651\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__31644\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__7201\ : CascadeMux
    port map (
            O => \N__31637\,
            I => \N__31634\
        );

    \I__7200\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31630\
        );

    \I__7199\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31627\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__31630\,
            I => \POWERLED.dutycycle_en_8\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__31627\,
            I => \POWERLED.dutycycle_en_8\
        );

    \I__7196\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31618\
        );

    \I__7195\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31615\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__31618\,
            I => \N__31610\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__31615\,
            I => \N__31610\
        );

    \I__7192\ : Span4Mux_v
    port map (
            O => \N__31610\,
            I => \N__31607\
        );

    \I__7191\ : Odrv4
    port map (
            O => \N__31607\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\
        );

    \I__7190\ : CascadeMux
    port map (
            O => \N__31604\,
            I => \N__31600\
        );

    \I__7189\ : InMux
    port map (
            O => \N__31603\,
            I => \N__31595\
        );

    \I__7188\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31595\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__31595\,
            I => \POWERLED.dutycycleZ1Z_3\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__31592\,
            I => \N__31576\
        );

    \I__7185\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31572\
        );

    \I__7184\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31569\
        );

    \I__7183\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31560\
        );

    \I__7182\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31557\
        );

    \I__7181\ : InMux
    port map (
            O => \N__31587\,
            I => \N__31554\
        );

    \I__7180\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31545\
        );

    \I__7179\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31545\
        );

    \I__7178\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31545\
        );

    \I__7177\ : InMux
    port map (
            O => \N__31583\,
            I => \N__31545\
        );

    \I__7176\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31540\
        );

    \I__7175\ : InMux
    port map (
            O => \N__31581\,
            I => \N__31540\
        );

    \I__7174\ : InMux
    port map (
            O => \N__31580\,
            I => \N__31535\
        );

    \I__7173\ : InMux
    port map (
            O => \N__31579\,
            I => \N__31535\
        );

    \I__7172\ : InMux
    port map (
            O => \N__31576\,
            I => \N__31530\
        );

    \I__7171\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31530\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__31572\,
            I => \N__31527\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__31569\,
            I => \N__31524\
        );

    \I__7168\ : InMux
    port map (
            O => \N__31568\,
            I => \N__31515\
        );

    \I__7167\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31515\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31515\
        );

    \I__7165\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31515\
        );

    \I__7164\ : InMux
    port map (
            O => \N__31564\,
            I => \N__31512\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__31563\,
            I => \N__31509\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__31560\,
            I => \N__31505\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__31557\,
            I => \N__31502\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31499\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__31545\,
            I => \N__31488\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__31540\,
            I => \N__31488\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__31535\,
            I => \N__31488\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__31530\,
            I => \N__31488\
        );

    \I__7155\ : Span4Mux_s3_h
    port map (
            O => \N__31527\,
            I => \N__31479\
        );

    \I__7154\ : Span4Mux_v
    port map (
            O => \N__31524\,
            I => \N__31479\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__31515\,
            I => \N__31479\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__31512\,
            I => \N__31479\
        );

    \I__7151\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31474\
        );

    \I__7150\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31474\
        );

    \I__7149\ : Span12Mux_s10_h
    port map (
            O => \N__31505\,
            I => \N__31471\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__31502\,
            I => \N__31468\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__31499\,
            I => \N__31465\
        );

    \I__7146\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31460\
        );

    \I__7145\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31460\
        );

    \I__7144\ : Span4Mux_s3_v
    port map (
            O => \N__31488\,
            I => \N__31453\
        );

    \I__7143\ : Span4Mux_v
    port map (
            O => \N__31479\,
            I => \N__31453\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__31474\,
            I => \N__31453\
        );

    \I__7141\ : Odrv12
    port map (
            O => \N__31471\,
            I => \POWERLED.N_421\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__31468\,
            I => \POWERLED.N_421\
        );

    \I__7139\ : Odrv4
    port map (
            O => \N__31465\,
            I => \POWERLED.N_421\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__31460\,
            I => \POWERLED.N_421\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__31453\,
            I => \POWERLED.N_421\
        );

    \I__7136\ : CascadeMux
    port map (
            O => \N__31442\,
            I => \POWERLED.dutycycleZ0Z_8_cascade_\
        );

    \I__7135\ : CascadeMux
    port map (
            O => \N__31439\,
            I => \POWERLED.un1_dutycycle_53_axb_3_1_cascade_\
        );

    \I__7134\ : CascadeMux
    port map (
            O => \N__31436\,
            I => \N__31427\
        );

    \I__7133\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31418\
        );

    \I__7132\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31413\
        );

    \I__7131\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31413\
        );

    \I__7130\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31410\
        );

    \I__7129\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31407\
        );

    \I__7128\ : CascadeMux
    port map (
            O => \N__31430\,
            I => \N__31402\
        );

    \I__7127\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31395\
        );

    \I__7126\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31392\
        );

    \I__7125\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31385\
        );

    \I__7124\ : InMux
    port map (
            O => \N__31424\,
            I => \N__31385\
        );

    \I__7123\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31385\
        );

    \I__7122\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31380\
        );

    \I__7121\ : InMux
    port map (
            O => \N__31421\,
            I => \N__31380\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__31418\,
            I => \N__31377\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__31413\,
            I => \N__31374\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31369\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__31407\,
            I => \N__31369\
        );

    \I__7116\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31358\
        );

    \I__7115\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31358\
        );

    \I__7114\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31358\
        );

    \I__7113\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31358\
        );

    \I__7112\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31358\
        );

    \I__7111\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31353\
        );

    \I__7110\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31353\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__31395\,
            I => \N__31348\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__31392\,
            I => \N__31348\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__31385\,
            I => \N__31345\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31340\
        );

    \I__7105\ : Span4Mux_s2_h
    port map (
            O => \N__31377\,
            I => \N__31340\
        );

    \I__7104\ : Span4Mux_s2_h
    port map (
            O => \N__31374\,
            I => \N__31337\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__31369\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__31358\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__31353\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__7100\ : Odrv4
    port map (
            O => \N__31348\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__7099\ : Odrv4
    port map (
            O => \N__31345\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__31340\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__7097\ : Odrv4
    port map (
            O => \N__31337\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__31322\,
            I => \N__31318\
        );

    \I__7095\ : InMux
    port map (
            O => \N__31321\,
            I => \N__31315\
        );

    \I__7094\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31311\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__31315\,
            I => \N__31302\
        );

    \I__7092\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31299\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__31311\,
            I => \N__31294\
        );

    \I__7090\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31291\
        );

    \I__7089\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31288\
        );

    \I__7088\ : InMux
    port map (
            O => \N__31308\,
            I => \N__31285\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__31307\,
            I => \N__31282\
        );

    \I__7086\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31277\
        );

    \I__7085\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31277\
        );

    \I__7084\ : Span4Mux_v
    port map (
            O => \N__31302\,
            I => \N__31273\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__31299\,
            I => \N__31270\
        );

    \I__7082\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31265\
        );

    \I__7081\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31265\
        );

    \I__7080\ : Span4Mux_h
    port map (
            O => \N__31294\,
            I => \N__31260\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31257\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31252\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__31285\,
            I => \N__31252\
        );

    \I__7076\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31249\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__31277\,
            I => \N__31244\
        );

    \I__7074\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31241\
        );

    \I__7073\ : Span4Mux_h
    port map (
            O => \N__31273\,
            I => \N__31238\
        );

    \I__7072\ : Span4Mux_v
    port map (
            O => \N__31270\,
            I => \N__31233\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__31265\,
            I => \N__31233\
        );

    \I__7070\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31230\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31227\
        );

    \I__7068\ : Span4Mux_v
    port map (
            O => \N__31260\,
            I => \N__31222\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__31257\,
            I => \N__31222\
        );

    \I__7066\ : Span4Mux_v
    port map (
            O => \N__31252\,
            I => \N__31217\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31217\
        );

    \I__7064\ : InMux
    port map (
            O => \N__31248\,
            I => \N__31212\
        );

    \I__7063\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31212\
        );

    \I__7062\ : Span4Mux_h
    port map (
            O => \N__31244\,
            I => \N__31199\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__31241\,
            I => \N__31199\
        );

    \I__7060\ : Span4Mux_s0_h
    port map (
            O => \N__31238\,
            I => \N__31199\
        );

    \I__7059\ : Span4Mux_h
    port map (
            O => \N__31233\,
            I => \N__31199\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__31230\,
            I => \N__31199\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31199\
        );

    \I__7056\ : Odrv4
    port map (
            O => \N__31222\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__31217\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__31212\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__31199\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__7052\ : CascadeMux
    port map (
            O => \N__31190\,
            I => \POWERLED.un1_i3_mux_cascade_\
        );

    \I__7051\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31183\
        );

    \I__7050\ : CascadeMux
    port map (
            O => \N__31186\,
            I => \N__31180\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31177\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31180\,
            I => \N__31174\
        );

    \I__7047\ : Odrv12
    port map (
            O => \N__31177\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__31174\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31166\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__31166\,
            I => \N__31163\
        );

    \I__7043\ : Span4Mux_h
    port map (
            O => \N__31163\,
            I => \N__31160\
        );

    \I__7042\ : Span4Mux_h
    port map (
            O => \N__31160\,
            I => \N__31157\
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__31157\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_5\
        );

    \I__7040\ : CascadeMux
    port map (
            O => \N__31154\,
            I => \N__31141\
        );

    \I__7039\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31133\
        );

    \I__7038\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31133\
        );

    \I__7037\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31133\
        );

    \I__7036\ : InMux
    port map (
            O => \N__31150\,
            I => \N__31128\
        );

    \I__7035\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31128\
        );

    \I__7034\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31123\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31123\
        );

    \I__7032\ : CascadeMux
    port map (
            O => \N__31146\,
            I => \N__31119\
        );

    \I__7031\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31116\
        );

    \I__7030\ : InMux
    port map (
            O => \N__31144\,
            I => \N__31109\
        );

    \I__7029\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31109\
        );

    \I__7028\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31109\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__31133\,
            I => \N__31106\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31097\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__31123\,
            I => \N__31097\
        );

    \I__7024\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31094\
        );

    \I__7023\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31091\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__31116\,
            I => \N__31084\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__31109\,
            I => \N__31079\
        );

    \I__7020\ : Span4Mux_s2_v
    port map (
            O => \N__31106\,
            I => \N__31079\
        );

    \I__7019\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31076\
        );

    \I__7018\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31069\
        );

    \I__7017\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31069\
        );

    \I__7016\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31069\
        );

    \I__7015\ : Span4Mux_v
    port map (
            O => \N__31097\,
            I => \N__31064\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__31094\,
            I => \N__31064\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__31091\,
            I => \N__31061\
        );

    \I__7012\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31056\
        );

    \I__7011\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31056\
        );

    \I__7010\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31051\
        );

    \I__7009\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31051\
        );

    \I__7008\ : Span4Mux_v
    port map (
            O => \N__31084\,
            I => \N__31046\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__31079\,
            I => \N__31046\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__31076\,
            I => \N__31039\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__31069\,
            I => \N__31039\
        );

    \I__7004\ : Span4Mux_h
    port map (
            O => \N__31064\,
            I => \N__31039\
        );

    \I__7003\ : Odrv12
    port map (
            O => \N__31061\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__31056\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__31051\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__31046\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__6999\ : Odrv4
    port map (
            O => \N__31039\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__6997\ : InMux
    port map (
            O => \N__31025\,
            I => \N__31015\
        );

    \I__6996\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31010\
        );

    \I__6995\ : InMux
    port map (
            O => \N__31023\,
            I => \N__31007\
        );

    \I__6994\ : CascadeMux
    port map (
            O => \N__31022\,
            I => \N__31004\
        );

    \I__6993\ : InMux
    port map (
            O => \N__31021\,
            I => \N__30999\
        );

    \I__6992\ : InMux
    port map (
            O => \N__31020\,
            I => \N__30994\
        );

    \I__6991\ : InMux
    port map (
            O => \N__31019\,
            I => \N__30994\
        );

    \I__6990\ : InMux
    port map (
            O => \N__31018\,
            I => \N__30991\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__31015\,
            I => \N__30988\
        );

    \I__6988\ : InMux
    port map (
            O => \N__31014\,
            I => \N__30983\
        );

    \I__6987\ : InMux
    port map (
            O => \N__31013\,
            I => \N__30983\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__30978\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__31007\,
            I => \N__30975\
        );

    \I__6984\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30968\
        );

    \I__6983\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30968\
        );

    \I__6982\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30968\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30963\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__30994\,
            I => \N__30963\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__30991\,
            I => \N__30960\
        );

    \I__6978\ : Span12Mux_s4_v
    port map (
            O => \N__30988\,
            I => \N__30955\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__30983\,
            I => \N__30955\
        );

    \I__6976\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30950\
        );

    \I__6975\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30950\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__30978\,
            I => \N__30945\
        );

    \I__6973\ : Span4Mux_h
    port map (
            O => \N__30975\,
            I => \N__30945\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__30968\,
            I => \N__30938\
        );

    \I__6971\ : Span4Mux_h
    port map (
            O => \N__30963\,
            I => \N__30938\
        );

    \I__6970\ : Span4Mux_h
    port map (
            O => \N__30960\,
            I => \N__30938\
        );

    \I__6969\ : Odrv12
    port map (
            O => \N__30955\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__30950\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6967\ : Odrv4
    port map (
            O => \N__30945\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__30938\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6965\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30921\
        );

    \I__6964\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30913\
        );

    \I__6963\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30906\
        );

    \I__6962\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30906\
        );

    \I__6961\ : InMux
    port map (
            O => \N__30925\,
            I => \N__30906\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__30924\,
            I => \N__30902\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30899\
        );

    \I__6958\ : CascadeMux
    port map (
            O => \N__30920\,
            I => \N__30896\
        );

    \I__6957\ : CascadeMux
    port map (
            O => \N__30919\,
            I => \N__30893\
        );

    \I__6956\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30886\
        );

    \I__6955\ : InMux
    port map (
            O => \N__30917\,
            I => \N__30886\
        );

    \I__6954\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30886\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30883\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__30906\,
            I => \N__30880\
        );

    \I__6951\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30875\
        );

    \I__6950\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30875\
        );

    \I__6949\ : Span12Mux_s6_v
    port map (
            O => \N__30899\,
            I => \N__30872\
        );

    \I__6948\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30867\
        );

    \I__6947\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30867\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__30886\,
            I => \N__30864\
        );

    \I__6945\ : Span4Mux_v
    port map (
            O => \N__30883\,
            I => \N__30857\
        );

    \I__6944\ : Span4Mux_v
    port map (
            O => \N__30880\,
            I => \N__30857\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__30875\,
            I => \N__30857\
        );

    \I__6942\ : Odrv12
    port map (
            O => \N__30872\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__30867\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__30864\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6939\ : Odrv4
    port map (
            O => \N__30857\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6938\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30845\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__30845\,
            I => \POWERLED.d_i3_mux\
        );

    \I__6936\ : CascadeMux
    port map (
            O => \N__30842\,
            I => \POWERLED.func_state_RNI_5Z0Z_1_cascade_\
        );

    \I__6935\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30836\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__30836\,
            I => \N__30832\
        );

    \I__6933\ : InMux
    port map (
            O => \N__30835\,
            I => \N__30829\
        );

    \I__6932\ : Odrv4
    port map (
            O => \N__30832\,
            I => \POWERLED.N_23_i\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__30829\,
            I => \POWERLED.N_23_i\
        );

    \I__6930\ : InMux
    port map (
            O => \N__30824\,
            I => \N__30821\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__30821\,
            I => \N__30818\
        );

    \I__6928\ : Span4Mux_s2_h
    port map (
            O => \N__30818\,
            I => \N__30815\
        );

    \I__6927\ : Odrv4
    port map (
            O => \N__30815\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\
        );

    \I__6926\ : InMux
    port map (
            O => \N__30812\,
            I => \N__30806\
        );

    \I__6925\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30806\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__30806\,
            I => \POWERLED.N_85\
        );

    \I__6923\ : InMux
    port map (
            O => \N__30803\,
            I => \N__30800\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__30800\,
            I => \N__30796\
        );

    \I__6921\ : InMux
    port map (
            O => \N__30799\,
            I => \N__30793\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__30796\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_5\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__30793\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_5\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__30788\,
            I => \POWERLED.func_state_RNI12ASZ0Z_1_cascade_\
        );

    \I__6917\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30778\
        );

    \I__6916\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30775\
        );

    \I__6915\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30770\
        );

    \I__6914\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30770\
        );

    \I__6913\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30766\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30759\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__30775\,
            I => \N__30759\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__30770\,
            I => \N__30759\
        );

    \I__6909\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30756\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__30766\,
            I => \N__30751\
        );

    \I__6907\ : Span4Mux_s1_h
    port map (
            O => \N__30759\,
            I => \N__30751\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30748\
        );

    \I__6905\ : Span4Mux_h
    port map (
            O => \N__30751\,
            I => \N__30745\
        );

    \I__6904\ : Odrv12
    port map (
            O => \N__30748\,
            I => \POWERLED.N_613\
        );

    \I__6903\ : Odrv4
    port map (
            O => \N__30745\,
            I => \POWERLED.N_613\
        );

    \I__6902\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30729\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__30739\,
            I => \N__30724\
        );

    \I__6900\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30713\
        );

    \I__6899\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30713\
        );

    \I__6898\ : InMux
    port map (
            O => \N__30736\,
            I => \N__30713\
        );

    \I__6897\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30710\
        );

    \I__6896\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30700\
        );

    \I__6895\ : InMux
    port map (
            O => \N__30733\,
            I => \N__30700\
        );

    \I__6894\ : InMux
    port map (
            O => \N__30732\,
            I => \N__30697\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__30729\,
            I => \N__30691\
        );

    \I__6892\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30688\
        );

    \I__6891\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30684\
        );

    \I__6890\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30681\
        );

    \I__6889\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30676\
        );

    \I__6888\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30676\
        );

    \I__6887\ : CascadeMux
    port map (
            O => \N__30721\,
            I => \N__30673\
        );

    \I__6886\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30667\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__30713\,
            I => \N__30659\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__30710\,
            I => \N__30659\
        );

    \I__6883\ : InMux
    port map (
            O => \N__30709\,
            I => \N__30656\
        );

    \I__6882\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30647\
        );

    \I__6881\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30647\
        );

    \I__6880\ : InMux
    port map (
            O => \N__30706\,
            I => \N__30647\
        );

    \I__6879\ : InMux
    port map (
            O => \N__30705\,
            I => \N__30647\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__30700\,
            I => \N__30642\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__30697\,
            I => \N__30642\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30639\
        );

    \I__6875\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30634\
        );

    \I__6874\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30634\
        );

    \I__6873\ : Span4Mux_s0_h
    port map (
            O => \N__30691\,
            I => \N__30629\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__30688\,
            I => \N__30629\
        );

    \I__6871\ : InMux
    port map (
            O => \N__30687\,
            I => \N__30626\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__30684\,
            I => \N__30619\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__30681\,
            I => \N__30619\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30619\
        );

    \I__6867\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30612\
        );

    \I__6866\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30612\
        );

    \I__6865\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30612\
        );

    \I__6864\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30609\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__30667\,
            I => \N__30606\
        );

    \I__6862\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30603\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__30665\,
            I => \N__30599\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__30664\,
            I => \N__30595\
        );

    \I__6859\ : Span4Mux_v
    port map (
            O => \N__30659\,
            I => \N__30588\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__30656\,
            I => \N__30588\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__30647\,
            I => \N__30588\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__30642\,
            I => \N__30581\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30581\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__30634\,
            I => \N__30581\
        );

    \I__6853\ : Span4Mux_v
    port map (
            O => \N__30629\,
            I => \N__30572\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__30626\,
            I => \N__30569\
        );

    \I__6851\ : Span4Mux_v
    port map (
            O => \N__30619\,
            I => \N__30564\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__30612\,
            I => \N__30564\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__30609\,
            I => \N__30557\
        );

    \I__6848\ : Span4Mux_v
    port map (
            O => \N__30606\,
            I => \N__30557\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__30603\,
            I => \N__30557\
        );

    \I__6846\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30554\
        );

    \I__6845\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30551\
        );

    \I__6844\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30545\
        );

    \I__6843\ : InMux
    port map (
            O => \N__30595\,
            I => \N__30545\
        );

    \I__6842\ : Span4Mux_v
    port map (
            O => \N__30588\,
            I => \N__30540\
        );

    \I__6841\ : Span4Mux_v
    port map (
            O => \N__30581\,
            I => \N__30540\
        );

    \I__6840\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30533\
        );

    \I__6839\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30533\
        );

    \I__6838\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30533\
        );

    \I__6837\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30526\
        );

    \I__6836\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30526\
        );

    \I__6835\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30526\
        );

    \I__6834\ : Span4Mux_v
    port map (
            O => \N__30572\,
            I => \N__30521\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__30569\,
            I => \N__30521\
        );

    \I__6832\ : Span4Mux_v
    port map (
            O => \N__30564\,
            I => \N__30514\
        );

    \I__6831\ : Span4Mux_h
    port map (
            O => \N__30557\,
            I => \N__30514\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__30554\,
            I => \N__30514\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__30551\,
            I => \N__30511\
        );

    \I__6828\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30508\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__30545\,
            I => \N__30501\
        );

    \I__6826\ : Sp12to4
    port map (
            O => \N__30540\,
            I => \N__30501\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__30533\,
            I => \N__30501\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__30526\,
            I => \N__30498\
        );

    \I__6823\ : Span4Mux_h
    port map (
            O => \N__30521\,
            I => \N__30493\
        );

    \I__6822\ : Span4Mux_v
    port map (
            O => \N__30514\,
            I => \N__30493\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__30511\,
            I => \N__30488\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__30508\,
            I => \N__30488\
        );

    \I__6819\ : Span12Mux_s8_h
    port map (
            O => \N__30501\,
            I => \N__30485\
        );

    \I__6818\ : Span12Mux_s8_h
    port map (
            O => \N__30498\,
            I => \N__30482\
        );

    \I__6817\ : IoSpan4Mux
    port map (
            O => \N__30493\,
            I => \N__30477\
        );

    \I__6816\ : IoSpan4Mux
    port map (
            O => \N__30488\,
            I => \N__30477\
        );

    \I__6815\ : Odrv12
    port map (
            O => \N__30485\,
            I => slp_s4n
        );

    \I__6814\ : Odrv12
    port map (
            O => \N__30482\,
            I => slp_s4n
        );

    \I__6813\ : Odrv4
    port map (
            O => \N__30477\,
            I => slp_s4n
        );

    \I__6812\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30464\
        );

    \I__6811\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30464\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__30464\,
            I => \N__30461\
        );

    \I__6809\ : Span4Mux_v
    port map (
            O => \N__30461\,
            I => \N__30458\
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__30458\,
            I => \POWERLED.func_state_RNI8AQHZ0Z_0\
        );

    \I__6807\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30452\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__30452\,
            I => \N__30449\
        );

    \I__6805\ : Span12Mux_s6_v
    port map (
            O => \N__30449\,
            I => \N__30446\
        );

    \I__6804\ : Odrv12
    port map (
            O => \N__30446\,
            I => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\
        );

    \I__6803\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30437\
        );

    \I__6802\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30437\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__30437\,
            I => \POWERLED.func_state_RNI12ASZ0Z_1\
        );

    \I__6800\ : InMux
    port map (
            O => \N__30434\,
            I => \N__30428\
        );

    \I__6799\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30428\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__30428\,
            I => \N__30425\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__30425\,
            I => \POWERLED.N_83\
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__30422\,
            I => \N__30417\
        );

    \I__6795\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30402\
        );

    \I__6794\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30402\
        );

    \I__6793\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30402\
        );

    \I__6792\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30395\
        );

    \I__6791\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30395\
        );

    \I__6790\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30395\
        );

    \I__6789\ : InMux
    port map (
            O => \N__30413\,
            I => \N__30390\
        );

    \I__6788\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30390\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__30411\,
            I => \N__30384\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__30410\,
            I => \N__30381\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__30409\,
            I => \N__30378\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30374\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__30395\,
            I => \N__30369\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__30390\,
            I => \N__30369\
        );

    \I__6781\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30364\
        );

    \I__6780\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30364\
        );

    \I__6779\ : InMux
    port map (
            O => \N__30387\,
            I => \N__30355\
        );

    \I__6778\ : InMux
    port map (
            O => \N__30384\,
            I => \N__30355\
        );

    \I__6777\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30355\
        );

    \I__6776\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30355\
        );

    \I__6775\ : CascadeMux
    port map (
            O => \N__30377\,
            I => \N__30349\
        );

    \I__6774\ : Span4Mux_h
    port map (
            O => \N__30374\,
            I => \N__30337\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__30369\,
            I => \N__30337\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__30364\,
            I => \N__30337\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__30355\,
            I => \N__30337\
        );

    \I__6770\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30332\
        );

    \I__6769\ : InMux
    port map (
            O => \N__30353\,
            I => \N__30332\
        );

    \I__6768\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30325\
        );

    \I__6767\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30325\
        );

    \I__6766\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30325\
        );

    \I__6765\ : CascadeMux
    port map (
            O => \N__30347\,
            I => \N__30322\
        );

    \I__6764\ : CascadeMux
    port map (
            O => \N__30346\,
            I => \N__30319\
        );

    \I__6763\ : Span4Mux_v
    port map (
            O => \N__30337\,
            I => \N__30311\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__30332\,
            I => \N__30306\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30325\,
            I => \N__30306\
        );

    \I__6760\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30299\
        );

    \I__6759\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30299\
        );

    \I__6758\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30299\
        );

    \I__6757\ : InMux
    port map (
            O => \N__30317\,
            I => \N__30296\
        );

    \I__6756\ : CascadeMux
    port map (
            O => \N__30316\,
            I => \N__30293\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__30315\,
            I => \N__30290\
        );

    \I__6754\ : CascadeMux
    port map (
            O => \N__30314\,
            I => \N__30285\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__30311\,
            I => \N__30281\
        );

    \I__6752\ : Span4Mux_v
    port map (
            O => \N__30306\,
            I => \N__30274\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__30299\,
            I => \N__30274\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__30296\,
            I => \N__30274\
        );

    \I__6749\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30267\
        );

    \I__6748\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30267\
        );

    \I__6747\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30267\
        );

    \I__6746\ : InMux
    port map (
            O => \N__30288\,
            I => \N__30259\
        );

    \I__6745\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30259\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__30284\,
            I => \N__30255\
        );

    \I__6743\ : IoSpan4Mux
    port map (
            O => \N__30281\,
            I => \N__30248\
        );

    \I__6742\ : Span4Mux_v
    port map (
            O => \N__30274\,
            I => \N__30248\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30248\
        );

    \I__6740\ : InMux
    port map (
            O => \N__30266\,
            I => \N__30245\
        );

    \I__6739\ : CascadeMux
    port map (
            O => \N__30265\,
            I => \N__30240\
        );

    \I__6738\ : CascadeMux
    port map (
            O => \N__30264\,
            I => \N__30236\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__30259\,
            I => \N__30232\
        );

    \I__6736\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30229\
        );

    \I__6735\ : InMux
    port map (
            O => \N__30255\,
            I => \N__30224\
        );

    \I__6734\ : IoSpan4Mux
    port map (
            O => \N__30248\,
            I => \N__30221\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__30245\,
            I => \N__30218\
        );

    \I__6732\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30213\
        );

    \I__6731\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30213\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30208\
        );

    \I__6729\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30208\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30205\
        );

    \I__6727\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30202\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__30232\,
            I => \N__30197\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30229\,
            I => \N__30197\
        );

    \I__6724\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30192\
        );

    \I__6723\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30192\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__30224\,
            I => \N__30189\
        );

    \I__6721\ : IoSpan4Mux
    port map (
            O => \N__30221\,
            I => \N__30186\
        );

    \I__6720\ : Span12Mux_s10_h
    port map (
            O => \N__30218\,
            I => \N__30177\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__30213\,
            I => \N__30177\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__30208\,
            I => \N__30177\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__30205\,
            I => \N__30177\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30202\,
            I => \N__30174\
        );

    \I__6715\ : Span4Mux_v
    port map (
            O => \N__30197\,
            I => \N__30169\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__30192\,
            I => \N__30169\
        );

    \I__6713\ : Odrv12
    port map (
            O => \N__30189\,
            I => slp_s3n
        );

    \I__6712\ : Odrv4
    port map (
            O => \N__30186\,
            I => slp_s3n
        );

    \I__6711\ : Odrv12
    port map (
            O => \N__30177\,
            I => slp_s3n
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__30174\,
            I => slp_s3n
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__30169\,
            I => slp_s3n
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__30158\,
            I => \N__30154\
        );

    \I__6707\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30134\
        );

    \I__6706\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30134\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30134\
        );

    \I__6704\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30134\
        );

    \I__6703\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30129\
        );

    \I__6702\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30129\
        );

    \I__6701\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30126\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__30148\,
            I => \N__30119\
        );

    \I__6699\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30112\
        );

    \I__6698\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30109\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__30145\,
            I => \N__30106\
        );

    \I__6696\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30102\
        );

    \I__6695\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30099\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30096\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__30129\,
            I => \N__30091\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__30126\,
            I => \N__30091\
        );

    \I__6691\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30086\
        );

    \I__6690\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30086\
        );

    \I__6689\ : InMux
    port map (
            O => \N__30123\,
            I => \N__30083\
        );

    \I__6688\ : InMux
    port map (
            O => \N__30122\,
            I => \N__30080\
        );

    \I__6687\ : InMux
    port map (
            O => \N__30119\,
            I => \N__30076\
        );

    \I__6686\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30070\
        );

    \I__6685\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30065\
        );

    \I__6684\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30065\
        );

    \I__6683\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30062\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30058\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__30109\,
            I => \N__30055\
        );

    \I__6680\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30050\
        );

    \I__6679\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30050\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30046\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__30099\,
            I => \N__30037\
        );

    \I__6676\ : Span4Mux_v
    port map (
            O => \N__30096\,
            I => \N__30037\
        );

    \I__6675\ : Span4Mux_s3_v
    port map (
            O => \N__30091\,
            I => \N__30037\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__30086\,
            I => \N__30037\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__30083\,
            I => \N__30032\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__30080\,
            I => \N__30032\
        );

    \I__6671\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30029\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__30076\,
            I => \N__30026\
        );

    \I__6669\ : InMux
    port map (
            O => \N__30075\,
            I => \N__30023\
        );

    \I__6668\ : CascadeMux
    port map (
            O => \N__30074\,
            I => \N__30019\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30015\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__30070\,
            I => \N__30005\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__30065\,
            I => \N__30005\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__30062\,
            I => \N__30005\
        );

    \I__6663\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30002\
        );

    \I__6662\ : Span4Mux_s2_h
    port map (
            O => \N__30058\,
            I => \N__29997\
        );

    \I__6661\ : Span4Mux_s2_h
    port map (
            O => \N__30055\,
            I => \N__29997\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__30050\,
            I => \N__29994\
        );

    \I__6659\ : InMux
    port map (
            O => \N__30049\,
            I => \N__29991\
        );

    \I__6658\ : Span4Mux_v
    port map (
            O => \N__30046\,
            I => \N__29982\
        );

    \I__6657\ : Span4Mux_v
    port map (
            O => \N__30037\,
            I => \N__29982\
        );

    \I__6656\ : Span4Mux_v
    port map (
            O => \N__30032\,
            I => \N__29982\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__30029\,
            I => \N__29982\
        );

    \I__6654\ : Span12Mux_s5_h
    port map (
            O => \N__30026\,
            I => \N__29977\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__30023\,
            I => \N__29974\
        );

    \I__6652\ : InMux
    port map (
            O => \N__30022\,
            I => \N__29969\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30019\,
            I => \N__29969\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30018\,
            I => \N__29966\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__30015\,
            I => \N__29963\
        );

    \I__6648\ : InMux
    port map (
            O => \N__30014\,
            I => \N__29960\
        );

    \I__6647\ : InMux
    port map (
            O => \N__30013\,
            I => \N__29955\
        );

    \I__6646\ : InMux
    port map (
            O => \N__30012\,
            I => \N__29955\
        );

    \I__6645\ : Span4Mux_v
    port map (
            O => \N__30005\,
            I => \N__29946\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29946\
        );

    \I__6643\ : Span4Mux_v
    port map (
            O => \N__29997\,
            I => \N__29946\
        );

    \I__6642\ : Span4Mux_s2_h
    port map (
            O => \N__29994\,
            I => \N__29946\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__29991\,
            I => \N__29941\
        );

    \I__6640\ : Span4Mux_h
    port map (
            O => \N__29982\,
            I => \N__29941\
        );

    \I__6639\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29936\
        );

    \I__6638\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29936\
        );

    \I__6637\ : Odrv12
    port map (
            O => \N__29977\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__29974\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__29969\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__29966\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__29963\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__29960\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__29955\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__29946\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6629\ : Odrv4
    port map (
            O => \N__29941\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__29936\,
            I => \func_state_RNIMJ6IF_0_1\
        );

    \I__6627\ : InMux
    port map (
            O => \N__29915\,
            I => \N__29909\
        );

    \I__6626\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29904\
        );

    \I__6625\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29904\
        );

    \I__6624\ : CascadeMux
    port map (
            O => \N__29912\,
            I => \N__29901\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__29909\,
            I => \N__29889\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__29904\,
            I => \N__29886\
        );

    \I__6621\ : InMux
    port map (
            O => \N__29901\,
            I => \N__29881\
        );

    \I__6620\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29881\
        );

    \I__6619\ : InMux
    port map (
            O => \N__29899\,
            I => \N__29876\
        );

    \I__6618\ : InMux
    port map (
            O => \N__29898\,
            I => \N__29876\
        );

    \I__6617\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29869\
        );

    \I__6616\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29869\
        );

    \I__6615\ : InMux
    port map (
            O => \N__29895\,
            I => \N__29869\
        );

    \I__6614\ : InMux
    port map (
            O => \N__29894\,
            I => \N__29866\
        );

    \I__6613\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29863\
        );

    \I__6612\ : InMux
    port map (
            O => \N__29892\,
            I => \N__29859\
        );

    \I__6611\ : Span4Mux_s3_v
    port map (
            O => \N__29889\,
            I => \N__29848\
        );

    \I__6610\ : Span4Mux_h
    port map (
            O => \N__29886\,
            I => \N__29848\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29848\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29848\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__29869\,
            I => \N__29848\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29845\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29841\
        );

    \I__6604\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29838\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__29859\,
            I => \N__29833\
        );

    \I__6602\ : Span4Mux_v
    port map (
            O => \N__29848\,
            I => \N__29833\
        );

    \I__6601\ : Span12Mux_s4_v
    port map (
            O => \N__29845\,
            I => \N__29830\
        );

    \I__6600\ : InMux
    port map (
            O => \N__29844\,
            I => \N__29827\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__29841\,
            I => \N__29820\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N__29820\
        );

    \I__6597\ : Span4Mux_h
    port map (
            O => \N__29833\,
            I => \N__29820\
        );

    \I__6596\ : Odrv12
    port map (
            O => \N__29830\,
            I => \RSMRSTn_rep2\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__29827\,
            I => \RSMRSTn_rep2\
        );

    \I__6594\ : Odrv4
    port map (
            O => \N__29820\,
            I => \RSMRSTn_rep2\
        );

    \I__6593\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29809\
        );

    \I__6592\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29806\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__29809\,
            I => \N__29802\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29799\
        );

    \I__6589\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29796\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__29802\,
            I => \POWERLED.N_531\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__29799\,
            I => \POWERLED.N_531\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__29796\,
            I => \POWERLED.N_531\
        );

    \I__6585\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29786\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__29786\,
            I => \N__29783\
        );

    \I__6583\ : Span4Mux_v
    port map (
            O => \N__29783\,
            I => \N__29780\
        );

    \I__6582\ : Sp12to4
    port map (
            O => \N__29780\,
            I => \N__29777\
        );

    \I__6581\ : Span12Mux_s3_h
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__6580\ : Odrv12
    port map (
            O => \N__29774\,
            I => \POWERLED.un1_clk_100khz_51_and_i_3_0\
        );

    \I__6579\ : CascadeMux
    port map (
            O => \N__29771\,
            I => \POWERLED.N_532_cascade_\
        );

    \I__6578\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29765\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__29765\,
            I => \POWERLED.N_530\
        );

    \I__6576\ : CascadeMux
    port map (
            O => \N__29762\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_5_cascade_\
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__29759\,
            I => \N__29754\
        );

    \I__6574\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29749\
        );

    \I__6573\ : InMux
    port map (
            O => \N__29757\,
            I => \N__29749\
        );

    \I__6572\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29745\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__29749\,
            I => \N__29739\
        );

    \I__6570\ : InMux
    port map (
            O => \N__29748\,
            I => \N__29736\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__29745\,
            I => \N__29733\
        );

    \I__6568\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29730\
        );

    \I__6567\ : CascadeMux
    port map (
            O => \N__29743\,
            I => \N__29727\
        );

    \I__6566\ : CascadeMux
    port map (
            O => \N__29742\,
            I => \N__29722\
        );

    \I__6565\ : Span4Mux_s3_v
    port map (
            O => \N__29739\,
            I => \N__29717\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__29736\,
            I => \N__29717\
        );

    \I__6563\ : Span4Mux_s3_v
    port map (
            O => \N__29733\,
            I => \N__29712\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__29730\,
            I => \N__29712\
        );

    \I__6561\ : InMux
    port map (
            O => \N__29727\,
            I => \N__29709\
        );

    \I__6560\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29706\
        );

    \I__6559\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29703\
        );

    \I__6558\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29700\
        );

    \I__6557\ : Span4Mux_v
    port map (
            O => \N__29717\,
            I => \N__29694\
        );

    \I__6556\ : Span4Mux_v
    port map (
            O => \N__29712\,
            I => \N__29694\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__29709\,
            I => \N__29691\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__29706\,
            I => \N__29688\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__29703\,
            I => \N__29683\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__29700\,
            I => \N__29683\
        );

    \I__6551\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29680\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__29694\,
            I => \POWERLED.N_251\
        );

    \I__6549\ : Odrv4
    port map (
            O => \N__29691\,
            I => \POWERLED.N_251\
        );

    \I__6548\ : Odrv12
    port map (
            O => \N__29688\,
            I => \POWERLED.N_251\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__29683\,
            I => \POWERLED.N_251\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__29680\,
            I => \POWERLED.N_251\
        );

    \I__6545\ : InMux
    port map (
            O => \N__29669\,
            I => \N__29665\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__29668\,
            I => \N__29662\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__29665\,
            I => \N__29659\
        );

    \I__6542\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29656\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__29659\,
            I => \N__29651\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__29656\,
            I => \N__29648\
        );

    \I__6539\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29645\
        );

    \I__6538\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29642\
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__29651\,
            I => \POWERLED.N_633\
        );

    \I__6536\ : Odrv4
    port map (
            O => \N__29648\,
            I => \POWERLED.N_633\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__29645\,
            I => \POWERLED.N_633\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__29642\,
            I => \POWERLED.N_633\
        );

    \I__6533\ : CascadeMux
    port map (
            O => \N__29633\,
            I => \POWERLED.func_state_RNIOGRSZ0Z_1_cascade_\
        );

    \I__6532\ : IoInMux
    port map (
            O => \N__29630\,
            I => \N__29627\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__29627\,
            I => \N__29623\
        );

    \I__6530\ : IoInMux
    port map (
            O => \N__29626\,
            I => \N__29620\
        );

    \I__6529\ : IoSpan4Mux
    port map (
            O => \N__29623\,
            I => \N__29614\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__29620\,
            I => \N__29611\
        );

    \I__6527\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29605\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__29618\,
            I => \N__29601\
        );

    \I__6525\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29597\
        );

    \I__6524\ : Span4Mux_s0_h
    port map (
            O => \N__29614\,
            I => \N__29594\
        );

    \I__6523\ : Span4Mux_s0_h
    port map (
            O => \N__29611\,
            I => \N__29591\
        );

    \I__6522\ : InMux
    port map (
            O => \N__29610\,
            I => \N__29586\
        );

    \I__6521\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29586\
        );

    \I__6520\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29583\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__29605\,
            I => \N__29580\
        );

    \I__6518\ : InMux
    port map (
            O => \N__29604\,
            I => \N__29577\
        );

    \I__6517\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29574\
        );

    \I__6516\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29569\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__29597\,
            I => \N__29566\
        );

    \I__6514\ : Sp12to4
    port map (
            O => \N__29594\,
            I => \N__29559\
        );

    \I__6513\ : Sp12to4
    port map (
            O => \N__29591\,
            I => \N__29559\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__29586\,
            I => \N__29559\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__29583\,
            I => \N__29554\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__29580\,
            I => \N__29547\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__29577\,
            I => \N__29547\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__29574\,
            I => \N__29547\
        );

    \I__6507\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29544\
        );

    \I__6506\ : InMux
    port map (
            O => \N__29572\,
            I => \N__29541\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__29569\,
            I => \N__29538\
        );

    \I__6504\ : Span4Mux_h
    port map (
            O => \N__29566\,
            I => \N__29533\
        );

    \I__6503\ : Span12Mux_s10_v
    port map (
            O => \N__29559\,
            I => \N__29530\
        );

    \I__6502\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29527\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29524\
        );

    \I__6500\ : Span4Mux_v
    port map (
            O => \N__29554\,
            I => \N__29521\
        );

    \I__6499\ : Span4Mux_v
    port map (
            O => \N__29547\,
            I => \N__29518\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__29544\,
            I => \N__29511\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29511\
        );

    \I__6496\ : Span4Mux_s3_h
    port map (
            O => \N__29538\,
            I => \N__29511\
        );

    \I__6495\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29506\
        );

    \I__6494\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29506\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__29533\,
            I => v5s_enn
        );

    \I__6492\ : Odrv12
    port map (
            O => \N__29530\,
            I => v5s_enn
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__29527\,
            I => v5s_enn
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__29524\,
            I => v5s_enn
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__29521\,
            I => v5s_enn
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__29518\,
            I => v5s_enn
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__29511\,
            I => v5s_enn
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__29506\,
            I => v5s_enn
        );

    \I__6485\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29486\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__29486\,
            I => \N__29481\
        );

    \I__6483\ : InMux
    port map (
            O => \N__29485\,
            I => \N__29476\
        );

    \I__6482\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29476\
        );

    \I__6481\ : Odrv12
    port map (
            O => \N__29481\,
            I => \POWERLED.N_413_N\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__29476\,
            I => \POWERLED.N_413_N\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__29471\,
            I => \N__29467\
        );

    \I__6478\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29462\
        );

    \I__6477\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29462\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__29462\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__6475\ : CascadeMux
    port map (
            O => \N__29459\,
            I => \POWERLED.dutycycleZ0Z_6_cascade_\
        );

    \I__6474\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29452\
        );

    \I__6473\ : InMux
    port map (
            O => \N__29455\,
            I => \N__29449\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__29452\,
            I => \N__29446\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__29449\,
            I => \N__29443\
        );

    \I__6470\ : Span4Mux_v
    port map (
            O => \N__29446\,
            I => \N__29437\
        );

    \I__6469\ : Span4Mux_s1_h
    port map (
            O => \N__29443\,
            I => \N__29437\
        );

    \I__6468\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29434\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__29437\,
            I => \N__29429\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__29434\,
            I => \N__29429\
        );

    \I__6465\ : Span4Mux_v
    port map (
            O => \N__29429\,
            I => \N__29426\
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__29426\,
            I => \POWERLED.N_612\
        );

    \I__6463\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29420\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29417\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__29417\,
            I => \N__29414\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__29414\,
            I => \POWERLED.N_672\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__29411\,
            I => \POWERLED.N_672_cascade_\
        );

    \I__6458\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29405\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__29405\,
            I => \N__29402\
        );

    \I__6456\ : Span4Mux_h
    port map (
            O => \N__29402\,
            I => \N__29399\
        );

    \I__6455\ : Odrv4
    port map (
            O => \N__29399\,
            I => \POWERLED.un1_dutycycle_168_0\
        );

    \I__6454\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29390\
        );

    \I__6453\ : InMux
    port map (
            O => \N__29395\,
            I => \N__29390\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__29390\,
            I => \N__29385\
        );

    \I__6451\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29380\
        );

    \I__6450\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29380\
        );

    \I__6449\ : Span4Mux_v
    port map (
            O => \N__29385\,
            I => \N__29377\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__29380\,
            I => \N__29374\
        );

    \I__6447\ : Odrv4
    port map (
            O => \N__29377\,
            I => \POWERLED.count_clk_RNIZ0Z_6\
        );

    \I__6446\ : Odrv12
    port map (
            O => \N__29374\,
            I => \POWERLED.count_clk_RNIZ0Z_6\
        );

    \I__6445\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29366\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29361\
        );

    \I__6443\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29356\
        );

    \I__6442\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29356\
        );

    \I__6441\ : Span4Mux_v
    port map (
            O => \N__29361\,
            I => \N__29352\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__29356\,
            I => \N__29349\
        );

    \I__6439\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29346\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__29352\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__29349\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__29346\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__29339\,
            I => \POWERLED.N_412_i_cascade_\
        );

    \I__6434\ : InMux
    port map (
            O => \N__29336\,
            I => \N__29332\
        );

    \I__6433\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29329\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29332\,
            I => \N__29326\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__29329\,
            I => \N__29323\
        );

    \I__6430\ : Span4Mux_v
    port map (
            O => \N__29326\,
            I => \N__29320\
        );

    \I__6429\ : Span4Mux_s2_v
    port map (
            O => \N__29323\,
            I => \N__29317\
        );

    \I__6428\ : Odrv4
    port map (
            O => \N__29320\,
            I => \POWERLED.N_604\
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__29317\,
            I => \POWERLED.N_604\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__29312\,
            I => \N__29309\
        );

    \I__6425\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29303\
        );

    \I__6424\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29303\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__29303\,
            I => \N__29300\
        );

    \I__6422\ : Span12Mux_s9_v
    port map (
            O => \N__29300\,
            I => \N__29297\
        );

    \I__6421\ : Odrv12
    port map (
            O => \N__29297\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_3\
        );

    \I__6420\ : CascadeMux
    port map (
            O => \N__29294\,
            I => \N__29288\
        );

    \I__6419\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29285\
        );

    \I__6418\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29282\
        );

    \I__6417\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29279\
        );

    \I__6416\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29276\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29271\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__29282\,
            I => \N__29268\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29264\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__29276\,
            I => \N__29261\
        );

    \I__6411\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29256\
        );

    \I__6410\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29256\
        );

    \I__6409\ : Span4Mux_s3_h
    port map (
            O => \N__29271\,
            I => \N__29253\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__29268\,
            I => \N__29250\
        );

    \I__6407\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29247\
        );

    \I__6406\ : Span4Mux_s3_h
    port map (
            O => \N__29264\,
            I => \N__29240\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__29261\,
            I => \N__29240\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29240\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__29253\,
            I => \POWERLED.N_435\
        );

    \I__6402\ : Odrv4
    port map (
            O => \N__29250\,
            I => \POWERLED.N_435\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__29247\,
            I => \POWERLED.N_435\
        );

    \I__6400\ : Odrv4
    port map (
            O => \N__29240\,
            I => \POWERLED.N_435\
        );

    \I__6399\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29227\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__29230\,
            I => \N__29224\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__29227\,
            I => \N__29219\
        );

    \I__6396\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29216\
        );

    \I__6395\ : CascadeMux
    port map (
            O => \N__29223\,
            I => \N__29213\
        );

    \I__6394\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29210\
        );

    \I__6393\ : Span4Mux_v
    port map (
            O => \N__29219\,
            I => \N__29206\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__29216\,
            I => \N__29203\
        );

    \I__6391\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29200\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29197\
        );

    \I__6389\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29194\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__29206\,
            I => \N__29187\
        );

    \I__6387\ : Span4Mux_h
    port map (
            O => \N__29203\,
            I => \N__29187\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29187\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__29197\,
            I => \POWERLED.N_412_i\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__29194\,
            I => \POWERLED.N_412_i\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__29187\,
            I => \POWERLED.N_412_i\
        );

    \I__6382\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29177\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29174\
        );

    \I__6380\ : Span4Mux_h
    port map (
            O => \N__29174\,
            I => \N__29170\
        );

    \I__6379\ : InMux
    port map (
            O => \N__29173\,
            I => \N__29167\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__29170\,
            I => \POWERLED.func_state_RNI_5Z0Z_1\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__29167\,
            I => \POWERLED.func_state_RNI_5Z0Z_1\
        );

    \I__6376\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29156\
        );

    \I__6375\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29156\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__6373\ : Odrv4
    port map (
            O => \N__29153\,
            I => \POWERLED.count_clk_1_13\
        );

    \I__6372\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29147\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__29147\,
            I => \POWERLED.count_clk_0_13\
        );

    \I__6370\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29138\
        );

    \I__6368\ : Odrv12
    port map (
            O => \N__29138\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__6367\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29126\
        );

    \I__6366\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29126\
        );

    \I__6365\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29126\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__29126\,
            I => \N__29123\
        );

    \I__6363\ : Odrv4
    port map (
            O => \N__29123\,
            I => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\
        );

    \I__6362\ : CascadeMux
    port map (
            O => \N__29120\,
            I => \N__29114\
        );

    \I__6361\ : CascadeMux
    port map (
            O => \N__29119\,
            I => \N__29111\
        );

    \I__6360\ : CEMux
    port map (
            O => \N__29118\,
            I => \N__29107\
        );

    \I__6359\ : CEMux
    port map (
            O => \N__29117\,
            I => \N__29100\
        );

    \I__6358\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29092\
        );

    \I__6357\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29092\
        );

    \I__6356\ : CEMux
    port map (
            O => \N__29110\,
            I => \N__29092\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__29107\,
            I => \N__29089\
        );

    \I__6354\ : CEMux
    port map (
            O => \N__29106\,
            I => \N__29086\
        );

    \I__6353\ : CascadeMux
    port map (
            O => \N__29105\,
            I => \N__29083\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__29104\,
            I => \N__29077\
        );

    \I__6351\ : CEMux
    port map (
            O => \N__29103\,
            I => \N__29071\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__29100\,
            I => \N__29066\
        );

    \I__6349\ : InMux
    port map (
            O => \N__29099\,
            I => \N__29063\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__29092\,
            I => \N__29057\
        );

    \I__6347\ : Span4Mux_v
    port map (
            O => \N__29089\,
            I => \N__29052\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__29086\,
            I => \N__29052\
        );

    \I__6345\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29047\
        );

    \I__6344\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29047\
        );

    \I__6343\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29040\
        );

    \I__6342\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29040\
        );

    \I__6341\ : InMux
    port map (
            O => \N__29077\,
            I => \N__29040\
        );

    \I__6340\ : CEMux
    port map (
            O => \N__29076\,
            I => \N__29034\
        );

    \I__6339\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29031\
        );

    \I__6338\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29028\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29025\
        );

    \I__6336\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29020\
        );

    \I__6335\ : CEMux
    port map (
            O => \N__29069\,
            I => \N__29020\
        );

    \I__6334\ : Span4Mux_v
    port map (
            O => \N__29066\,
            I => \N__29017\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29014\
        );

    \I__6332\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29007\
        );

    \I__6331\ : InMux
    port map (
            O => \N__29061\,
            I => \N__29007\
        );

    \I__6330\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29007\
        );

    \I__6329\ : Span4Mux_v
    port map (
            O => \N__29057\,
            I => \N__29000\
        );

    \I__6328\ : Span4Mux_s3_v
    port map (
            O => \N__29052\,
            I => \N__29000\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__29047\,
            I => \N__29000\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__29040\,
            I => \N__28997\
        );

    \I__6325\ : InMux
    port map (
            O => \N__29039\,
            I => \N__28992\
        );

    \I__6324\ : InMux
    port map (
            O => \N__29038\,
            I => \N__28992\
        );

    \I__6323\ : InMux
    port map (
            O => \N__29037\,
            I => \N__28987\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__29034\,
            I => \N__28984\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__29031\,
            I => \N__28977\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__29028\,
            I => \N__28977\
        );

    \I__6319\ : Span4Mux_h
    port map (
            O => \N__29025\,
            I => \N__28977\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__29020\,
            I => \N__28970\
        );

    \I__6317\ : Span4Mux_h
    port map (
            O => \N__29017\,
            I => \N__28970\
        );

    \I__6316\ : Span4Mux_v
    port map (
            O => \N__29014\,
            I => \N__28970\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__29007\,
            I => \N__28961\
        );

    \I__6314\ : Span4Mux_s0_h
    port map (
            O => \N__29000\,
            I => \N__28961\
        );

    \I__6313\ : Span4Mux_s3_v
    port map (
            O => \N__28997\,
            I => \N__28961\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__28992\,
            I => \N__28961\
        );

    \I__6311\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28956\
        );

    \I__6310\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28956\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__28987\,
            I => \POWERLED.count_clk_en\
        );

    \I__6308\ : Odrv12
    port map (
            O => \N__28984\,
            I => \POWERLED.count_clk_en\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__28977\,
            I => \POWERLED.count_clk_en\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__28970\,
            I => \POWERLED.count_clk_en\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__28961\,
            I => \POWERLED.count_clk_en\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__28956\,
            I => \POWERLED.count_clk_en\
        );

    \I__6303\ : CascadeMux
    port map (
            O => \N__28943\,
            I => \POWERLED.count_clkZ0Z_13_cascade_\
        );

    \I__6302\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28934\
        );

    \I__6301\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28934\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__28934\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__6299\ : InMux
    port map (
            O => \N__28931\,
            I => \N__28928\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__28928\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_0\
        );

    \I__6297\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28920\
        );

    \I__6296\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28915\
        );

    \I__6295\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28915\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__28920\,
            I => \N__28912\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__28915\,
            I => \N__28909\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__28912\,
            I => \N__28905\
        );

    \I__6291\ : Span4Mux_v
    port map (
            O => \N__28909\,
            I => \N__28902\
        );

    \I__6290\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28899\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__28905\,
            I => \POWERLED.N_676\
        );

    \I__6288\ : Odrv4
    port map (
            O => \N__28902\,
            I => \POWERLED.N_676\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__28899\,
            I => \POWERLED.N_676\
        );

    \I__6286\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28889\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__28889\,
            I => \POWERLED.N_492\
        );

    \I__6284\ : CascadeMux
    port map (
            O => \N__28886\,
            I => \N__28882\
        );

    \I__6283\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28877\
        );

    \I__6282\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28877\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__28877\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__6280\ : InMux
    port map (
            O => \N__28874\,
            I => \N__28868\
        );

    \I__6279\ : InMux
    port map (
            O => \N__28873\,
            I => \N__28868\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__28868\,
            I => \N__28865\
        );

    \I__6277\ : Span4Mux_s2_h
    port map (
            O => \N__28865\,
            I => \N__28862\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__28862\,
            I => \POWERLED.func_state_RNIS28SBZ0Z_1\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__28859\,
            I => \POWERLED.dutycycleZ1Z_5_cascade_\
        );

    \I__6274\ : CascadeMux
    port map (
            O => \N__28856\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_5_cascade_\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__28853\,
            I => \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_a2_0_cascade_\
        );

    \I__6272\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28836\
        );

    \I__6271\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28836\
        );

    \I__6270\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28833\
        );

    \I__6269\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28829\
        );

    \I__6268\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28824\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28845\,
            I => \N__28824\
        );

    \I__6266\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28817\
        );

    \I__6265\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28817\
        );

    \I__6264\ : InMux
    port map (
            O => \N__28842\,
            I => \N__28817\
        );

    \I__6263\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28810\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__28836\,
            I => \N__28805\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__28833\,
            I => \N__28805\
        );

    \I__6260\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28802\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__28829\,
            I => \N__28797\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28792\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__28817\,
            I => \N__28792\
        );

    \I__6256\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28787\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28782\
        );

    \I__6254\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28782\
        );

    \I__6253\ : InMux
    port map (
            O => \N__28813\,
            I => \N__28779\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__28810\,
            I => \N__28772\
        );

    \I__6251\ : Span4Mux_s3_h
    port map (
            O => \N__28805\,
            I => \N__28772\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28772\
        );

    \I__6249\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28767\
        );

    \I__6248\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28767\
        );

    \I__6247\ : Span4Mux_v
    port map (
            O => \N__28797\,
            I => \N__28762\
        );

    \I__6246\ : Span4Mux_v
    port map (
            O => \N__28792\,
            I => \N__28762\
        );

    \I__6245\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28757\
        );

    \I__6244\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28757\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__28787\,
            I => \N__28754\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__28782\,
            I => \func_state_RNI_2_0\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__28779\,
            I => \func_state_RNI_2_0\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__28772\,
            I => \func_state_RNI_2_0\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__28767\,
            I => \func_state_RNI_2_0\
        );

    \I__6238\ : Odrv4
    port map (
            O => \N__28762\,
            I => \func_state_RNI_2_0\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__28757\,
            I => \func_state_RNI_2_0\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__28754\,
            I => \func_state_RNI_2_0\
        );

    \I__6235\ : InMux
    port map (
            O => \N__28739\,
            I => \N__28736\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__28736\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_ns_1\
        );

    \I__6233\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28730\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__28730\,
            I => \POWERLED.count_clk_0_0\
        );

    \I__6231\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28724\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__28724\,
            I => \POWERLED.count_clk_RNI_0Z0Z_0\
        );

    \I__6229\ : InMux
    port map (
            O => \N__28721\,
            I => \N__28718\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__28718\,
            I => \N__28711\
        );

    \I__6227\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28702\
        );

    \I__6226\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28702\
        );

    \I__6225\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28702\
        );

    \I__6224\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28702\
        );

    \I__6223\ : Odrv4
    port map (
            O => \N__28711\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__28702\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__6221\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28688\
        );

    \I__6220\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28688\
        );

    \I__6219\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28688\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__28688\,
            I => \POWERLED.count_clk_1_14\
        );

    \I__6217\ : CascadeMux
    port map (
            O => \N__28685\,
            I => \POWERLED.count_clkZ0Z_0_cascade_\
        );

    \I__6216\ : InMux
    port map (
            O => \N__28682\,
            I => \N__28676\
        );

    \I__6215\ : InMux
    port map (
            O => \N__28681\,
            I => \N__28676\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__28676\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28669\
        );

    \I__6212\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28666\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__28669\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__28666\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__6209\ : CascadeMux
    port map (
            O => \N__28661\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_1_cascade_\
        );

    \I__6208\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28655\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__28655\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_2\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__28652\,
            I => \N__28649\
        );

    \I__6205\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28645\
        );

    \I__6204\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28642\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__28645\,
            I => \POWERLED.count_clk_RNISLCE7Z0Z_10\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__28642\,
            I => \POWERLED.count_clk_RNISLCE7Z0Z_10\
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__28637\,
            I => \N__28634\
        );

    \I__6200\ : InMux
    port map (
            O => \N__28634\,
            I => \N__28631\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__28631\,
            I => \POWERLED.count_clk_en_917_0\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__28628\,
            I => \N__28625\
        );

    \I__6197\ : InMux
    port map (
            O => \N__28625\,
            I => \N__28618\
        );

    \I__6196\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28618\
        );

    \I__6195\ : InMux
    port map (
            O => \N__28623\,
            I => \N__28615\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__28618\,
            I => \N__28612\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__28615\,
            I => \N__28609\
        );

    \I__6192\ : Span4Mux_v
    port map (
            O => \N__28612\,
            I => \N__28604\
        );

    \I__6191\ : Span4Mux_s3_h
    port map (
            O => \N__28609\,
            I => \N__28604\
        );

    \I__6190\ : Odrv4
    port map (
            O => \N__28604\,
            I => \POWERLED.func_state_RNIBVNS_2Z0Z_0\
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__28601\,
            I => \POWERLED.count_clk_en_1_cascade_\
        );

    \I__6188\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28594\
        );

    \I__6187\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28591\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__28594\,
            I => \N__28585\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__28591\,
            I => \N__28585\
        );

    \I__6184\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28582\
        );

    \I__6183\ : Span4Mux_s3_h
    port map (
            O => \N__28585\,
            I => \N__28579\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__28582\,
            I => \POWERLED.N_617\
        );

    \I__6181\ : Odrv4
    port map (
            O => \N__28579\,
            I => \POWERLED.N_617\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__28574\,
            I => \POWERLED.count_clk_en_cascade_\
        );

    \I__6179\ : CascadeMux
    port map (
            O => \N__28571\,
            I => \N__28568\
        );

    \I__6178\ : InMux
    port map (
            O => \N__28568\,
            I => \N__28565\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__28565\,
            I => \N__28562\
        );

    \I__6176\ : Odrv4
    port map (
            O => \N__28562\,
            I => \POWERLED.un1_count_clk_2_axb_12\
        );

    \I__6175\ : InMux
    port map (
            O => \N__28559\,
            I => \POWERLED.un1_count_clk_2_cry_12\
        );

    \I__6174\ : InMux
    port map (
            O => \N__28556\,
            I => \POWERLED.un1_count_clk_2_cry_13_cZ0\
        );

    \I__6173\ : InMux
    port map (
            O => \N__28553\,
            I => \N__28533\
        );

    \I__6172\ : InMux
    port map (
            O => \N__28552\,
            I => \N__28533\
        );

    \I__6171\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28533\
        );

    \I__6170\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28524\
        );

    \I__6169\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28524\
        );

    \I__6168\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28524\
        );

    \I__6167\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28524\
        );

    \I__6166\ : CascadeMux
    port map (
            O => \N__28546\,
            I => \N__28517\
        );

    \I__6165\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28509\
        );

    \I__6164\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28509\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28543\,
            I => \N__28509\
        );

    \I__6162\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28502\
        );

    \I__6161\ : InMux
    port map (
            O => \N__28541\,
            I => \N__28502\
        );

    \I__6160\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28502\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__28533\,
            I => \N__28497\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28497\
        );

    \I__6157\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28484\
        );

    \I__6156\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28484\
        );

    \I__6155\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28484\
        );

    \I__6154\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28484\
        );

    \I__6153\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28484\
        );

    \I__6152\ : InMux
    port map (
            O => \N__28516\,
            I => \N__28484\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__28509\,
            I => \POWERLED.func_state_RNI2VV9A_0_0\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__28502\,
            I => \POWERLED.func_state_RNI2VV9A_0_0\
        );

    \I__6149\ : Odrv4
    port map (
            O => \N__28497\,
            I => \POWERLED.func_state_RNI2VV9A_0_0\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__28484\,
            I => \POWERLED.func_state_RNI2VV9A_0_0\
        );

    \I__6147\ : InMux
    port map (
            O => \N__28475\,
            I => \POWERLED.un1_count_clk_2_cry_14\
        );

    \I__6146\ : InMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__6144\ : Odrv12
    port map (
            O => \N__28466\,
            I => \POWERLED.count_clk_0_15\
        );

    \I__6143\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28460\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__28460\,
            I => \N__28456\
        );

    \I__6141\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28453\
        );

    \I__6140\ : Odrv12
    port map (
            O => \N__28456\,
            I => \POWERLED.count_clk_1_15\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__28453\,
            I => \POWERLED.count_clk_1_15\
        );

    \I__6138\ : InMux
    port map (
            O => \N__28448\,
            I => \N__28444\
        );

    \I__6137\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28441\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__28444\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__28441\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__6134\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__6132\ : Span4Mux_v
    port map (
            O => \N__28430\,
            I => \N__28425\
        );

    \I__6131\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28420\
        );

    \I__6130\ : InMux
    port map (
            O => \N__28428\,
            I => \N__28420\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__28425\,
            I => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__28420\,
            I => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\
        );

    \I__6127\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28409\
        );

    \I__6126\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28409\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__28409\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__6124\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28403\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__28403\,
            I => \POWERLED.un1_count_clk_2_axb_10\
        );

    \I__6122\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28397\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__28397\,
            I => \POWERLED.un1_count_clk_2_axb_14\
        );

    \I__6120\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28388\
        );

    \I__6119\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28388\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__28388\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__6117\ : InMux
    port map (
            O => \N__28385\,
            I => \POWERLED.un1_count_clk_2_cry_3\
        );

    \I__6116\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28378\
        );

    \I__6115\ : CascadeMux
    port map (
            O => \N__28381\,
            I => \N__28374\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__28378\,
            I => \N__28371\
        );

    \I__6113\ : InMux
    port map (
            O => \N__28377\,
            I => \N__28368\
        );

    \I__6112\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28365\
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__28371\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__28368\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__28365\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__6108\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28352\
        );

    \I__6107\ : InMux
    port map (
            O => \N__28357\,
            I => \N__28352\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__28352\,
            I => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\
        );

    \I__6105\ : InMux
    port map (
            O => \N__28349\,
            I => \POWERLED.un1_count_clk_2_cry_4\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28346\,
            I => \N__28339\
        );

    \I__6103\ : InMux
    port map (
            O => \N__28345\,
            I => \N__28339\
        );

    \I__6102\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28336\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__28339\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__28336\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__6099\ : InMux
    port map (
            O => \N__28331\,
            I => \N__28325\
        );

    \I__6098\ : InMux
    port map (
            O => \N__28330\,
            I => \N__28325\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__28325\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__6096\ : InMux
    port map (
            O => \N__28322\,
            I => \POWERLED.un1_count_clk_2_cry_5\
        );

    \I__6095\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28315\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__28318\,
            I => \N__28311\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__28315\,
            I => \N__28307\
        );

    \I__6092\ : InMux
    port map (
            O => \N__28314\,
            I => \N__28304\
        );

    \I__6091\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28301\
        );

    \I__6090\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28297\
        );

    \I__6089\ : Span4Mux_s2_h
    port map (
            O => \N__28307\,
            I => \N__28294\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__28304\,
            I => \N__28291\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__28301\,
            I => \N__28288\
        );

    \I__6086\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28285\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28282\
        );

    \I__6084\ : Span4Mux_h
    port map (
            O => \N__28294\,
            I => \N__28277\
        );

    \I__6083\ : Span4Mux_s2_h
    port map (
            O => \N__28291\,
            I => \N__28277\
        );

    \I__6082\ : Span4Mux_s2_h
    port map (
            O => \N__28288\,
            I => \N__28274\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__28285\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__6080\ : Odrv12
    port map (
            O => \N__28282\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__28277\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__28274\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__6077\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28259\
        );

    \I__6076\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28259\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__28259\,
            I => \N__28256\
        );

    \I__6074\ : Span4Mux_h
    port map (
            O => \N__28256\,
            I => \N__28253\
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__28253\,
            I => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\
        );

    \I__6072\ : InMux
    port map (
            O => \N__28250\,
            I => \POWERLED.un1_count_clk_2_cry_6\
        );

    \I__6071\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28242\
        );

    \I__6070\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28237\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28237\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__28242\,
            I => \N__28234\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__28237\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__6066\ : Odrv4
    port map (
            O => \N__28234\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__6065\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28223\
        );

    \I__6064\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28223\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__28223\,
            I => \N__28220\
        );

    \I__6062\ : Odrv4
    port map (
            O => \N__28220\,
            I => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\
        );

    \I__6061\ : InMux
    port map (
            O => \N__28217\,
            I => \POWERLED.un1_count_clk_2_cry_7\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28210\
        );

    \I__6059\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28206\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28203\
        );

    \I__6057\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28200\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__28206\,
            I => \N__28193\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__28203\,
            I => \N__28193\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__28200\,
            I => \N__28193\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__28193\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__6052\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28186\
        );

    \I__6051\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28183\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__28186\,
            I => \N__28178\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__28183\,
            I => \N__28178\
        );

    \I__6048\ : Odrv4
    port map (
            O => \N__28178\,
            I => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\
        );

    \I__6047\ : InMux
    port map (
            O => \N__28175\,
            I => \bfn_12_6_0_\
        );

    \I__6046\ : InMux
    port map (
            O => \N__28172\,
            I => \POWERLED.un1_count_clk_2_cry_9\
        );

    \I__6045\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28163\
        );

    \I__6044\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28163\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__28163\,
            I => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\
        );

    \I__6042\ : InMux
    port map (
            O => \N__28160\,
            I => \POWERLED.un1_count_clk_2_cry_10\
        );

    \I__6041\ : InMux
    port map (
            O => \N__28157\,
            I => \POWERLED.un1_count_clk_2_cry_11_cZ0\
        );

    \I__6040\ : CascadeMux
    port map (
            O => \N__28154\,
            I => \POWERLED.count_clkZ0Z_3_cascade_\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__28151\,
            I => \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_\
        );

    \I__6038\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28142\
        );

    \I__6037\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28142\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__28142\,
            I => \N__28139\
        );

    \I__6035\ : Odrv4
    port map (
            O => \N__28139\,
            I => \POWERLED.count_clk_0_3\
        );

    \I__6034\ : CascadeMux
    port map (
            O => \N__28136\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_\
        );

    \I__6033\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28129\
        );

    \I__6032\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__28129\,
            I => \N__28123\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__28126\,
            I => \N__28120\
        );

    \I__6029\ : Span4Mux_h
    port map (
            O => \N__28123\,
            I => \N__28117\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__28120\,
            I => \POWERLED.N_625\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__28117\,
            I => \POWERLED.N_625\
        );

    \I__6026\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28107\
        );

    \I__6025\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28102\
        );

    \I__6024\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28102\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__28107\,
            I => \N__28099\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28096\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__28099\,
            I => \POWERLED.count_clk_RNIZ0Z_1\
        );

    \I__6020\ : Odrv4
    port map (
            O => \N__28096\,
            I => \POWERLED.count_clk_RNIZ0Z_1\
        );

    \I__6019\ : CascadeMux
    port map (
            O => \N__28091\,
            I => \POWERLED.N_625_cascade_\
        );

    \I__6018\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28085\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__28085\,
            I => \N__28082\
        );

    \I__6016\ : Span4Mux_v
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__28079\,
            I => \POWERLED.count_clk_RNIPGQN2_5Z0Z_3\
        );

    \I__6014\ : CascadeMux
    port map (
            O => \N__28076\,
            I => \N__28072\
        );

    \I__6013\ : CascadeMux
    port map (
            O => \N__28075\,
            I => \N__28067\
        );

    \I__6012\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28064\
        );

    \I__6011\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28059\
        );

    \I__6010\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28059\
        );

    \I__6009\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28056\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__28064\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__28059\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__28056\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6005\ : CascadeMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__6004\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28041\
        );

    \I__6003\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28036\
        );

    \I__6002\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28036\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__28041\,
            I => \N__28033\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__28036\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__5999\ : Odrv4
    port map (
            O => \N__28033\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__5998\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28022\
        );

    \I__5997\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28022\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__28022\,
            I => \N__28019\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__28019\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__5994\ : InMux
    port map (
            O => \N__28016\,
            I => \POWERLED.un1_count_clk_2_cry_1\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__5992\ : InMux
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__28007\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__5990\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27995\
        );

    \I__5989\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27995\
        );

    \I__5988\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27995\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__27995\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__5986\ : InMux
    port map (
            O => \N__27992\,
            I => \POWERLED.un1_count_clk_2_cry_2\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__27989\,
            I => \N__27984\
        );

    \I__5984\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27981\
        );

    \I__5983\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27978\
        );

    \I__5982\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27975\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__27981\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__27978\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__27975\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__5978\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__27965\,
            I => \POWERLED.N_529\
        );

    \I__5976\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27956\
        );

    \I__5975\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27956\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__27953\,
            I => \POWERLED.dutycycle_en_12\
        );

    \I__5972\ : InMux
    port map (
            O => \N__27950\,
            I => \N__27947\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__27947\,
            I => \POWERLED.count_clk_0_8\
        );

    \I__5970\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27941\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__27941\,
            I => \POWERLED.count_clk_0_9\
        );

    \I__5968\ : InMux
    port map (
            O => \N__27938\,
            I => \N__27935\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__27935\,
            I => \POWERLED.count_clk_0_2\
        );

    \I__5966\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27929\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27926\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__27926\,
            I => \N__27923\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__27923\,
            I => \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_d\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__27920\,
            I => \POWERLED.N_526_cascade_\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__27917\,
            I => \N__27914\
        );

    \I__5960\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27908\
        );

    \I__5959\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27908\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__27908\,
            I => \N__27905\
        );

    \I__5957\ : Odrv12
    port map (
            O => \N__27905\,
            I => \POWERLED.dutycycle_RNI36306Z0Z_14\
        );

    \I__5956\ : CascadeMux
    port map (
            O => \N__27902\,
            I => \N__27898\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__27901\,
            I => \N__27894\
        );

    \I__5954\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27886\
        );

    \I__5953\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27886\
        );

    \I__5952\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27881\
        );

    \I__5951\ : InMux
    port map (
            O => \N__27893\,
            I => \N__27881\
        );

    \I__5950\ : CascadeMux
    port map (
            O => \N__27892\,
            I => \N__27875\
        );

    \I__5949\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27872\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27867\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__27881\,
            I => \N__27867\
        );

    \I__5946\ : InMux
    port map (
            O => \N__27880\,
            I => \N__27862\
        );

    \I__5945\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27862\
        );

    \I__5944\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27856\
        );

    \I__5943\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27856\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__27872\,
            I => \N__27849\
        );

    \I__5941\ : Span4Mux_s3_v
    port map (
            O => \N__27867\,
            I => \N__27849\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__27862\,
            I => \N__27849\
        );

    \I__5939\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27846\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__27856\,
            I => \N__27841\
        );

    \I__5937\ : Span4Mux_v
    port map (
            O => \N__27849\,
            I => \N__27841\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__27846\,
            I => \POWERLED.func_state_RNI_8Z0Z_1\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__27841\,
            I => \POWERLED.func_state_RNI_8Z0Z_1\
        );

    \I__5934\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27826\
        );

    \I__5933\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27826\
        );

    \I__5932\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27820\
        );

    \I__5931\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27820\
        );

    \I__5930\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27814\
        );

    \I__5929\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27814\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__27826\,
            I => \N__27811\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__27825\,
            I => \N__27807\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__27820\,
            I => \N__27804\
        );

    \I__5925\ : InMux
    port map (
            O => \N__27819\,
            I => \N__27801\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__27814\,
            I => \N__27798\
        );

    \I__5923\ : Span4Mux_s2_v
    port map (
            O => \N__27811\,
            I => \N__27795\
        );

    \I__5922\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27792\
        );

    \I__5921\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27789\
        );

    \I__5920\ : Span4Mux_h
    port map (
            O => \N__27804\,
            I => \N__27786\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__27801\,
            I => \N__27779\
        );

    \I__5918\ : Span4Mux_s2_v
    port map (
            O => \N__27798\,
            I => \N__27779\
        );

    \I__5917\ : Span4Mux_h
    port map (
            O => \N__27795\,
            I => \N__27779\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__27792\,
            I => \POWERLED.N_203\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__27789\,
            I => \POWERLED.N_203\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__27786\,
            I => \POWERLED.N_203\
        );

    \I__5913\ : Odrv4
    port map (
            O => \N__27779\,
            I => \POWERLED.N_203\
        );

    \I__5912\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27764\
        );

    \I__5911\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27756\
        );

    \I__5910\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27756\
        );

    \I__5909\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27756\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__27764\,
            I => \N__27751\
        );

    \I__5907\ : CascadeMux
    port map (
            O => \N__27763\,
            I => \N__27748\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__27756\,
            I => \N__27740\
        );

    \I__5905\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27737\
        );

    \I__5904\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27734\
        );

    \I__5903\ : Span4Mux_s3_h
    port map (
            O => \N__27751\,
            I => \N__27731\
        );

    \I__5902\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27726\
        );

    \I__5901\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27726\
        );

    \I__5900\ : InMux
    port map (
            O => \N__27746\,
            I => \N__27721\
        );

    \I__5899\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27721\
        );

    \I__5898\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27716\
        );

    \I__5897\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27716\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__27740\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__27737\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__27734\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__27731\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__27726\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__27721\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__27716\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__27701\,
            I => \POWERLED.N_524_cascade_\
        );

    \I__5888\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27695\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__27695\,
            I => \POWERLED.un1_clk_100khz_47_and_i_1\
        );

    \I__5886\ : IoInMux
    port map (
            O => \N__27692\,
            I => \N__27689\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__27689\,
            I => \N__27684\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__27688\,
            I => \N__27681\
        );

    \I__5883\ : CascadeMux
    port map (
            O => \N__27687\,
            I => \N__27678\
        );

    \I__5882\ : IoSpan4Mux
    port map (
            O => \N__27684\,
            I => \N__27674\
        );

    \I__5881\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27667\
        );

    \I__5880\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27667\
        );

    \I__5879\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27660\
        );

    \I__5878\ : Span4Mux_s2_v
    port map (
            O => \N__27674\,
            I => \N__27657\
        );

    \I__5877\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27654\
        );

    \I__5876\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27651\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__27667\,
            I => \N__27648\
        );

    \I__5874\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27645\
        );

    \I__5873\ : CascadeMux
    port map (
            O => \N__27665\,
            I => \N__27641\
        );

    \I__5872\ : CascadeMux
    port map (
            O => \N__27664\,
            I => \N__27637\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__27663\,
            I => \N__27634\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__27660\,
            I => \N__27631\
        );

    \I__5869\ : Span4Mux_h
    port map (
            O => \N__27657\,
            I => \N__27626\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__27654\,
            I => \N__27626\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__27651\,
            I => \N__27618\
        );

    \I__5866\ : Span4Mux_v
    port map (
            O => \N__27648\,
            I => \N__27612\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__27645\,
            I => \N__27612\
        );

    \I__5864\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27609\
        );

    \I__5863\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27600\
        );

    \I__5862\ : InMux
    port map (
            O => \N__27640\,
            I => \N__27600\
        );

    \I__5861\ : InMux
    port map (
            O => \N__27637\,
            I => \N__27600\
        );

    \I__5860\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27600\
        );

    \I__5859\ : Span4Mux_s2_v
    port map (
            O => \N__27631\,
            I => \N__27595\
        );

    \I__5858\ : Span4Mux_h
    port map (
            O => \N__27626\,
            I => \N__27595\
        );

    \I__5857\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27590\
        );

    \I__5856\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27590\
        );

    \I__5855\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27583\
        );

    \I__5854\ : InMux
    port map (
            O => \N__27622\,
            I => \N__27583\
        );

    \I__5853\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27583\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__27618\,
            I => \N__27579\
        );

    \I__5851\ : CascadeMux
    port map (
            O => \N__27617\,
            I => \N__27576\
        );

    \I__5850\ : Span4Mux_v
    port map (
            O => \N__27612\,
            I => \N__27569\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__27609\,
            I => \N__27569\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27566\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__27595\,
            I => \N__27559\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__27590\,
            I => \N__27559\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__27583\,
            I => \N__27559\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__27582\,
            I => \N__27556\
        );

    \I__5843\ : Span4Mux_v
    port map (
            O => \N__27579\,
            I => \N__27553\
        );

    \I__5842\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27546\
        );

    \I__5841\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27546\
        );

    \I__5840\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27546\
        );

    \I__5839\ : Span4Mux_h
    port map (
            O => \N__27569\,
            I => \N__27543\
        );

    \I__5838\ : Span4Mux_v
    port map (
            O => \N__27566\,
            I => \N__27538\
        );

    \I__5837\ : Span4Mux_v
    port map (
            O => \N__27559\,
            I => \N__27538\
        );

    \I__5836\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27535\
        );

    \I__5835\ : Odrv4
    port map (
            O => \N__27553\,
            I => rsmrstn
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__27546\,
            I => rsmrstn
        );

    \I__5833\ : Odrv4
    port map (
            O => \N__27543\,
            I => rsmrstn
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__27538\,
            I => rsmrstn
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__27535\,
            I => rsmrstn
        );

    \I__5830\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27521\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27516\
        );

    \I__5828\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27513\
        );

    \I__5827\ : CascadeMux
    port map (
            O => \N__27519\,
            I => \N__27507\
        );

    \I__5826\ : Span4Mux_v
    port map (
            O => \N__27516\,
            I => \N__27503\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__27513\,
            I => \N__27500\
        );

    \I__5824\ : InMux
    port map (
            O => \N__27512\,
            I => \N__27497\
        );

    \I__5823\ : InMux
    port map (
            O => \N__27511\,
            I => \N__27492\
        );

    \I__5822\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27492\
        );

    \I__5821\ : InMux
    port map (
            O => \N__27507\,
            I => \N__27487\
        );

    \I__5820\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27487\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__27503\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__5818\ : Odrv12
    port map (
            O => \N__27500\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__27497\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__27492\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__27487\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__27476\,
            I => \N__27472\
        );

    \I__5813\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27467\
        );

    \I__5812\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27467\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__27467\,
            I => \N__27464\
        );

    \I__5810\ : Odrv12
    port map (
            O => \N__27464\,
            I => \POWERLED.N_2381_i\
        );

    \I__5809\ : CascadeMux
    port map (
            O => \N__27461\,
            I => \N__27453\
        );

    \I__5808\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27446\
        );

    \I__5807\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27446\
        );

    \I__5806\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27443\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__27457\,
            I => \N__27439\
        );

    \I__5804\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27436\
        );

    \I__5803\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27431\
        );

    \I__5802\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27431\
        );

    \I__5801\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27428\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27425\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__27443\,
            I => \N__27422\
        );

    \I__5798\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27419\
        );

    \I__5797\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27416\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27413\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__27431\,
            I => \N__27410\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__27428\,
            I => \N__27401\
        );

    \I__5793\ : Span4Mux_v
    port map (
            O => \N__27425\,
            I => \N__27401\
        );

    \I__5792\ : Span4Mux_v
    port map (
            O => \N__27422\,
            I => \N__27401\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__27419\,
            I => \N__27401\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__27416\,
            I => \N__27396\
        );

    \I__5789\ : Span4Mux_s2_h
    port map (
            O => \N__27413\,
            I => \N__27396\
        );

    \I__5788\ : Span4Mux_v
    port map (
            O => \N__27410\,
            I => \N__27391\
        );

    \I__5787\ : Span4Mux_v
    port map (
            O => \N__27401\,
            I => \N__27391\
        );

    \I__5786\ : Span4Mux_v
    port map (
            O => \N__27396\,
            I => \N__27388\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__27391\,
            I => \POWERLED.N_91_1_N\
        );

    \I__5784\ : Odrv4
    port map (
            O => \N__27388\,
            I => \POWERLED.N_91_1_N\
        );

    \I__5783\ : CascadeMux
    port map (
            O => \N__27383\,
            I => \POWERLED.N_527_cascade_\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__27380\,
            I => \POWERLED.un1_clk_100khz_48_and_i_1_cascade_\
        );

    \I__5781\ : CascadeMux
    port map (
            O => \N__27377\,
            I => \N__27365\
        );

    \I__5780\ : CascadeMux
    port map (
            O => \N__27376\,
            I => \N__27361\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__27375\,
            I => \N__27356\
        );

    \I__5778\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27347\
        );

    \I__5777\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27347\
        );

    \I__5776\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27347\
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__27371\,
            I => \N__27337\
        );

    \I__5774\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27328\
        );

    \I__5773\ : InMux
    port map (
            O => \N__27369\,
            I => \N__27328\
        );

    \I__5772\ : InMux
    port map (
            O => \N__27368\,
            I => \N__27328\
        );

    \I__5771\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27328\
        );

    \I__5770\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27325\
        );

    \I__5769\ : InMux
    port map (
            O => \N__27361\,
            I => \N__27316\
        );

    \I__5768\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27316\
        );

    \I__5767\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27316\
        );

    \I__5766\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27316\
        );

    \I__5765\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27313\
        );

    \I__5764\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27310\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__27347\,
            I => \N__27307\
        );

    \I__5762\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27302\
        );

    \I__5761\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27302\
        );

    \I__5760\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27299\
        );

    \I__5759\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27290\
        );

    \I__5758\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27290\
        );

    \I__5757\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27290\
        );

    \I__5756\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27290\
        );

    \I__5755\ : InMux
    port map (
            O => \N__27337\,
            I => \N__27287\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__27328\,
            I => \N__27280\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27280\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__27316\,
            I => \N__27280\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__27313\,
            I => \N__27275\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__27310\,
            I => \N__27275\
        );

    \I__5749\ : Odrv12
    port map (
            O => \N__27307\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__27302\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__27299\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__27290\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__27287\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__27280\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__27275\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__27260\,
            I => \POWERLED.un1_clk_100khz_30_and_i_0_a2_5_0_0_cascade_\
        );

    \I__5741\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27254\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__27254\,
            I => \POWERLED.dutycycle_eena_2_0_0_tz_1\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__27251\,
            I => \POWERLED.dutycycle_eena_2_d_0_cascade_\
        );

    \I__5738\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27242\
        );

    \I__5737\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27242\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27239\
        );

    \I__5735\ : Odrv12
    port map (
            O => \N__27239\,
            I => \POWERLED.dutycycle_RNIRUFD6Z0Z_9\
        );

    \I__5734\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27229\
        );

    \I__5733\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__5732\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27224\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27221\
        );

    \I__5730\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27216\
        );

    \I__5729\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27216\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__27224\,
            I => \N__27213\
        );

    \I__5727\ : Span4Mux_s3_v
    port map (
            O => \N__27221\,
            I => \N__27210\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__27216\,
            I => \N__27207\
        );

    \I__5725\ : Span4Mux_h
    port map (
            O => \N__27213\,
            I => \N__27202\
        );

    \I__5724\ : Span4Mux_h
    port map (
            O => \N__27210\,
            I => \N__27197\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__27207\,
            I => \N__27197\
        );

    \I__5722\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27192\
        );

    \I__5721\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27192\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__27202\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__27197\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__27192\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__27185\,
            I => \N__27181\
        );

    \I__5716\ : InMux
    port map (
            O => \N__27184\,
            I => \N__27178\
        );

    \I__5715\ : InMux
    port map (
            O => \N__27181\,
            I => \N__27168\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__27178\,
            I => \N__27165\
        );

    \I__5713\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27160\
        );

    \I__5712\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27160\
        );

    \I__5711\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27157\
        );

    \I__5710\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27152\
        );

    \I__5709\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27152\
        );

    \I__5708\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27146\
        );

    \I__5707\ : InMux
    port map (
            O => \N__27171\,
            I => \N__27146\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__27168\,
            I => \N__27141\
        );

    \I__5705\ : Span4Mux_v
    port map (
            O => \N__27165\,
            I => \N__27141\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__27138\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__27157\,
            I => \N__27133\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__27152\,
            I => \N__27133\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__27151\,
            I => \N__27130\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__27146\,
            I => \N__27127\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__27141\,
            I => \N__27122\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__27138\,
            I => \N__27122\
        );

    \I__5697\ : Span4Mux_h
    port map (
            O => \N__27133\,
            I => \N__27119\
        );

    \I__5696\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27116\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__27127\,
            I => \RSMRSTn_rep1\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__27122\,
            I => \RSMRSTn_rep1\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__27119\,
            I => \RSMRSTn_rep1\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__27116\,
            I => \RSMRSTn_rep1\
        );

    \I__5691\ : CascadeMux
    port map (
            O => \N__27107\,
            I => \N__27100\
        );

    \I__5690\ : CascadeMux
    port map (
            O => \N__27106\,
            I => \N__27093\
        );

    \I__5689\ : CascadeMux
    port map (
            O => \N__27105\,
            I => \N__27090\
        );

    \I__5688\ : CascadeMux
    port map (
            O => \N__27104\,
            I => \N__27086\
        );

    \I__5687\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27082\
        );

    \I__5686\ : InMux
    port map (
            O => \N__27100\,
            I => \N__27079\
        );

    \I__5685\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27076\
        );

    \I__5684\ : CascadeMux
    port map (
            O => \N__27098\,
            I => \N__27070\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__27097\,
            I => \N__27067\
        );

    \I__5682\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27058\
        );

    \I__5681\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27058\
        );

    \I__5680\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27058\
        );

    \I__5679\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27051\
        );

    \I__5678\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27051\
        );

    \I__5677\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27051\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__27082\,
            I => \N__27046\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__27079\,
            I => \N__27046\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__27076\,
            I => \N__27043\
        );

    \I__5673\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27040\
        );

    \I__5672\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27033\
        );

    \I__5671\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27033\
        );

    \I__5670\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27033\
        );

    \I__5669\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27028\
        );

    \I__5668\ : InMux
    port map (
            O => \N__27066\,
            I => \N__27028\
        );

    \I__5667\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27025\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__27058\,
            I => \N__27020\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__27051\,
            I => \N__27020\
        );

    \I__5664\ : Span4Mux_v
    port map (
            O => \N__27046\,
            I => \N__27015\
        );

    \I__5663\ : Span4Mux_v
    port map (
            O => \N__27043\,
            I => \N__27015\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27040\,
            I => \N__27004\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__27033\,
            I => \N__27004\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__27028\,
            I => \N__27004\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__27025\,
            I => \N__27004\
        );

    \I__5658\ : Span4Mux_s3_v
    port map (
            O => \N__27020\,
            I => \N__27004\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__27015\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__27004\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__26999\,
            I => \POWERLED.N_520_cascade_\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__26996\,
            I => \N__26993\
        );

    \I__5653\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26989\
        );

    \I__5652\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26986\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__26989\,
            I => \N__26981\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__26986\,
            I => \N__26981\
        );

    \I__5649\ : Odrv4
    port map (
            O => \N__26981\,
            I => \POWERLED.dutycycle_RNIRUFD6Z0Z_12\
        );

    \I__5648\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26970\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__26977\,
            I => \N__26964\
        );

    \I__5646\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26956\
        );

    \I__5645\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26956\
        );

    \I__5644\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26956\
        );

    \I__5643\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26953\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__26970\,
            I => \N__26949\
        );

    \I__5641\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26942\
        );

    \I__5640\ : InMux
    port map (
            O => \N__26968\,
            I => \N__26942\
        );

    \I__5639\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26942\
        );

    \I__5638\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26939\
        );

    \I__5637\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26936\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__26956\,
            I => \N__26931\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__26953\,
            I => \N__26931\
        );

    \I__5634\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26928\
        );

    \I__5633\ : Span4Mux_h
    port map (
            O => \N__26949\,
            I => \N__26923\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__26942\,
            I => \N__26923\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__26939\,
            I => \N__26920\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__26936\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5629\ : Odrv12
    port map (
            O => \N__26931\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__26928\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__26923\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__26920\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5625\ : CascadeMux
    port map (
            O => \N__26909\,
            I => \POWERLED.N_518_cascade_\
        );

    \I__5624\ : InMux
    port map (
            O => \N__26906\,
            I => \N__26903\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__26903\,
            I => \POWERLED.un1_clk_100khz_42_and_i_1\
        );

    \I__5622\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26897\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__26897\,
            I => \N__26894\
        );

    \I__5620\ : Span4Mux_h
    port map (
            O => \N__26894\,
            I => \N__26891\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__26891\,
            I => \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_0_3_1\
        );

    \I__5618\ : CascadeMux
    port map (
            O => \N__26888\,
            I => \POWERLED.N_203_cascade_\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__26885\,
            I => \POWERLED.N_521_cascade_\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__26882\,
            I => \POWERLED.un1_clk_100khz_43_and_i_1_cascade_\
        );

    \I__5615\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__26876\,
            I => \POWERLED.N_523\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__26873\,
            I => \POWERLED.N_503_cascade_\
        );

    \I__5612\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26864\
        );

    \I__5611\ : InMux
    port map (
            O => \N__26869\,
            I => \N__26864\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__26864\,
            I => \N__26861\
        );

    \I__5609\ : Odrv12
    port map (
            O => \N__26861\,
            I => \POWERLED.dutycycle_1_0_0\
        );

    \I__5608\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26855\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__26855\,
            I => \POWERLED.dutycycle_eena\
        );

    \I__5606\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26846\
        );

    \I__5605\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26846\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__26846\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__5603\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26840\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26837\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__26837\,
            I => \N__26834\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__26834\,
            I => \POWERLED.N_510\
        );

    \I__5599\ : CascadeMux
    port map (
            O => \N__26831\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_a2_c_cascade_\
        );

    \I__5598\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26825\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26817\
        );

    \I__5596\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26806\
        );

    \I__5595\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26806\
        );

    \I__5594\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26806\
        );

    \I__5593\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26806\
        );

    \I__5592\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26806\
        );

    \I__5591\ : Span12Mux_s10_v
    port map (
            O => \N__26817\,
            I => \N__26799\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__26806\,
            I => \N__26799\
        );

    \I__5589\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26796\
        );

    \I__5588\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26793\
        );

    \I__5587\ : Odrv12
    port map (
            O => \N__26799\,
            I => rsmrst_pwrgd_signal
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__26796\,
            I => rsmrst_pwrgd_signal
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__26793\,
            I => rsmrst_pwrgd_signal
        );

    \I__5584\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__26783\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_a2_d\
        );

    \I__5582\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__26777\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_0_2\
        );

    \I__5580\ : CascadeMux
    port map (
            O => \N__26774\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d_cascade_\
        );

    \I__5579\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26765\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26765\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__5576\ : Span4Mux_h
    port map (
            O => \N__26762\,
            I => \N__26759\
        );

    \I__5575\ : Odrv4
    port map (
            O => \N__26759\,
            I => \POWERLED.dutycycle_eena_5\
        );

    \I__5574\ : CascadeMux
    port map (
            O => \N__26756\,
            I => \N__26749\
        );

    \I__5573\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26739\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__26754\,
            I => \N__26736\
        );

    \I__5571\ : InMux
    port map (
            O => \N__26753\,
            I => \N__26731\
        );

    \I__5570\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26728\
        );

    \I__5569\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26721\
        );

    \I__5568\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26721\
        );

    \I__5567\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26721\
        );

    \I__5566\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26718\
        );

    \I__5565\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26715\
        );

    \I__5564\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26710\
        );

    \I__5563\ : InMux
    port map (
            O => \N__26743\,
            I => \N__26710\
        );

    \I__5562\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26704\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__26739\,
            I => \N__26701\
        );

    \I__5560\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26694\
        );

    \I__5559\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26694\
        );

    \I__5558\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26694\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26691\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__26728\,
            I => \N__26682\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__26721\,
            I => \N__26682\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26682\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__26715\,
            I => \N__26682\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__26710\,
            I => \N__26679\
        );

    \I__5551\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26676\
        );

    \I__5550\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26671\
        );

    \I__5549\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26671\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__26704\,
            I => \N__26668\
        );

    \I__5547\ : Span4Mux_v
    port map (
            O => \N__26701\,
            I => \N__26663\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26663\
        );

    \I__5545\ : Span4Mux_v
    port map (
            O => \N__26691\,
            I => \N__26658\
        );

    \I__5544\ : Span4Mux_v
    port map (
            O => \N__26682\,
            I => \N__26658\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__26679\,
            I => \N__26651\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__26676\,
            I => \N__26651\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__26671\,
            I => \N__26651\
        );

    \I__5540\ : Span12Mux_v
    port map (
            O => \N__26668\,
            I => \N__26648\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__26663\,
            I => \N__26645\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__26658\,
            I => \N__26640\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__26651\,
            I => \N__26640\
        );

    \I__5536\ : Odrv12
    port map (
            O => \N__26648\,
            I => gpio_fpga_soc_4
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__26645\,
            I => gpio_fpga_soc_4
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__26640\,
            I => gpio_fpga_soc_4
        );

    \I__5533\ : CascadeMux
    port map (
            O => \N__26633\,
            I => \POWERLED.N_249_cascade_\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__26630\,
            I => \POWERLED.N_546_cascade_\
        );

    \I__5531\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26620\
        );

    \I__5529\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26617\
        );

    \I__5528\ : Span4Mux_h
    port map (
            O => \N__26620\,
            I => \N__26614\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__5526\ : Odrv4
    port map (
            O => \N__26614\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_0\
        );

    \I__5525\ : Odrv12
    port map (
            O => \N__26611\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_0\
        );

    \I__5524\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__26603\,
            I => \POWERLED.N_482\
        );

    \I__5522\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26597\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__26597\,
            I => \N__26594\
        );

    \I__5520\ : Odrv12
    port map (
            O => \N__26594\,
            I => \POWERLED.g0_i_m2_rn_1_0\
        );

    \I__5519\ : CascadeMux
    port map (
            O => \N__26591\,
            I => \POWERLED.dutycycleZ0Z_1_cascade_\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__26588\,
            I => \N__26585\
        );

    \I__5517\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__26582\,
            I => \POWERLED.dutycycle_eena_0_0\
        );

    \I__5515\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26575\
        );

    \I__5514\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26572\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__26575\,
            I => \N__26569\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__26572\,
            I => \POWERLED.g0_1\
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__26569\,
            I => \POWERLED.g0_1\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__26564\,
            I => \POWERLED.dutycycle_eena_0_0_cascade_\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__26561\,
            I => \POWERLED.dutycycle_eena_cascade_\
        );

    \I__5508\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26554\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__26557\,
            I => \N__26549\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__26554\,
            I => \N__26544\
        );

    \I__5505\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26541\
        );

    \I__5504\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26537\
        );

    \I__5503\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26532\
        );

    \I__5502\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26532\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__26547\,
            I => \N__26529\
        );

    \I__5500\ : Span4Mux_h
    port map (
            O => \N__26544\,
            I => \N__26526\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__26541\,
            I => \N__26523\
        );

    \I__5498\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26519\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26516\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__26532\,
            I => \N__26513\
        );

    \I__5495\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26510\
        );

    \I__5494\ : Span4Mux_h
    port map (
            O => \N__26526\,
            I => \N__26505\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__26523\,
            I => \N__26502\
        );

    \I__5492\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26499\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__26519\,
            I => \N__26496\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__26516\,
            I => \N__26489\
        );

    \I__5489\ : Span4Mux_v
    port map (
            O => \N__26513\,
            I => \N__26489\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__26510\,
            I => \N__26489\
        );

    \I__5487\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26484\
        );

    \I__5486\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26484\
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__26505\,
            I => \POWERLED.dutycycle\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__26502\,
            I => \POWERLED.dutycycle\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__26499\,
            I => \POWERLED.dutycycle\
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__26496\,
            I => \POWERLED.dutycycle\
        );

    \I__5481\ : Odrv4
    port map (
            O => \N__26489\,
            I => \POWERLED.dutycycle\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__26484\,
            I => \POWERLED.dutycycle\
        );

    \I__5479\ : CascadeMux
    port map (
            O => \N__26471\,
            I => \N__26467\
        );

    \I__5478\ : InMux
    port map (
            O => \N__26470\,
            I => \N__26462\
        );

    \I__5477\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26462\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__26462\,
            I => \POWERLED.g0_i_m2_sn\
        );

    \I__5475\ : CascadeMux
    port map (
            O => \N__26459\,
            I => \N__26450\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__26458\,
            I => \N__26447\
        );

    \I__5473\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26441\
        );

    \I__5472\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26441\
        );

    \I__5471\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26436\
        );

    \I__5470\ : InMux
    port map (
            O => \N__26454\,
            I => \N__26436\
        );

    \I__5469\ : InMux
    port map (
            O => \N__26453\,
            I => \N__26431\
        );

    \I__5468\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26431\
        );

    \I__5467\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26426\
        );

    \I__5466\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26426\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__26441\,
            I => \N__26416\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__26436\,
            I => \N__26416\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__26431\,
            I => \N__26416\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__26426\,
            I => \N__26416\
        );

    \I__5461\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26413\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__26416\,
            I => \N__26410\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__26413\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5458\ : Odrv4
    port map (
            O => \N__26410\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5457\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26399\
        );

    \I__5456\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26399\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__26399\,
            I => \POWERLED.g0_i_m2_rn_1\
        );

    \I__5454\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__26393\,
            I => \POWERLED.dutycycleZ1Z_1\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__5451\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26380\
        );

    \I__5450\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26377\
        );

    \I__5449\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26372\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26372\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__26383\,
            I => \N__26368\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__26380\,
            I => \N__26358\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__26377\,
            I => \N__26358\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26358\
        );

    \I__5443\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26353\
        );

    \I__5442\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26353\
        );

    \I__5441\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26350\
        );

    \I__5440\ : InMux
    port map (
            O => \N__26366\,
            I => \N__26346\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__26365\,
            I => \N__26343\
        );

    \I__5438\ : Span4Mux_v
    port map (
            O => \N__26358\,
            I => \N__26339\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__26353\,
            I => \N__26334\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__26350\,
            I => \N__26334\
        );

    \I__5435\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26331\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26328\
        );

    \I__5433\ : InMux
    port map (
            O => \N__26343\,
            I => \N__26325\
        );

    \I__5432\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26322\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__26339\,
            I => \N_247\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__26334\,
            I => \N_247\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__26331\,
            I => \N_247\
        );

    \I__5428\ : Odrv4
    port map (
            O => \N__26328\,
            I => \N_247\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__26325\,
            I => \N_247\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__26322\,
            I => \N_247\
        );

    \I__5425\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__26306\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_2\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__26303\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_1_cascade_\
        );

    \I__5422\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26297\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__26297\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_4\
        );

    \I__5420\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26288\
        );

    \I__5419\ : InMux
    port map (
            O => \N__26293\,
            I => \N__26288\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__26288\,
            I => \POWERLED.func_state_RNI_0Z0Z_1\
        );

    \I__5417\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26282\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__26282\,
            I => \N__26277\
        );

    \I__5415\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26272\
        );

    \I__5414\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26269\
        );

    \I__5413\ : Span4Mux_v
    port map (
            O => \N__26277\,
            I => \N__26266\
        );

    \I__5412\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26261\
        );

    \I__5411\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26261\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__26272\,
            I => \N__26256\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__26269\,
            I => \N__26256\
        );

    \I__5408\ : Span4Mux_v
    port map (
            O => \N__26266\,
            I => \N__26253\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26250\
        );

    \I__5406\ : Span4Mux_h
    port map (
            O => \N__26256\,
            I => \N__26247\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__26253\,
            I => \func_state_RNI_4_1\
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__26250\,
            I => \func_state_RNI_4_1\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__26247\,
            I => \func_state_RNI_4_1\
        );

    \I__5402\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26236\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__26239\,
            I => \N__26232\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__26236\,
            I => \N__26227\
        );

    \I__5399\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26224\
        );

    \I__5398\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26219\
        );

    \I__5397\ : InMux
    port map (
            O => \N__26231\,
            I => \N__26219\
        );

    \I__5396\ : InMux
    port map (
            O => \N__26230\,
            I => \N__26216\
        );

    \I__5395\ : Span4Mux_h
    port map (
            O => \N__26227\,
            I => \N__26213\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__26224\,
            I => \N__26210\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__26219\,
            I => \N__26205\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__26216\,
            I => \N__26205\
        );

    \I__5391\ : Span4Mux_s1_h
    port map (
            O => \N__26213\,
            I => \N__26200\
        );

    \I__5390\ : Span4Mux_h
    port map (
            O => \N__26210\,
            I => \N__26200\
        );

    \I__5389\ : Span4Mux_v
    port map (
            O => \N__26205\,
            I => \N__26197\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__26200\,
            I => \func_state_RNI_0_0\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__26197\,
            I => \func_state_RNI_0_0\
        );

    \I__5386\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26186\
        );

    \I__5385\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26186\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__26186\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_0\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__26183\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_0_cascade_\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__26180\,
            I => \N__26176\
        );

    \I__5381\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26171\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26164\
        );

    \I__5379\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26164\
        );

    \I__5378\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26164\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26161\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26164\,
            I => \N__26158\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__26161\,
            I => \N__26155\
        );

    \I__5374\ : Span4Mux_s3_h
    port map (
            O => \N__26158\,
            I => \N__26152\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__26155\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__26152\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__5371\ : CascadeMux
    port map (
            O => \N__26147\,
            I => \POWERLED.N_668_cascade_\
        );

    \I__5370\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26141\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__26141\,
            I => \N__26138\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__26138\,
            I => \POWERLED.N_490\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__26135\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_\
        );

    \I__5366\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26114\
        );

    \I__5365\ : InMux
    port map (
            O => \N__26131\,
            I => \N__26114\
        );

    \I__5364\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26107\
        );

    \I__5363\ : InMux
    port map (
            O => \N__26129\,
            I => \N__26107\
        );

    \I__5362\ : InMux
    port map (
            O => \N__26128\,
            I => \N__26107\
        );

    \I__5361\ : InMux
    port map (
            O => \N__26127\,
            I => \N__26102\
        );

    \I__5360\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26102\
        );

    \I__5359\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26087\
        );

    \I__5358\ : InMux
    port map (
            O => \N__26124\,
            I => \N__26087\
        );

    \I__5357\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26087\
        );

    \I__5356\ : InMux
    port map (
            O => \N__26122\,
            I => \N__26087\
        );

    \I__5355\ : InMux
    port map (
            O => \N__26121\,
            I => \N__26080\
        );

    \I__5354\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26080\
        );

    \I__5353\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26080\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__26114\,
            I => \N__26077\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26072\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26072\
        );

    \I__5349\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26059\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26100\,
            I => \N__26059\
        );

    \I__5347\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26059\
        );

    \I__5346\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26059\
        );

    \I__5345\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26059\
        );

    \I__5344\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26059\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__26087\,
            I => \N__26056\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__26080\,
            I => \N__26053\
        );

    \I__5341\ : Span4Mux_s2_v
    port map (
            O => \N__26077\,
            I => \N__26046\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__26072\,
            I => \N__26046\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__26059\,
            I => \N__26046\
        );

    \I__5338\ : Span4Mux_v
    port map (
            O => \N__26056\,
            I => \N__26041\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__26053\,
            I => \N__26041\
        );

    \I__5336\ : Span4Mux_v
    port map (
            O => \N__26046\,
            I => \N__26038\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__26041\,
            I => \POWERLED.N_123\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__26038\,
            I => \POWERLED.N_123\
        );

    \I__5333\ : InMux
    port map (
            O => \N__26033\,
            I => \N__26030\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__26030\,
            I => \N__26026\
        );

    \I__5331\ : InMux
    port map (
            O => \N__26029\,
            I => \N__26023\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__26026\,
            I => \N__26020\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__26023\,
            I => \POWERLED.N_443\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__26020\,
            I => \POWERLED.N_443\
        );

    \I__5327\ : CascadeMux
    port map (
            O => \N__26015\,
            I => \N__26011\
        );

    \I__5326\ : CascadeMux
    port map (
            O => \N__26014\,
            I => \N__26007\
        );

    \I__5325\ : InMux
    port map (
            O => \N__26011\,
            I => \N__26004\
        );

    \I__5324\ : InMux
    port map (
            O => \N__26010\,
            I => \N__25999\
        );

    \I__5323\ : InMux
    port map (
            O => \N__26007\,
            I => \N__25999\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__26004\,
            I => \N__25996\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__25999\,
            I => \N__25991\
        );

    \I__5320\ : Span4Mux_h
    port map (
            O => \N__25996\,
            I => \N__25991\
        );

    \I__5319\ : Odrv4
    port map (
            O => \N__25991\,
            I => \POWERLED.count_off_RNIH9TEZ0Z_10\
        );

    \I__5318\ : InMux
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__25985\,
            I => \N__25982\
        );

    \I__5316\ : Odrv12
    port map (
            O => \N__25982\,
            I => \POWERLED.un1_func_state25_6_0_0_0_2_1\
        );

    \I__5315\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25973\
        );

    \I__5314\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25973\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__25973\,
            I => \POWERLED.N_668\
        );

    \I__5312\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25966\
        );

    \I__5311\ : CascadeMux
    port map (
            O => \N__25969\,
            I => \N__25963\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__25966\,
            I => \N__25960\
        );

    \I__5309\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25957\
        );

    \I__5308\ : Span12Mux_s3_h
    port map (
            O => \N__25960\,
            I => \N__25954\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25951\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__25954\,
            I => \POWERLED.count_off_1_sqmuxa\
        );

    \I__5305\ : Odrv12
    port map (
            O => \N__25951\,
            I => \POWERLED.count_off_1_sqmuxa\
        );

    \I__5304\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25943\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__25940\,
            I => \POWERLED.un1_dutycycle_172_m0\
        );

    \I__5301\ : CascadeMux
    port map (
            O => \N__25937\,
            I => \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_\
        );

    \I__5300\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25931\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__25931\,
            I => \N__25928\
        );

    \I__5298\ : Span4Mux_v
    port map (
            O => \N__25928\,
            I => \N__25925\
        );

    \I__5297\ : Odrv4
    port map (
            O => \N__25925\,
            I => \POWERLED.un1_dutycycle_172_m1\
        );

    \I__5296\ : CascadeMux
    port map (
            O => \N__25922\,
            I => \N__25918\
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__25921\,
            I => \N__25915\
        );

    \I__5294\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25912\
        );

    \I__5293\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25909\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25904\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__25909\,
            I => \N__25904\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__25904\,
            I => \N__25901\
        );

    \I__5289\ : Odrv4
    port map (
            O => \N__25901\,
            I => \POWERLED.func_state_RNI_3Z0Z_1\
        );

    \I__5288\ : CascadeMux
    port map (
            O => \N__25898\,
            I => \POWERLED.count_clk_RNIZ0Z_0_cascade_\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__25895\,
            I => \POWERLED.count_clkZ0Z_1_cascade_\
        );

    \I__5286\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25889\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__25889\,
            I => \POWERLED.count_clk_0_1\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__25886\,
            I => \N__25883\
        );

    \I__5283\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25880\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__25880\,
            I => \N__25877\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__25877\,
            I => \POWERLED.count_clk_0_11\
        );

    \I__5280\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25868\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__25873\,
            I => \N__25861\
        );

    \I__5278\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25858\
        );

    \I__5277\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25855\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__25868\,
            I => \N__25852\
        );

    \I__5275\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25847\
        );

    \I__5274\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25847\
        );

    \I__5273\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25844\
        );

    \I__5272\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25839\
        );

    \I__5271\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25839\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25836\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25833\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__25852\,
            I => \N__25830\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__25847\,
            I => \N__25823\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__25844\,
            I => \N__25823\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__25839\,
            I => \N__25823\
        );

    \I__5264\ : Span4Mux_s2_h
    port map (
            O => \N__25836\,
            I => \N__25820\
        );

    \I__5263\ : Span4Mux_s2_h
    port map (
            O => \N__25833\,
            I => \N__25817\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__25830\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__5261\ : Odrv4
    port map (
            O => \N__25823\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__25820\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__25817\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__25808\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3_cascade_\
        );

    \I__5257\ : SRMux
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25797\
        );

    \I__5255\ : SRMux
    port map (
            O => \N__25801\,
            I => \N__25794\
        );

    \I__5254\ : SRMux
    port map (
            O => \N__25800\,
            I => \N__25791\
        );

    \I__5253\ : Span4Mux_v
    port map (
            O => \N__25797\,
            I => \N__25786\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__25794\,
            I => \N__25786\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__25791\,
            I => \N__25783\
        );

    \I__5250\ : Span4Mux_s2_v
    port map (
            O => \N__25786\,
            I => \N__25778\
        );

    \I__5249\ : Span4Mux_s1_h
    port map (
            O => \N__25783\,
            I => \N__25778\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__25778\,
            I => \G_30\
        );

    \I__5247\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__25772\,
            I => \POWERLED.count_clk_0_4\
        );

    \I__5245\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__25766\,
            I => \POWERLED.count_clk_0_5\
        );

    \I__5243\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25760\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__25760\,
            I => \POWERLED.count_clk_0_6\
        );

    \I__5241\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25727\
        );

    \I__5240\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25727\
        );

    \I__5239\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25718\
        );

    \I__5238\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25718\
        );

    \I__5237\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25718\
        );

    \I__5236\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25718\
        );

    \I__5235\ : InMux
    port map (
            O => \N__25751\,
            I => \N__25709\
        );

    \I__5234\ : InMux
    port map (
            O => \N__25750\,
            I => \N__25709\
        );

    \I__5233\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25709\
        );

    \I__5232\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25709\
        );

    \I__5231\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25702\
        );

    \I__5230\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25702\
        );

    \I__5229\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25702\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__25744\,
            I => \N__25699\
        );

    \I__5227\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25694\
        );

    \I__5226\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25687\
        );

    \I__5225\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25687\
        );

    \I__5224\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25687\
        );

    \I__5223\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25684\
        );

    \I__5222\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25673\
        );

    \I__5221\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25673\
        );

    \I__5220\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25673\
        );

    \I__5219\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25673\
        );

    \I__5218\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25673\
        );

    \I__5217\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25668\
        );

    \I__5216\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25668\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__25727\,
            I => \N__25659\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__25718\,
            I => \N__25659\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25659\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__25702\,
            I => \N__25659\
        );

    \I__5211\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25648\
        );

    \I__5210\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25648\
        );

    \I__5209\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25648\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__25694\,
            I => \N__25635\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__25687\,
            I => \N__25635\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__25684\,
            I => \N__25635\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25635\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__25668\,
            I => \N__25635\
        );

    \I__5203\ : Span4Mux_v
    port map (
            O => \N__25659\,
            I => \N__25635\
        );

    \I__5202\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25631\
        );

    \I__5201\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25624\
        );

    \I__5200\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25624\
        );

    \I__5199\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25624\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__25648\,
            I => \N__25621\
        );

    \I__5197\ : Span4Mux_v
    port map (
            O => \N__25635\,
            I => \N__25616\
        );

    \I__5196\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25613\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__25631\,
            I => \N__25610\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__25624\,
            I => \N__25605\
        );

    \I__5193\ : Span12Mux_s6_h
    port map (
            O => \N__25621\,
            I => \N__25605\
        );

    \I__5192\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25600\
        );

    \I__5191\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25600\
        );

    \I__5190\ : Sp12to4
    port map (
            O => \N__25616\,
            I => \N__25595\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__25613\,
            I => \N__25595\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__25610\,
            I => \clk_100Khz_signalkeep_3\
        );

    \I__5187\ : Odrv12
    port map (
            O => \N__25605\,
            I => \clk_100Khz_signalkeep_3\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__25600\,
            I => \clk_100Khz_signalkeep_3\
        );

    \I__5185\ : Odrv12
    port map (
            O => \N__25595\,
            I => \clk_100Khz_signalkeep_3\
        );

    \I__5184\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25583\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__25583\,
            I => \N__25574\
        );

    \I__5182\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25569\
        );

    \I__5181\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25569\
        );

    \I__5180\ : InMux
    port map (
            O => \N__25580\,
            I => \N__25566\
        );

    \I__5179\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25561\
        );

    \I__5178\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25561\
        );

    \I__5177\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25558\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__25574\,
            I => \N__25553\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__25569\,
            I => \N__25553\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__25566\,
            I => \clk_100Khz_signalkeep_3_rep1\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__25561\,
            I => \clk_100Khz_signalkeep_3_rep1\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__25558\,
            I => \clk_100Khz_signalkeep_3_rep1\
        );

    \I__5171\ : Odrv4
    port map (
            O => \N__25553\,
            I => \clk_100Khz_signalkeep_3_rep1\
        );

    \I__5170\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25540\
        );

    \I__5169\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25537\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__25540\,
            I => \N__25534\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__25537\,
            I => \N__25529\
        );

    \I__5166\ : Span4Mux_s2_v
    port map (
            O => \N__25534\,
            I => \N__25529\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__25529\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__5164\ : InMux
    port map (
            O => \N__25526\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__5162\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25513\
        );

    \I__5160\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25510\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__25513\,
            I => \N__25507\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__25510\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__25507\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__5156\ : InMux
    port map (
            O => \N__25502\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__25499\,
            I => \N__25496\
        );

    \I__5154\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25493\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__25493\,
            I => \N__25489\
        );

    \I__5152\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25486\
        );

    \I__5151\ : Span4Mux_s2_v
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__25486\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__5149\ : Odrv4
    port map (
            O => \N__25483\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__5148\ : InMux
    port map (
            O => \N__25478\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__5147\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25472\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__25472\,
            I => \N__25468\
        );

    \I__5145\ : InMux
    port map (
            O => \N__25471\,
            I => \N__25465\
        );

    \I__5144\ : Span4Mux_s2_v
    port map (
            O => \N__25468\,
            I => \N__25462\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__25465\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__25462\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__5141\ : InMux
    port map (
            O => \N__25457\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__5140\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25451\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25447\
        );

    \I__5138\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25444\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__25447\,
            I => \N__25441\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__25444\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__25441\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__5134\ : InMux
    port map (
            O => \N__25436\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__5133\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25390\
        );

    \I__5132\ : InMux
    port map (
            O => \N__25432\,
            I => \N__25390\
        );

    \I__5131\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25390\
        );

    \I__5130\ : InMux
    port map (
            O => \N__25430\,
            I => \N__25390\
        );

    \I__5129\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25381\
        );

    \I__5128\ : InMux
    port map (
            O => \N__25428\,
            I => \N__25381\
        );

    \I__5127\ : InMux
    port map (
            O => \N__25427\,
            I => \N__25381\
        );

    \I__5126\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25381\
        );

    \I__5125\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25372\
        );

    \I__5124\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25372\
        );

    \I__5123\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25372\
        );

    \I__5122\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25372\
        );

    \I__5121\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25363\
        );

    \I__5120\ : InMux
    port map (
            O => \N__25420\,
            I => \N__25363\
        );

    \I__5119\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25363\
        );

    \I__5118\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25363\
        );

    \I__5117\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25356\
        );

    \I__5116\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25356\
        );

    \I__5115\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25356\
        );

    \I__5114\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25347\
        );

    \I__5113\ : InMux
    port map (
            O => \N__25413\,
            I => \N__25347\
        );

    \I__5112\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25347\
        );

    \I__5111\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25347\
        );

    \I__5110\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25340\
        );

    \I__5109\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25340\
        );

    \I__5108\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25340\
        );

    \I__5107\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25331\
        );

    \I__5106\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25331\
        );

    \I__5105\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25331\
        );

    \I__5104\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25331\
        );

    \I__5103\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25328\
        );

    \I__5102\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25325\
        );

    \I__5101\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25320\
        );

    \I__5100\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25320\
        );

    \I__5099\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25317\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25305\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__25381\,
            I => \N__25302\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__25372\,
            I => \N__25299\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__25363\,
            I => \N__25296\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__25356\,
            I => \N__25293\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25290\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__25340\,
            I => \N__25287\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__25331\,
            I => \N__25284\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__25328\,
            I => \N__25281\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__25325\,
            I => \N__25278\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__25320\,
            I => \N__25275\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25272\
        );

    \I__5086\ : CEMux
    port map (
            O => \N__25316\,
            I => \N__25229\
        );

    \I__5085\ : CEMux
    port map (
            O => \N__25315\,
            I => \N__25229\
        );

    \I__5084\ : CEMux
    port map (
            O => \N__25314\,
            I => \N__25229\
        );

    \I__5083\ : CEMux
    port map (
            O => \N__25313\,
            I => \N__25229\
        );

    \I__5082\ : CEMux
    port map (
            O => \N__25312\,
            I => \N__25229\
        );

    \I__5081\ : CEMux
    port map (
            O => \N__25311\,
            I => \N__25229\
        );

    \I__5080\ : CEMux
    port map (
            O => \N__25310\,
            I => \N__25229\
        );

    \I__5079\ : CEMux
    port map (
            O => \N__25309\,
            I => \N__25229\
        );

    \I__5078\ : CEMux
    port map (
            O => \N__25308\,
            I => \N__25229\
        );

    \I__5077\ : Glb2LocalMux
    port map (
            O => \N__25305\,
            I => \N__25229\
        );

    \I__5076\ : Glb2LocalMux
    port map (
            O => \N__25302\,
            I => \N__25229\
        );

    \I__5075\ : Glb2LocalMux
    port map (
            O => \N__25299\,
            I => \N__25229\
        );

    \I__5074\ : Glb2LocalMux
    port map (
            O => \N__25296\,
            I => \N__25229\
        );

    \I__5073\ : Glb2LocalMux
    port map (
            O => \N__25293\,
            I => \N__25229\
        );

    \I__5072\ : Glb2LocalMux
    port map (
            O => \N__25290\,
            I => \N__25229\
        );

    \I__5071\ : Glb2LocalMux
    port map (
            O => \N__25287\,
            I => \N__25229\
        );

    \I__5070\ : Glb2LocalMux
    port map (
            O => \N__25284\,
            I => \N__25229\
        );

    \I__5069\ : Glb2LocalMux
    port map (
            O => \N__25281\,
            I => \N__25229\
        );

    \I__5068\ : Glb2LocalMux
    port map (
            O => \N__25278\,
            I => \N__25229\
        );

    \I__5067\ : Glb2LocalMux
    port map (
            O => \N__25275\,
            I => \N__25229\
        );

    \I__5066\ : Glb2LocalMux
    port map (
            O => \N__25272\,
            I => \N__25229\
        );

    \I__5065\ : GlobalMux
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__5064\ : gio2CtrlBuf
    port map (
            O => \N__25226\,
            I => \N_92_g\
        );

    \I__5063\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25219\
        );

    \I__5062\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25216\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__25219\,
            I => \N__25213\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__25216\,
            I => \N__25208\
        );

    \I__5059\ : Span4Mux_s2_v
    port map (
            O => \N__25213\,
            I => \N__25208\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__25208\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__5057\ : InMux
    port map (
            O => \N__25205\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__5056\ : IoInMux
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__5054\ : IoSpan4Mux
    port map (
            O => \N__25196\,
            I => \N__25190\
        );

    \I__5053\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25187\
        );

    \I__5052\ : InMux
    port map (
            O => \N__25194\,
            I => \N__25184\
        );

    \I__5051\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25177\
        );

    \I__5050\ : IoSpan4Mux
    port map (
            O => \N__25190\,
            I => \N__25174\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25169\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__25184\,
            I => \N__25169\
        );

    \I__5047\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25166\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25163\
        );

    \I__5045\ : IoInMux
    port map (
            O => \N__25181\,
            I => \N__25160\
        );

    \I__5044\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25157\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25154\
        );

    \I__5042\ : Span4Mux_s0_h
    port map (
            O => \N__25174\,
            I => \N__25151\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__25169\,
            I => \N__25148\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25143\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__25163\,
            I => \N__25143\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__25160\,
            I => \N__25140\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__25157\,
            I => \N__25137\
        );

    \I__5036\ : Span12Mux_s2_h
    port map (
            O => \N__25154\,
            I => \N__25134\
        );

    \I__5035\ : Span4Mux_h
    port map (
            O => \N__25151\,
            I => \N__25127\
        );

    \I__5034\ : Span4Mux_s2_v
    port map (
            O => \N__25148\,
            I => \N__25127\
        );

    \I__5033\ : Span4Mux_v
    port map (
            O => \N__25143\,
            I => \N__25127\
        );

    \I__5032\ : IoSpan4Mux
    port map (
            O => \N__25140\,
            I => \N__25124\
        );

    \I__5031\ : Span12Mux_v
    port map (
            O => \N__25137\,
            I => \N__25121\
        );

    \I__5030\ : Span12Mux_v
    port map (
            O => \N__25134\,
            I => \N__25118\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__25127\,
            I => \N__25113\
        );

    \I__5028\ : IoSpan4Mux
    port map (
            O => \N__25124\,
            I => \N__25113\
        );

    \I__5027\ : Odrv12
    port map (
            O => \N__25121\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5026\ : Odrv12
    port map (
            O => \N__25118\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__25113\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5024\ : InMux
    port map (
            O => \N__25106\,
            I => \bfn_11_4_0_\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__25103\,
            I => \N__25100\
        );

    \I__5022\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25097\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__25097\,
            I => \N__25093\
        );

    \I__5020\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25090\
        );

    \I__5019\ : Span4Mux_h
    port map (
            O => \N__25093\,
            I => \N__25087\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__25090\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__25087\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__5016\ : CEMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__5014\ : Span4Mux_s2_h
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__5013\ : Odrv4
    port map (
            O => \N__25073\,
            I => \VPP_VDDQ.N_92_0\
        );

    \I__5012\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25066\
        );

    \I__5011\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25063\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__25063\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__25060\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__5007\ : InMux
    port map (
            O => \N__25055\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__5006\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25048\
        );

    \I__5005\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25045\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__25048\,
            I => \N__25042\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__25045\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__25042\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__5001\ : InMux
    port map (
            O => \N__25037\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__5000\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25030\
        );

    \I__4999\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25027\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__25024\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25027\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__25024\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4995\ : InMux
    port map (
            O => \N__25019\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__4994\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25012\
        );

    \I__4993\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__25012\,
            I => \N__25006\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__25009\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__25006\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4989\ : InMux
    port map (
            O => \N__25001\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__4988\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24994\
        );

    \I__4987\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24991\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__24994\,
            I => \N__24988\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__24991\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__24988\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__4983\ : InMux
    port map (
            O => \N__24983\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__4982\ : InMux
    port map (
            O => \N__24980\,
            I => \N__24976\
        );

    \I__4981\ : InMux
    port map (
            O => \N__24979\,
            I => \N__24973\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__24976\,
            I => \N__24970\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__24973\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__4978\ : Odrv12
    port map (
            O => \N__24970\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__4977\ : InMux
    port map (
            O => \N__24965\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__4975\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24955\
        );

    \I__4974\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24952\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__24955\,
            I => \N__24949\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__24952\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__24949\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4970\ : InMux
    port map (
            O => \N__24944\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__4969\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24937\
        );

    \I__4968\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24934\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__24937\,
            I => \N__24931\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__24934\,
            I => \N__24926\
        );

    \I__4965\ : Span4Mux_s2_v
    port map (
            O => \N__24931\,
            I => \N__24926\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__24926\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__4963\ : InMux
    port map (
            O => \N__24923\,
            I => \bfn_11_3_0_\
        );

    \I__4962\ : InMux
    port map (
            O => \N__24920\,
            I => \N__24914\
        );

    \I__4961\ : InMux
    port map (
            O => \N__24919\,
            I => \N__24914\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__24914\,
            I => \N__24911\
        );

    \I__4959\ : Odrv12
    port map (
            O => \N__24911\,
            I => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__24908\,
            I => \N__24905\
        );

    \I__4957\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24899\
        );

    \I__4956\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24899\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__4954\ : Span12Mux_s5_h
    port map (
            O => \N__24896\,
            I => \N__24893\
        );

    \I__4953\ : Odrv12
    port map (
            O => \N__24893\,
            I => \POWERLED.dutycycle_en_4\
        );

    \I__4952\ : CascadeMux
    port map (
            O => \N__24890\,
            I => \N__24887\
        );

    \I__4951\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24881\
        );

    \I__4950\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24881\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__24881\,
            I => \POWERLED.dutycycleZ1Z_10\
        );

    \I__4948\ : CascadeMux
    port map (
            O => \N__24878\,
            I => \POWERLED.dutycycleZ0Z_2_cascade_\
        );

    \I__4947\ : InMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__24869\,
            I => \POWERLED.un2_count_clk_17_0_0_a2_0_0\
        );

    \I__4944\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__24863\,
            I => \POWERLED.un1_dutycycle_53_50_0_0\
        );

    \I__4942\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24853\
        );

    \I__4941\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24850\
        );

    \I__4940\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24843\
        );

    \I__4939\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24843\
        );

    \I__4938\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24843\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__24853\,
            I => \N__24840\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__24850\,
            I => \POWERLED.un1_dutycycle_53_4_0\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__24843\,
            I => \POWERLED.un1_dutycycle_53_4_0\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__24840\,
            I => \POWERLED.un1_dutycycle_53_4_0\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__24833\,
            I => \POWERLED.un1_dutycycle_53_10_2_cascade_\
        );

    \I__4932\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24827\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__24827\,
            I => \N__24824\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__24824\,
            I => \POWERLED.un1_dutycycle_53_10_3\
        );

    \I__4929\ : InMux
    port map (
            O => \N__24821\,
            I => \N__24818\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__24818\,
            I => \POWERLED.un1_dutycycle_53_9_a1_0\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \N__24810\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__24814\,
            I => \N__24806\
        );

    \I__4925\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24803\
        );

    \I__4924\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24800\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__24809\,
            I => \N__24797\
        );

    \I__4922\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24790\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__24803\,
            I => \N__24785\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__24800\,
            I => \N__24785\
        );

    \I__4919\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24782\
        );

    \I__4918\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24779\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__24795\,
            I => \N__24774\
        );

    \I__4916\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24771\
        );

    \I__4915\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24768\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__24790\,
            I => \N__24762\
        );

    \I__4913\ : Span4Mux_h
    port map (
            O => \N__24785\,
            I => \N__24762\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__24782\,
            I => \N__24757\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24757\
        );

    \I__4910\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24750\
        );

    \I__4909\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24750\
        );

    \I__4908\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24750\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__24771\,
            I => \N__24743\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__24768\,
            I => \N__24740\
        );

    \I__4905\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24737\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__24762\,
            I => \N__24732\
        );

    \I__4903\ : Span4Mux_h
    port map (
            O => \N__24757\,
            I => \N__24732\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24729\
        );

    \I__4901\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24720\
        );

    \I__4900\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24720\
        );

    \I__4899\ : InMux
    port map (
            O => \N__24747\,
            I => \N__24720\
        );

    \I__4898\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24720\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__24743\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4896\ : Odrv12
    port map (
            O => \N__24740\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__24737\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4894\ : Odrv4
    port map (
            O => \N__24732\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__24729\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__24720\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__24707\,
            I => \N__24697\
        );

    \I__4890\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24692\
        );

    \I__4889\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24689\
        );

    \I__4888\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24682\
        );

    \I__4887\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24682\
        );

    \I__4886\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24682\
        );

    \I__4885\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24679\
        );

    \I__4884\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24673\
        );

    \I__4883\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24670\
        );

    \I__4882\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24665\
        );

    \I__4881\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24665\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__24692\,
            I => \N__24660\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__24689\,
            I => \N__24660\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__24682\,
            I => \N__24657\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__24679\,
            I => \N__24654\
        );

    \I__4876\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24649\
        );

    \I__4875\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24649\
        );

    \I__4874\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24646\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__24673\,
            I => \N__24637\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__24670\,
            I => \N__24637\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__24665\,
            I => \N__24637\
        );

    \I__4870\ : Span4Mux_v
    port map (
            O => \N__24660\,
            I => \N__24637\
        );

    \I__4869\ : Span4Mux_v
    port map (
            O => \N__24657\,
            I => \N__24634\
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__24654\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__24649\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__24646\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4865\ : Odrv4
    port map (
            O => \N__24637\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__24634\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4863\ : CascadeMux
    port map (
            O => \N__24623\,
            I => \N__24620\
        );

    \I__4862\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24615\
        );

    \I__4861\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24609\
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__24618\,
            I => \N__24600\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__24615\,
            I => \N__24596\
        );

    \I__4858\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24591\
        );

    \I__4857\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24591\
        );

    \I__4856\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24588\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24585\
        );

    \I__4854\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24582\
        );

    \I__4853\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24579\
        );

    \I__4852\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24574\
        );

    \I__4851\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24574\
        );

    \I__4850\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24569\
        );

    \I__4849\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24569\
        );

    \I__4848\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24564\
        );

    \I__4847\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24564\
        );

    \I__4846\ : Span4Mux_h
    port map (
            O => \N__24596\,
            I => \N__24557\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__24591\,
            I => \N__24557\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24557\
        );

    \I__4843\ : Odrv4
    port map (
            O => \N__24585\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__24582\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__24579\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__24574\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__24569\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__24564\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__24557\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4836\ : CascadeMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__4835\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__24536\,
            I => \POWERLED.un1_dutycycle_53_50_3_0\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__24533\,
            I => \N__24529\
        );

    \I__4832\ : InMux
    port map (
            O => \N__24532\,
            I => \N__24526\
        );

    \I__4831\ : InMux
    port map (
            O => \N__24529\,
            I => \N__24523\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__24526\,
            I => \N__24520\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__24523\,
            I => \N__24517\
        );

    \I__4828\ : Span4Mux_s2_v
    port map (
            O => \N__24520\,
            I => \N__24512\
        );

    \I__4827\ : Span4Mux_s2_v
    port map (
            O => \N__24517\,
            I => \N__24512\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__24512\,
            I => \VPP_VDDQ.N_64_i\
        );

    \I__4825\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24505\
        );

    \I__4824\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24502\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__24505\,
            I => \N__24499\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__24502\,
            I => \N__24494\
        );

    \I__4821\ : Span4Mux_s1_v
    port map (
            O => \N__24499\,
            I => \N__24494\
        );

    \I__4820\ : Odrv4
    port map (
            O => \N__24494\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__4819\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__24488\,
            I => \POWERLED.un1_dutycycle_53_45_0\
        );

    \I__4817\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__24479\,
            I => \POWERLED.dutycycle_RNIZ0Z_4\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__24476\,
            I => \POWERLED.un1_dutycycle_53_35_1_cascade_\
        );

    \I__4813\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24469\
        );

    \I__4812\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24464\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__24469\,
            I => \N__24461\
        );

    \I__4810\ : InMux
    port map (
            O => \N__24468\,
            I => \N__24456\
        );

    \I__4809\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24456\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__24464\,
            I => \POWERLED.un1_dutycycle_53_22\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__24461\,
            I => \POWERLED.un1_dutycycle_53_22\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__24456\,
            I => \POWERLED.un1_dutycycle_53_22\
        );

    \I__4805\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__24446\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_6\
        );

    \I__4803\ : InMux
    port map (
            O => \N__24443\,
            I => \N__24438\
        );

    \I__4802\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24435\
        );

    \I__4801\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24431\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__24438\,
            I => \N__24428\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__24435\,
            I => \N__24422\
        );

    \I__4798\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24419\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__24431\,
            I => \N__24416\
        );

    \I__4796\ : Span4Mux_s3_v
    port map (
            O => \N__24428\,
            I => \N__24413\
        );

    \I__4795\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24410\
        );

    \I__4794\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24407\
        );

    \I__4793\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24404\
        );

    \I__4792\ : Span4Mux_s1_v
    port map (
            O => \N__24422\,
            I => \N__24397\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__24419\,
            I => \N__24397\
        );

    \I__4790\ : Span4Mux_h
    port map (
            O => \N__24416\,
            I => \N__24397\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__24413\,
            I => \POWERLED.dutycycle_RNI_10_8\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__24410\,
            I => \POWERLED.dutycycle_RNI_10_8\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__24407\,
            I => \POWERLED.dutycycle_RNI_10_8\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__24404\,
            I => \POWERLED.dutycycle_RNI_10_8\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__24397\,
            I => \POWERLED.dutycycle_RNI_10_8\
        );

    \I__4784\ : InMux
    port map (
            O => \N__24386\,
            I => \N__24383\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__24383\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__24380\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_\
        );

    \I__4781\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24371\
        );

    \I__4780\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24371\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__24371\,
            I => \POWERLED.un1_dutycycle_53_35_1\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__4777\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24361\
        );

    \I__4776\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24358\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__24361\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_6\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__24358\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_6\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__24353\,
            I => \N__24350\
        );

    \I__4772\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24345\
        );

    \I__4771\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24340\
        );

    \I__4770\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24340\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__24345\,
            I => \POWERLED.un1_dutycycle_53_50_a0_0\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__24340\,
            I => \POWERLED.un1_dutycycle_53_50_a0_0\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__24335\,
            I => \POWERLED.un1_dutycycle_53_50_a0_0_cascade_\
        );

    \I__4766\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__24329\,
            I => \POWERLED.un1_dutycycle_53_50_a0_0_0\
        );

    \I__4764\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24323\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__24323\,
            I => \POWERLED.un1_dutycycle_53_9_4_0\
        );

    \I__4762\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__24317\,
            I => \POWERLED.un1_dutycycle_53_9_4_1\
        );

    \I__4760\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24310\
        );

    \I__4759\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24307\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__24310\,
            I => \N__24302\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__24307\,
            I => \N__24302\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__24302\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__24299\,
            I => \N__24295\
        );

    \I__4754\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24290\
        );

    \I__4753\ : InMux
    port map (
            O => \N__24295\,
            I => \N__24290\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__24287\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__24284\,
            I => \POWERLED.dutycycleZ0Z_7_cascade_\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__24281\,
            I => \POWERLED.un1_dutycycle_53_9_a0_0_cascade_\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__24278\,
            I => \N__24275\
        );

    \I__4747\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__24269\,
            I => \POWERLED.un1_dutycycle_53_10_4\
        );

    \I__4744\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__24263\,
            I => \POWERLED.un1_dutycycle_53_40_0\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__24260\,
            I => \POWERLED.un1_dutycycle_53_axb_11_1_cascade_\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__24257\,
            I => \POWERLED.un1_dutycycle_53_axb_11_cascade_\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__24254\,
            I => \N__24251\
        );

    \I__4739\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__4737\ : Odrv4
    port map (
            O => \N__24245\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_14\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__24242\,
            I => \POWERLED.dutycycleZ0Z_5_cascade_\
        );

    \I__4735\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__24236\,
            I => \POWERLED.dutycycle_RNIF86R3Z0Z_4\
        );

    \I__4733\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24230\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__24230\,
            I => \POWERLED.dutycycle_RNIP1UTZ0Z_4\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__24227\,
            I => \POWERLED.dutycycle_RNIF86R3Z0Z_4_cascade_\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24215\
        );

    \I__4729\ : InMux
    port map (
            O => \N__24223\,
            I => \N__24215\
        );

    \I__4728\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24215\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__24215\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__24212\,
            I => \POWERLED.un1_dutycycle_53_31_0_0_cascade_\
        );

    \I__4725\ : InMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__24206\,
            I => \POWERLED.un1_dutycycle_53_9_3\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__24203\,
            I => \N__24200\
        );

    \I__4722\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__24191\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_11\
        );

    \I__4718\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24182\
        );

    \I__4717\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24182\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__24182\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__4714\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24170\
        );

    \I__4713\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24170\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24167\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__24167\,
            I => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\
        );

    \I__4710\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24158\
        );

    \I__4709\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24158\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__24158\,
            I => \N__24155\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__24155\,
            I => \N__24152\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__24152\,
            I => \POWERLED.dutycycle_RNIRT5H5Z0Z_8\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__24149\,
            I => \POWERLED.dutycycleZ0Z_3_cascade_\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__24146\,
            I => \POWERLED.dutycycle_RNI_10_8_cascade_\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24140\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__24140\,
            I => \POWERLED.un1_dutycycle_53_9_4\
        );

    \I__4701\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24131\
        );

    \I__4700\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24131\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__24131\,
            I => \N__24128\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__24128\,
            I => \N__24125\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__24125\,
            I => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\
        );

    \I__4696\ : InMux
    port map (
            O => \N__24122\,
            I => \POWERLED.un1_dutycycle_94_cry_10\
        );

    \I__4695\ : InMux
    port map (
            O => \N__24119\,
            I => \POWERLED.un1_dutycycle_94_cry_11_cZ0\
        );

    \I__4694\ : InMux
    port map (
            O => \N__24116\,
            I => \N__24108\
        );

    \I__4693\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24103\
        );

    \I__4692\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24103\
        );

    \I__4691\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24098\
        );

    \I__4690\ : InMux
    port map (
            O => \N__24112\,
            I => \N__24098\
        );

    \I__4689\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24095\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24090\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__24103\,
            I => \N__24085\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__24098\,
            I => \N__24085\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__24095\,
            I => \N__24082\
        );

    \I__4684\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24079\
        );

    \I__4683\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24076\
        );

    \I__4682\ : Span4Mux_h
    port map (
            O => \N__24090\,
            I => \N__24071\
        );

    \I__4681\ : Span4Mux_s1_v
    port map (
            O => \N__24085\,
            I => \N__24071\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__24082\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__24079\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__24076\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__24071\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4676\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24056\
        );

    \I__4675\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24056\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__24056\,
            I => \N__24053\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__24053\,
            I => \N__24050\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__24050\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\
        );

    \I__4671\ : InMux
    port map (
            O => \N__24047\,
            I => \POWERLED.un1_dutycycle_94_cry_12\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__24044\,
            I => \N__24033\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__24043\,
            I => \N__24030\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__24042\,
            I => \N__24026\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__24041\,
            I => \N__24023\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__24040\,
            I => \N__24018\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__24039\,
            I => \N__24015\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__24038\,
            I => \N__24011\
        );

    \I__4663\ : CascadeMux
    port map (
            O => \N__24037\,
            I => \N__24007\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__24036\,
            I => \N__24004\
        );

    \I__4661\ : InMux
    port map (
            O => \N__24033\,
            I => \N__23999\
        );

    \I__4660\ : InMux
    port map (
            O => \N__24030\,
            I => \N__23999\
        );

    \I__4659\ : InMux
    port map (
            O => \N__24029\,
            I => \N__23994\
        );

    \I__4658\ : InMux
    port map (
            O => \N__24026\,
            I => \N__23994\
        );

    \I__4657\ : InMux
    port map (
            O => \N__24023\,
            I => \N__23983\
        );

    \I__4656\ : InMux
    port map (
            O => \N__24022\,
            I => \N__23983\
        );

    \I__4655\ : InMux
    port map (
            O => \N__24021\,
            I => \N__23983\
        );

    \I__4654\ : InMux
    port map (
            O => \N__24018\,
            I => \N__23983\
        );

    \I__4653\ : InMux
    port map (
            O => \N__24015\,
            I => \N__23983\
        );

    \I__4652\ : InMux
    port map (
            O => \N__24014\,
            I => \N__23972\
        );

    \I__4651\ : InMux
    port map (
            O => \N__24011\,
            I => \N__23972\
        );

    \I__4650\ : InMux
    port map (
            O => \N__24010\,
            I => \N__23972\
        );

    \I__4649\ : InMux
    port map (
            O => \N__24007\,
            I => \N__23972\
        );

    \I__4648\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23972\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23963\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__23994\,
            I => \N__23963\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23963\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__23972\,
            I => \N__23963\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__23963\,
            I => \POWERLED.N_435_i\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__23960\,
            I => \N__23957\
        );

    \I__4641\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23951\
        );

    \I__4640\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23951\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__4638\ : Span4Mux_s3_v
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__23945\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\
        );

    \I__4636\ : InMux
    port map (
            O => \N__23942\,
            I => \POWERLED.un1_dutycycle_94_cry_13_cZ0\
        );

    \I__4635\ : InMux
    port map (
            O => \N__23939\,
            I => \POWERLED.un1_dutycycle_94_cry_14\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__23936\,
            I => \N__23932\
        );

    \I__4633\ : InMux
    port map (
            O => \N__23935\,
            I => \N__23927\
        );

    \I__4632\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23927\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__4630\ : Span4Mux_s2_v
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__23921\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\
        );

    \I__4628\ : IoInMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__23915\,
            I => \N__23912\
        );

    \I__4626\ : IoSpan4Mux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__4625\ : Span4Mux_s3_h
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__4624\ : Span4Mux_h
    port map (
            O => \N__23906\,
            I => \N__23903\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__23903\,
            I => vccst_en
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__23900\,
            I => \N__23897\
        );

    \I__4621\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23894\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__23891\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__23888\,
            I => \POWERLED.dutycycle_RNIP1UTZ0Z_4_cascade_\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__23885\,
            I => \N__23882\
        );

    \I__4616\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__23879\,
            I => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\
        );

    \I__4614\ : InMux
    port map (
            O => \N__23876\,
            I => \POWERLED.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__4613\ : InMux
    port map (
            O => \N__23873\,
            I => \POWERLED.un1_dutycycle_94_cry_2_cZ0\
        );

    \I__4612\ : InMux
    port map (
            O => \N__23870\,
            I => \POWERLED.un1_dutycycle_94_cry_3_cZ0\
        );

    \I__4611\ : InMux
    port map (
            O => \N__23867\,
            I => \POWERLED.un1_dutycycle_94_cry_4\
        );

    \I__4610\ : InMux
    port map (
            O => \N__23864\,
            I => \POWERLED.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__4609\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23858\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__23858\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\
        );

    \I__4607\ : InMux
    port map (
            O => \N__23855\,
            I => \POWERLED.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__4606\ : InMux
    port map (
            O => \N__23852\,
            I => \bfn_9_11_0_\
        );

    \I__4605\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23843\
        );

    \I__4604\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23843\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__23843\,
            I => \N__23840\
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__23840\,
            I => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\
        );

    \I__4601\ : InMux
    port map (
            O => \N__23837\,
            I => \POWERLED.un1_dutycycle_94_cry_8\
        );

    \I__4600\ : InMux
    port map (
            O => \N__23834\,
            I => \POWERLED.un1_dutycycle_94_cry_9\
        );

    \I__4599\ : CascadeMux
    port map (
            O => \N__23831\,
            I => \N__23828\
        );

    \I__4598\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23825\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__23825\,
            I => \POWERLED.func_state_1_m2s2_i_0_a2_1_0\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__23822\,
            I => \POWERLED.un1_dutycycle_96_0_a3_0_a2_1_cascade_\
        );

    \I__4595\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23816\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__23816\,
            I => \N__23812\
        );

    \I__4593\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23809\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__23812\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__23809\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__23804\,
            I => \POWERLED.N_251_cascade_\
        );

    \I__4589\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23795\
        );

    \I__4587\ : Odrv4
    port map (
            O => \N__23795\,
            I => \POWERLED.N_506\
        );

    \I__4586\ : InMux
    port map (
            O => \N__23792\,
            I => \POWERLED.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__23789\,
            I => \POWERLED.N_448_cascade_\
        );

    \I__4584\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23783\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__23780\,
            I => \POWERLED.N_656_0\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__23777\,
            I => \POWERLED.N_133_cascade_\
        );

    \I__4580\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23771\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__23771\,
            I => \POWERLED.un1_dutycycle_172_m4\
        );

    \I__4578\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23765\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__23765\,
            I => \N__23762\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__23762\,
            I => \POWERLED.dutycycle_eena_14_c\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__23759\,
            I => \POWERLED.N_488_cascade_\
        );

    \I__4574\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__23753\,
            I => \POWERLED.un1_dutycycle_172_m2\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__23750\,
            I => \POWERLED.un1_clk_100khz_30_and_i_0_0_sx_cascade_\
        );

    \I__4571\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__23744\,
            I => \POWERLED.un1_dutycycle_164_0_a3_0_a2_0\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__23741\,
            I => \POWERLED.count_clkZ0Z_7_cascade_\
        );

    \I__4568\ : InMux
    port map (
            O => \N__23738\,
            I => \N__23735\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__23735\,
            I => \N__23732\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__23732\,
            I => \POWERLED.un1_func_state25_6_0_o_N_4\
        );

    \I__4565\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23723\
        );

    \I__4564\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23723\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__23723\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_9_0\
        );

    \I__4562\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23717\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__23717\,
            I => \POWERLED.count_clk_0_7\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__23714\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_\
        );

    \I__4559\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__23705\,
            I => \POWERLED.un1_dutycycle_172_m3\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__23702\,
            I => \POWERLED.un1_clk_100khz_52_and_i_0_m2_ns_1_cascade_\
        );

    \I__4555\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23696\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__23696\,
            I => \POWERLED_g2_1_0_0\
        );

    \I__4553\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23690\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__4551\ : Span4Mux_v
    port map (
            O => \N__23687\,
            I => \N__23684\
        );

    \I__4550\ : Odrv4
    port map (
            O => \N__23684\,
            I => \POWERLED.N_74\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__23681\,
            I => \POWERLED.N_4_0_cascade_\
        );

    \I__4548\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23672\
        );

    \I__4547\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23672\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__23672\,
            I => \POWERLED.func_state_1_m2_0_0_0\
        );

    \I__4545\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__23666\,
            I => \POWERLED.g1_0_0\
        );

    \I__4543\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__23660\,
            I => \POWERLED.func_state_1_m2_N_3_7_1\
        );

    \I__4541\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23649\
        );

    \I__4540\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23649\
        );

    \I__4539\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23644\
        );

    \I__4538\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23644\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__23649\,
            I => \clk_100Khz_signalkeep_3_fast\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__23644\,
            I => \clk_100Khz_signalkeep_3_fast\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__4534\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__23633\,
            I => \POWERLED.N_671_0\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__23630\,
            I => \G_7_i_a4_1_0_cascade_\
        );

    \I__4531\ : InMux
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__23624\,
            I => \RSMRST_PWRGD.G_7_i_0\
        );

    \I__4529\ : CascadeMux
    port map (
            O => \N__23621\,
            I => \POWERLED.N_533_cascade_\
        );

    \I__4528\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__23615\,
            I => \POWERLED.N_533\
        );

    \I__4526\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__23609\,
            I => \POWERLED.un1_clk_100khz_51_and_i_3_0_sx\
        );

    \I__4524\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23599\
        );

    \I__4522\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23596\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__23599\,
            I => \N__23593\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__23596\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__23593\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__4518\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23584\
        );

    \I__4517\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23581\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__23584\,
            I => \N__23576\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__23581\,
            I => \N__23576\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__23573\,
            I => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\
        );

    \I__4512\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__23567\,
            I => \POWERLED.count_off_0_4\
        );

    \I__4510\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23558\
        );

    \I__4509\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23558\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23555\
        );

    \I__4507\ : Odrv4
    port map (
            O => \N__23555\,
            I => \POWERLED.count_off_RNIZ0Z_1\
        );

    \I__4506\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__23549\,
            I => \POWERLED.count_off_0_1\
        );

    \I__4504\ : CEMux
    port map (
            O => \N__23546\,
            I => \N__23534\
        );

    \I__4503\ : CEMux
    port map (
            O => \N__23545\,
            I => \N__23531\
        );

    \I__4502\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23522\
        );

    \I__4501\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23522\
        );

    \I__4500\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23522\
        );

    \I__4499\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23522\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__23540\,
            I => \N__23515\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__23539\,
            I => \N__23512\
        );

    \I__4496\ : CEMux
    port map (
            O => \N__23538\,
            I => \N__23508\
        );

    \I__4495\ : CEMux
    port map (
            O => \N__23537\,
            I => \N__23505\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23502\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23499\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__23522\,
            I => \N__23496\
        );

    \I__4491\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23491\
        );

    \I__4490\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23491\
        );

    \I__4489\ : CEMux
    port map (
            O => \N__23519\,
            I => \N__23480\
        );

    \I__4488\ : CEMux
    port map (
            O => \N__23518\,
            I => \N__23477\
        );

    \I__4487\ : InMux
    port map (
            O => \N__23515\,
            I => \N__23474\
        );

    \I__4486\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23469\
        );

    \I__4485\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23469\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__23508\,
            I => \N__23466\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__23505\,
            I => \N__23461\
        );

    \I__4482\ : Span4Mux_s2_v
    port map (
            O => \N__23502\,
            I => \N__23461\
        );

    \I__4481\ : Span4Mux_s2_v
    port map (
            O => \N__23499\,
            I => \N__23456\
        );

    \I__4480\ : Span4Mux_s2_v
    port map (
            O => \N__23496\,
            I => \N__23456\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23453\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23442\
        );

    \I__4477\ : CEMux
    port map (
            O => \N__23489\,
            I => \N__23442\
        );

    \I__4476\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23442\
        );

    \I__4475\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23442\
        );

    \I__4474\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23442\
        );

    \I__4473\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23435\
        );

    \I__4472\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23435\
        );

    \I__4471\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23435\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__23480\,
            I => \N__23432\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__23477\,
            I => \N__23429\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__23474\,
            I => \N__23424\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__23469\,
            I => \N__23424\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__23466\,
            I => \N__23415\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__23461\,
            I => \N__23415\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__23456\,
            I => \N__23415\
        );

    \I__4463\ : Span4Mux_v
    port map (
            O => \N__23453\,
            I => \N__23415\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__23442\,
            I => \N__23410\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__23435\,
            I => \N__23410\
        );

    \I__4460\ : Span4Mux_s3_h
    port map (
            O => \N__23432\,
            I => \N__23403\
        );

    \I__4459\ : Span4Mux_s3_v
    port map (
            O => \N__23429\,
            I => \N__23403\
        );

    \I__4458\ : Span4Mux_s3_h
    port map (
            O => \N__23424\,
            I => \N__23403\
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__23415\,
            I => \POWERLED.func_state_RNI7LSV8Z0Z_0\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__23410\,
            I => \POWERLED.func_state_RNI7LSV8Z0Z_0\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__23403\,
            I => \POWERLED.func_state_RNI7LSV8Z0Z_0\
        );

    \I__4454\ : InMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23388\
        );

    \I__4452\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23383\
        );

    \I__4451\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23383\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__23388\,
            I => \N__23380\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23377\
        );

    \I__4448\ : Odrv4
    port map (
            O => \N__23380\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__23377\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__23372\,
            I => \N_7_cascade_\
        );

    \I__4445\ : CascadeMux
    port map (
            O => \N__23369\,
            I => \N_8_0_cascade_\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__23366\,
            I => \POWERLED.g0_5Z0Z_1_cascade_\
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__23363\,
            I => \POWERLED.G_30Z0Z_0_cascade_\
        );

    \I__4442\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23356\
        );

    \I__4441\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23353\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__23356\,
            I => \VPP_VDDQ_un6_count\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__23353\,
            I => \VPP_VDDQ_un6_count\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__23348\,
            I => \G_30_cascade_\
        );

    \I__4437\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23335\
        );

    \I__4435\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23326\
        );

    \I__4434\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23326\
        );

    \I__4433\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23326\
        );

    \I__4432\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23326\
        );

    \I__4431\ : Span4Mux_v
    port map (
            O => \N__23335\,
            I => \N__23323\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__23326\,
            I => \N__23320\
        );

    \I__4429\ : Span4Mux_h
    port map (
            O => \N__23323\,
            I => \N__23315\
        );

    \I__4428\ : Span4Mux_s3_h
    port map (
            O => \N__23320\,
            I => \N__23315\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__23315\,
            I => \N_626\
        );

    \I__4426\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23306\
        );

    \I__4425\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23306\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__23303\,
            I => \N__23298\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__23302\,
            I => \N__23293\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__23301\,
            I => \N__23290\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__23298\,
            I => \N__23286\
        );

    \I__4419\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23283\
        );

    \I__4418\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23274\
        );

    \I__4417\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23274\
        );

    \I__4416\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23274\
        );

    \I__4415\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23274\
        );

    \I__4414\ : Odrv4
    port map (
            O => \N__23286\,
            I => \VPP_VDDQ_curr_state_1\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__23283\,
            I => \VPP_VDDQ_curr_state_1\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__23274\,
            I => \VPP_VDDQ_curr_state_1\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__23267\,
            I => \N__23264\
        );

    \I__4410\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__4408\ : Span4Mux_h
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__4407\ : Span4Mux_h
    port map (
            O => \N__23255\,
            I => \N__23248\
        );

    \I__4406\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23239\
        );

    \I__4405\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23239\
        );

    \I__4404\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23239\
        );

    \I__4403\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23239\
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__23248\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__23239\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__4400\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__23231\,
            I => \POWERLED.count_off_0_3\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__23228\,
            I => \N__23225\
        );

    \I__4397\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23219\
        );

    \I__4396\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23219\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__23213\,
            I => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\
        );

    \I__4392\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__4390\ : Span4Mux_s3_v
    port map (
            O => \N__23204\,
            I => \N__23201\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__23201\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__4388\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__23195\,
            I => \N__23192\
        );

    \I__4386\ : Span4Mux_v
    port map (
            O => \N__23192\,
            I => \N__23188\
        );

    \I__4385\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23185\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__23188\,
            I => \N__23182\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23179\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__23182\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__4381\ : Odrv12
    port map (
            O => \N__23179\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__23174\,
            I => \POWERLED.count_offZ0Z_3_cascade_\
        );

    \I__4379\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23164\
        );

    \I__4377\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23161\
        );

    \I__4376\ : Span4Mux_v
    port map (
            O => \N__23164\,
            I => \N__23158\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__23161\,
            I => \N__23155\
        );

    \I__4374\ : Span4Mux_v
    port map (
            O => \N__23158\,
            I => \N__23152\
        );

    \I__4373\ : Span4Mux_v
    port map (
            O => \N__23155\,
            I => \N__23149\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__23152\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__23149\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__4370\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__23141\,
            I => \POWERLED.un34_clk_100khz_10\
        );

    \I__4368\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23135\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__4366\ : Span12Mux_s5_h
    port map (
            O => \N__23132\,
            I => \N__23129\
        );

    \I__4365\ : Odrv12
    port map (
            O => \N__23129\,
            I => \POWERLED.un34_clk_100khz_11\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__23126\,
            I => \POWERLED.un34_clk_100khz_8_cascade_\
        );

    \I__4363\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23120\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__23117\,
            I => \POWERLED.un34_clk_100khz_9\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__23114\,
            I => \POWERLED.dutycycleZ0Z_9_cascade_\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__23111\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__23108\,
            I => \N__23105\
        );

    \I__4357\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23102\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__23102\,
            I => \POWERLED.un1_dutycycle_53_2_1\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \POWERLED.un1_dutycycle_53_2_1_cascade_\
        );

    \I__4354\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23090\
        );

    \I__4353\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23090\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__23090\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_13\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__23087\,
            I => \VPP_VDDQ.un6_count_8_cascade_\
        );

    \I__4350\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23081\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__23081\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__4348\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23075\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__23075\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__4346\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__23069\,
            I => \VPP_VDDQ.un6_count_9\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__23066\,
            I => \POWERLED.dutycycle_RNI_12Z0Z_8_cascade_\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__4342\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23057\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__23057\,
            I => \POWERLED.dutycycle_RNIZ0Z_15\
        );

    \I__4340\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23051\
        );

    \I__4339\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23045\
        );

    \I__4338\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23045\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__23045\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__23042\,
            I => \POWERLED.dutycycleZ0Z_14_cascade_\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__23039\,
            I => \POWERLED.N_2381_i_cascade_\
        );

    \I__4334\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__23033\,
            I => \POWERLED.un2_count_clk_17_0_0_a2_0_5\
        );

    \I__4332\ : InMux
    port map (
            O => \N__23030\,
            I => \N__23027\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__23027\,
            I => \N__23024\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__23024\,
            I => \POWERLED.dutycycle_RNIZ0Z_13\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__23021\,
            I => \N__23017\
        );

    \I__4328\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23012\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23012\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__23012\,
            I => \POWERLED.dutycycleZ1Z_11\
        );

    \I__4325\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23003\
        );

    \I__4324\ : InMux
    port map (
            O => \N__23008\,
            I => \N__23003\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__4322\ : Span4Mux_v
    port map (
            O => \N__23000\,
            I => \N__22997\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__22997\,
            I => \POWERLED.dutycycle_en_7\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_8_cascade_\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__22991\,
            I => \POWERLED.dutycycle_RNIZ0Z_6_cascade_\
        );

    \I__4318\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__22985\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_7\
        );

    \I__4316\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__22979\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_8\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__4313\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__22970\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_5\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__22967\,
            I => \POWERLED.un1_dutycycle_53_31_a4_1_cascade_\
        );

    \I__4310\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__22961\,
            I => \POWERLED.un1_dutycycle_53_31_a5_1\
        );

    \I__4308\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22955\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__22955\,
            I => \POWERLED.un1_dutycycle_53_31_a0_2\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__22952\,
            I => \N__22949\
        );

    \I__4305\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22946\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__22946\,
            I => \POWERLED.dutycycle_RNIZ0Z_12\
        );

    \I__4303\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22937\
        );

    \I__4302\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22937\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__22937\,
            I => \POWERLED.dutycycleZ1Z_14\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__4299\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22925\
        );

    \I__4298\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22925\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22922\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__22922\,
            I => \POWERLED.dutycycle_en_10\
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__4294\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22910\
        );

    \I__4293\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22910\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__22910\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4291\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22904\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__22904\,
            I => \POWERLED.un1_dutycycle_53_41_0\
        );

    \I__4289\ : CascadeMux
    port map (
            O => \N__22901\,
            I => \POWERLED.un1_dutycycle_53_40_0_cascade_\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__4287\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22892\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__22892\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_13\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__22889\,
            I => \N__22885\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__22888\,
            I => \N__22882\
        );

    \I__4283\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22877\
        );

    \I__4282\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22877\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__22877\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__22874\,
            I => \POWERLED.dutycycleZ0Z_4_cascade_\
        );

    \I__4279\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22866\
        );

    \I__4278\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22863\
        );

    \I__4277\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22860\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__22866\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__22863\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__22860\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__4272\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__22847\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__4270\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22841\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__22841\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_0\
        );

    \I__4268\ : CascadeMux
    port map (
            O => \N__22838\,
            I => \POWERLED.dutycycle_RNIZ0Z_3_cascade_\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__4266\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22829\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__22829\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__4263\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__22820\,
            I => \POWERLED.dutycycle_RNIZ0Z_2\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__4260\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22808\
        );

    \I__4259\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22801\
        );

    \I__4258\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22801\
        );

    \I__4257\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22801\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__22808\,
            I => \N__22798\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__22801\,
            I => \N__22795\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__22798\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__4253\ : Odrv12
    port map (
            O => \N__22795\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__22790\,
            I => \N__22786\
        );

    \I__4251\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22780\
        );

    \I__4250\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22780\
        );

    \I__4249\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22777\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22774\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__22777\,
            I => \N__22771\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__22774\,
            I => \N__22768\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__22771\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__22768\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__4242\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__22757\,
            I => \POWERLED.mult1_un47_sum_axb_4\
        );

    \I__4240\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22751\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__22748\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__4237\ : CascadeMux
    port map (
            O => \N__22745\,
            I => \N__22741\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__22744\,
            I => \N__22738\
        );

    \I__4235\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22735\
        );

    \I__4234\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22732\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22729\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__22732\,
            I => \N__22724\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__22729\,
            I => \N__22724\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__22724\,
            I => \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__4228\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__22715\,
            I => \POWERLED.un1_dutycycle_53_i_29\
        );

    \I__4226\ : InMux
    port map (
            O => \N__22712\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__4224\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__22703\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__4222\ : InMux
    port map (
            O => \N__22700\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__4220\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22691\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__22691\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__4217\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22682\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__22682\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__4215\ : InMux
    port map (
            O => \N__22679\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__4213\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22670\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__22670\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_5\
        );

    \I__4211\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22660\
        );

    \I__4210\ : InMux
    port map (
            O => \N__22666\,
            I => \N__22660\
        );

    \I__4209\ : InMux
    port map (
            O => \N__22665\,
            I => \N__22657\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__22660\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__22657\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__4206\ : InMux
    port map (
            O => \N__22652\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__4204\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__22643\,
            I => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__4202\ : InMux
    port map (
            O => \N__22640\,
            I => \POWERLED.mult1_un47_sum_cry_6\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__22637\,
            I => \N__22633\
        );

    \I__4200\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22627\
        );

    \I__4199\ : InMux
    port map (
            O => \N__22633\,
            I => \N__22627\
        );

    \I__4198\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22624\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__22627\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__22624\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \POWERLED.mult1_un54_sum_s_8_cascade_\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__22616\,
            I => \N__22612\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__22615\,
            I => \N__22608\
        );

    \I__4192\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22601\
        );

    \I__4191\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22601\
        );

    \I__4190\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22601\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__22601\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__22598\,
            I => \POWERLED.N_71_cascade_\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__22595\,
            I => \POWERLED.dutycycleZ0Z_0_cascade_\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__4185\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__4183\ : Span4Mux_h
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__22580\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__22577\,
            I => \POWERLED.N_426_i_cascade_\
        );

    \I__4180\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__22571\,
            I => \POWERLED.dutycycle_eena_1\
        );

    \I__4178\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__22565\,
            I => \POWERLED.N_71\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__22562\,
            I => \POWERLED.dutycycle_eena_1_cascade_\
        );

    \I__4175\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22553\
        );

    \I__4174\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22553\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__22553\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__22550\,
            I => \N__22544\
        );

    \I__4171\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22540\
        );

    \I__4170\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22528\
        );

    \I__4169\ : InMux
    port map (
            O => \N__22547\,
            I => \N__22528\
        );

    \I__4168\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22528\
        );

    \I__4167\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22528\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__22540\,
            I => \N__22525\
        );

    \I__4165\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22514\
        );

    \I__4164\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22514\
        );

    \I__4163\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22514\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__22528\,
            I => \N__22511\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__22525\,
            I => \N__22508\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__22524\,
            I => \N__22505\
        );

    \I__4159\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22500\
        );

    \I__4158\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22497\
        );

    \I__4157\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22494\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__22514\,
            I => \N__22491\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__22511\,
            I => \N__22486\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__22508\,
            I => \N__22486\
        );

    \I__4153\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22481\
        );

    \I__4152\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22481\
        );

    \I__4151\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22478\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__22500\,
            I => \N__22475\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__22497\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__22494\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4147\ : Odrv12
    port map (
            O => \N__22491\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__22486\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__22481\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__22478\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4143\ : Odrv12
    port map (
            O => \N__22475\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4142\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22457\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__22457\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0\
        );

    \I__4140\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22448\
        );

    \I__4139\ : InMux
    port map (
            O => \N__22453\,
            I => \N__22448\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__22448\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__22445\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0_cascade_\
        );

    \I__4136\ : InMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__22439\,
            I => \POWERLED.N_540_1\
        );

    \I__4134\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22433\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__22433\,
            I => \POWERLED.N_542\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22427\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__22427\,
            I => \N__22423\
        );

    \I__4130\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22420\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__22423\,
            I => \POWERLED.N_673\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__22420\,
            I => \POWERLED.N_673\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__22415\,
            I => \POWERLED.func_state_1_m2s2_i_0_1_cascade_\
        );

    \I__4126\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__22409\,
            I => \POWERLED.N_6_1\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__22406\,
            I => \POWERLED.N_74_cascade_\
        );

    \I__4123\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__22400\,
            I => \POWERLED.func_state_1_m2_ns_1_1\
        );

    \I__4121\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22391\
        );

    \I__4120\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22391\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__22391\,
            I => \POWERLED.func_state_1_m2_1\
        );

    \I__4118\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22384\
        );

    \I__4117\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22381\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__22384\,
            I => \N__22378\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__22381\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_0\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__22378\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_0\
        );

    \I__4113\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__22370\,
            I => \POWERLED.N_6_2\
        );

    \I__4111\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__22364\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_a2_0_1_2\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__22361\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_0_2_cascade_\
        );

    \I__4108\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__22355\,
            I => \POWERLED.un1_func_state25_6_0_0_0_2\
        );

    \I__4106\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22346\
        );

    \I__4105\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22346\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__4103\ : Span4Mux_s2_v
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__4102\ : Span4Mux_v
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__22337\,
            I => \POWERLED.func_state_RNI5SKJ1Z0Z_1\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__22334\,
            I => \N__22327\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__22333\,
            I => \N__22324\
        );

    \I__4098\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22319\
        );

    \I__4097\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22312\
        );

    \I__4096\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22312\
        );

    \I__4095\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22312\
        );

    \I__4094\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22305\
        );

    \I__4093\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22305\
        );

    \I__4092\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22305\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22302\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__22312\,
            I => \N__22297\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__22305\,
            I => \N__22297\
        );

    \I__4088\ : Span4Mux_v
    port map (
            O => \N__22302\,
            I => \N__22294\
        );

    \I__4087\ : Span12Mux_v
    port map (
            O => \N__22297\,
            I => \N__22291\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__4085\ : Odrv12
    port map (
            O => \N__22291\,
            I => vddq_ok
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__22288\,
            I => vddq_ok
        );

    \I__4083\ : CascadeMux
    port map (
            O => \N__22283\,
            I => \func_state_RNI_2_0_cascade_\
        );

    \I__4082\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__22277\,
            I => \POWERLED.func_state_1_m0_1_1\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__22274\,
            I => \v5s_enn_cascade_\
        );

    \I__4079\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__22268\,
            I => \POWERLED.func_state_en_0_0\
        );

    \I__4077\ : InMux
    port map (
            O => \N__22265\,
            I => \N__22259\
        );

    \I__4076\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22259\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__22259\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__22256\,
            I => \POWERLED.func_state_en_0_0_cascade_\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__22253\,
            I => \N__22248\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__22252\,
            I => \N__22245\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__22251\,
            I => \N__22242\
        );

    \I__4070\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22237\
        );

    \I__4069\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22237\
        );

    \I__4068\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22234\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__22237\,
            I => \RSMRSTn_fast\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__22234\,
            I => \RSMRSTn_fast\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__22229\,
            I => \N__22226\
        );

    \I__4064\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__22217\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__4059\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__22208\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__4056\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__22199\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__4054\ : CascadeMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__4053\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__4051\ : Span4Mux_h
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__22184\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__4048\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__4046\ : Span4Mux_h
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__22169\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__4044\ : InMux
    port map (
            O => \N__22166\,
            I => \bfn_8_5_0_\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__22163\,
            I => \POWERLED.N_673_0_cascade_\
        );

    \I__4042\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__22157\,
            I => \POWERLED.N_423_0\
        );

    \I__4040\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22148\
        );

    \I__4039\ : InMux
    port map (
            O => \N__22153\,
            I => \N__22148\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__22148\,
            I => \POWERLED.count_off_1_14\
        );

    \I__4037\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__22142\,
            I => \POWERLED.count_off_0_14\
        );

    \I__4035\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22133\
        );

    \I__4034\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22133\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__22133\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNIPGZ0Z497\
        );

    \I__4032\ : InMux
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__22127\,
            I => \POWERLED.count_off_0_15\
        );

    \I__4030\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__22121\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__4028\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22114\
        );

    \I__4027\ : InMux
    port map (
            O => \N__22117\,
            I => \N__22111\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__22114\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__22111\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__4024\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22102\
        );

    \I__4023\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22099\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__22102\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__22099\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__22094\,
            I => \POWERLED.count_offZ0Z_15_cascade_\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__22091\,
            I => \N__22086\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__22090\,
            I => \N__22082\
        );

    \I__4017\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22079\
        );

    \I__4016\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22074\
        );

    \I__4015\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22074\
        );

    \I__4014\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22071\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__22079\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__22074\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__22071\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__4010\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__22055\,
            I => \POWERLED.count_off_0_6\
        );

    \I__4006\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__22049\,
            I => \N__22045\
        );

    \I__4004\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22042\
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__22045\,
            I => \POWERLED.count_off_1_6\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__22042\,
            I => \POWERLED.count_off_1_6\
        );

    \I__4001\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22033\
        );

    \I__4000\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22030\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__22033\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__22030\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__3996\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22019\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22016\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__22016\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__22013\,
            I => \N__22010\
        );

    \I__3992\ : InMux
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__3990\ : Odrv12
    port map (
            O => \N__22004\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__3988\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__3986\ : Odrv4
    port map (
            O => \N__21992\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__3985\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21983\
        );

    \I__3983\ : Span4Mux_h
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__21980\,
            I => \POWERLED.count_off_0_5\
        );

    \I__3981\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__3979\ : Span4Mux_s0_v
    port map (
            O => \N__21971\,
            I => \N__21967\
        );

    \I__3978\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21964\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__21967\,
            I => \POWERLED.count_off_1_5\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__21964\,
            I => \POWERLED.count_off_1_5\
        );

    \I__3975\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__21956\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__21953\,
            I => \POWERLED.count_offZ0Z_5_cascade_\
        );

    \I__3972\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__21947\,
            I => \POWERLED.count_off_0_0\
        );

    \I__3970\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__21941\,
            I => \POWERLED.count_off_1_0\
        );

    \I__3968\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__21935\,
            I => \POWERLED.count_off_0_2\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__3965\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21923\
        );

    \I__3964\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21923\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__21923\,
            I => \POWERLED.count_off_1_2\
        );

    \I__3962\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21916\
        );

    \I__3961\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__21916\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__21913\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__3958\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21902\
        );

    \I__3957\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21902\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__21902\,
            I => \POWERLED.count_off_1_13\
        );

    \I__3955\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__21896\,
            I => \POWERLED.count_off_0_13\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__21893\,
            I => \POWERLED.N_598_cascade_\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__21890\,
            I => \POWERLED.N_450_cascade_\
        );

    \I__3951\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__21884\,
            I => \POWERLED.N_599\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__21881\,
            I => \POWERLED.N_449_cascade_\
        );

    \I__3948\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__21875\,
            I => \POWERLED.N_2376_i\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__21872\,
            I => \POWERLED.N_2376_i_cascade_\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__21869\,
            I => \POWERLED.count_offZ0Z_0_cascade_\
        );

    \I__3944\ : InMux
    port map (
            O => \N__21866\,
            I => \POWERLED.un1_dutycycle_53_cry_14\
        );

    \I__3943\ : InMux
    port map (
            O => \N__21863\,
            I => \bfn_7_15_0_\
        );

    \I__3942\ : InMux
    port map (
            O => \N__21860\,
            I => \POWERLED.CO2\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__3940\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21848\
        );

    \I__3939\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21848\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__21842\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__3934\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__21833\,
            I => \POWERLED.dutycycle_RNIZ0Z_14\
        );

    \I__3932\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21826\
        );

    \I__3931\ : InMux
    port map (
            O => \N__21829\,
            I => \N__21823\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__21826\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__21823\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__3928\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__21815\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__3926\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__21809\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_15\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21799\
        );

    \I__3922\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21796\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__21799\,
            I => \N__21793\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__21796\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__21793\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__3918\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__21782\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__3915\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21775\
        );

    \I__3914\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21772\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21769\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__21772\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__21769\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__3910\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__21761\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__3908\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21754\
        );

    \I__3907\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21751\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__21754\,
            I => \N__21748\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__21751\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__21748\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__3903\ : InMux
    port map (
            O => \N__21743\,
            I => \POWERLED.un1_dutycycle_53_cry_5\
        );

    \I__3902\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21736\
        );

    \I__3901\ : InMux
    port map (
            O => \N__21739\,
            I => \N__21733\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__21736\,
            I => \N__21730\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__21733\,
            I => \N__21727\
        );

    \I__3898\ : Span4Mux_h
    port map (
            O => \N__21730\,
            I => \N__21724\
        );

    \I__3897\ : Odrv12
    port map (
            O => \N__21727\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__21724\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__3895\ : InMux
    port map (
            O => \N__21719\,
            I => \POWERLED.un1_dutycycle_53_cry_6\
        );

    \I__3894\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21712\
        );

    \I__3893\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21709\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21704\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__21709\,
            I => \N__21704\
        );

    \I__3890\ : Span4Mux_s2_v
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__21701\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__3888\ : InMux
    port map (
            O => \N__21698\,
            I => \bfn_7_14_0_\
        );

    \I__3887\ : InMux
    port map (
            O => \N__21695\,
            I => \POWERLED.un1_dutycycle_53_cry_8\
        );

    \I__3886\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21689\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__21689\,
            I => \N__21685\
        );

    \I__3884\ : InMux
    port map (
            O => \N__21688\,
            I => \N__21682\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__21685\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__21682\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__3881\ : InMux
    port map (
            O => \N__21677\,
            I => \POWERLED.un1_dutycycle_53_cry_9\
        );

    \I__3880\ : InMux
    port map (
            O => \N__21674\,
            I => \POWERLED.un1_dutycycle_53_cry_10\
        );

    \I__3879\ : InMux
    port map (
            O => \N__21671\,
            I => \POWERLED.un1_dutycycle_53_cry_11\
        );

    \I__3878\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__3876\ : Span4Mux_v
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__21659\,
            I => \N__21655\
        );

    \I__3874\ : InMux
    port map (
            O => \N__21658\,
            I => \N__21652\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__21655\,
            I => \N__21647\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__21652\,
            I => \N__21647\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__21647\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__3870\ : InMux
    port map (
            O => \N__21644\,
            I => \POWERLED.un1_dutycycle_53_cry_12\
        );

    \I__3869\ : InMux
    port map (
            O => \N__21641\,
            I => \POWERLED.un1_dutycycle_53_cry_13\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__3867\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__21632\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__3865\ : InMux
    port map (
            O => \N__21629\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__21626\,
            I => \N__21622\
        );

    \I__3863\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21617\
        );

    \I__3862\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21617\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__21617\,
            I => \N__21611\
        );

    \I__3860\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21608\
        );

    \I__3859\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21603\
        );

    \I__3858\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21603\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__21611\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__21608\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__21603\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__21596\,
            I => \N__21593\
        );

    \I__3853\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__21590\,
            I => \POWERLED.un1_dutycycle_53_i_28\
        );

    \I__3851\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__3849\ : Span4Mux_v
    port map (
            O => \N__21581\,
            I => \N__21577\
        );

    \I__3848\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21574\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__21577\,
            I => \POWERLED.un1_dutycycle_53_axb_0\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__21574\,
            I => \POWERLED.un1_dutycycle_53_axb_0\
        );

    \I__3845\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21566\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__21566\,
            I => \N__21562\
        );

    \I__3843\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21559\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__21562\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__21559\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__3840\ : InMux
    port map (
            O => \N__21554\,
            I => \POWERLED.un1_dutycycle_53_cry_0\
        );

    \I__3839\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__21548\,
            I => \N__21545\
        );

    \I__3837\ : Span4Mux_v
    port map (
            O => \N__21545\,
            I => \N__21541\
        );

    \I__3836\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21538\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__21541\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__21538\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__3833\ : InMux
    port map (
            O => \N__21533\,
            I => \POWERLED.un1_dutycycle_53_cry_1\
        );

    \I__3832\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__3830\ : Span4Mux_v
    port map (
            O => \N__21524\,
            I => \N__21520\
        );

    \I__3829\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__21520\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__21517\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__3826\ : InMux
    port map (
            O => \N__21512\,
            I => \POWERLED.un1_dutycycle_53_cry_2\
        );

    \I__3825\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21506\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21503\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__21503\,
            I => \N__21499\
        );

    \I__3822\ : InMux
    port map (
            O => \N__21502\,
            I => \N__21496\
        );

    \I__3821\ : Span4Mux_v
    port map (
            O => \N__21499\,
            I => \N__21491\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21491\
        );

    \I__3819\ : Span4Mux_v
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__21488\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__3817\ : InMux
    port map (
            O => \N__21485\,
            I => \POWERLED.un1_dutycycle_53_cry_3\
        );

    \I__3816\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21475\
        );

    \I__3814\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21472\
        );

    \I__3813\ : Span4Mux_h
    port map (
            O => \N__21475\,
            I => \N__21469\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__21472\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__21469\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__3810\ : InMux
    port map (
            O => \N__21464\,
            I => \POWERLED.un1_dutycycle_53_cry_4\
        );

    \I__3809\ : InMux
    port map (
            O => \N__21461\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__3808\ : InMux
    port map (
            O => \N__21458\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__21455\,
            I => \N__21452\
        );

    \I__3806\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21449\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__21449\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__3804\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21443\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21440\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__3801\ : Span4Mux_v
    port map (
            O => \N__21437\,
            I => \N__21434\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__21434\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__21431\,
            I => \N__21428\
        );

    \I__3798\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__21422\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__3795\ : InMux
    port map (
            O => \N__21419\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__3793\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__21410\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__3791\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21404\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__21401\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__3788\ : InMux
    port map (
            O => \N__21398\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__3787\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__21392\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__21389\,
            I => \N__21386\
        );

    \I__3784\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21383\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__21380\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__3781\ : InMux
    port map (
            O => \N__21377\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__3779\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__21368\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__3777\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__3775\ : Span4Mux_h
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__21356\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__3773\ : InMux
    port map (
            O => \N__21353\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__3772\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21347\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__21347\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__3770\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__3768\ : Odrv4
    port map (
            O => \N__21338\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__3767\ : InMux
    port map (
            O => \N__21335\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__3766\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21326\
        );

    \I__3765\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21326\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__21326\,
            I => \N__21323\
        );

    \I__3763\ : Odrv12
    port map (
            O => \N__21323\,
            I => \POWERLED.count_off_1_8\
        );

    \I__3762\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21317\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__21317\,
            I => \POWERLED.count_off_0_8\
        );

    \I__3760\ : InMux
    port map (
            O => \N__21314\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__3759\ : InMux
    port map (
            O => \N__21311\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__3758\ : InMux
    port map (
            O => \N__21308\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__3757\ : InMux
    port map (
            O => \N__21305\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__21302\,
            I => \POWERLED.N_512_cascade_\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__21299\,
            I => \POWERLED.un1_clk_100khz_39_and_i_1_cascade_\
        );

    \I__3754\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21293\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__21293\,
            I => \POWERLED.N_514\
        );

    \I__3752\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21287\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__21287\,
            I => \POWERLED.N_508\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__21284\,
            I => \POWERLED.un1_clk_100khz_33_and_i_1_cascade_\
        );

    \I__3749\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21275\
        );

    \I__3748\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21275\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__3746\ : Span4Mux_v
    port map (
            O => \N__21272\,
            I => \N__21269\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__21269\,
            I => \POWERLED.count_off_1_7\
        );

    \I__3744\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__21263\,
            I => \POWERLED.count_off_0_7\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__21260\,
            I => \POWERLED.func_state_1_ss0_i_0_0_1_1_cascade_\
        );

    \I__3741\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__21254\,
            I => \POWERLED.N_423\
        );

    \I__3739\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__21248\,
            I => \POWERLED.N_671\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__21245\,
            I => \N__21242\
        );

    \I__3736\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21236\
        );

    \I__3735\ : InMux
    port map (
            O => \N__21241\,
            I => \N__21236\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__3733\ : Odrv12
    port map (
            O => \N__21233\,
            I => \POWERLED.func_state_enZ0\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__21230\,
            I => \N__21226\
        );

    \I__3731\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21221\
        );

    \I__3730\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21221\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__21221\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3728\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21208\
        );

    \I__3727\ : InMux
    port map (
            O => \N__21217\,
            I => \N__21208\
        );

    \I__3726\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21199\
        );

    \I__3725\ : InMux
    port map (
            O => \N__21215\,
            I => \N__21199\
        );

    \I__3724\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21199\
        );

    \I__3723\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21199\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__21208\,
            I => \N__21190\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21190\
        );

    \I__3720\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21183\
        );

    \I__3719\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21183\
        );

    \I__3718\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21183\
        );

    \I__3717\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21180\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__21190\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__21183\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__21180\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__3713\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__21170\,
            I => \N__21164\
        );

    \I__3711\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21161\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21156\
        );

    \I__3709\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21156\
        );

    \I__3708\ : Span4Mux_s1_v
    port map (
            O => \N__21164\,
            I => \N__21153\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__21161\,
            I => \N__21145\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__21156\,
            I => \N__21140\
        );

    \I__3705\ : Span4Mux_v
    port map (
            O => \N__21153\,
            I => \N__21140\
        );

    \I__3704\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21129\
        );

    \I__3703\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21129\
        );

    \I__3702\ : InMux
    port map (
            O => \N__21150\,
            I => \N__21129\
        );

    \I__3701\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21129\
        );

    \I__3700\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21129\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__21145\,
            I => \N__21124\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__21140\,
            I => \N__21124\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__21129\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__21124\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__21119\,
            I => \VCCST_EN_i_1_cascade_\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__21116\,
            I => \POWERLED.un1_func_state25_6_0_o_N_5_cascade_\
        );

    \I__3693\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__21110\,
            I => \POWERLED.N_432\
        );

    \I__3691\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__21104\,
            I => \POWERLED.un1_func_state25_6_0_o_N_7_2\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21101\,
            I => \POWERLED.un3_count_off_1_cry_14\
        );

    \I__3688\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21094\
        );

    \I__3687\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21091\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__21088\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__21091\,
            I => \POWERLED.count_off_1_12\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__21088\,
            I => \POWERLED.count_off_1_12\
        );

    \I__3683\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__21077\,
            I => \POWERLED.count_off_0_12\
        );

    \I__3680\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21070\
        );

    \I__3679\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21067\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__21070\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__21067\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3676\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21058\
        );

    \I__3675\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21055\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__21058\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__21055\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__21050\,
            I => \N__21046\
        );

    \I__3671\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21043\
        );

    \I__3670\ : InMux
    port map (
            O => \N__21046\,
            I => \N__21040\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__21043\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__21040\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21031\
        );

    \I__3666\ : InMux
    port map (
            O => \N__21034\,
            I => \N__21028\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__21031\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__21028\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3663\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21019\
        );

    \I__3662\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21016\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__21019\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__21016\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3659\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21007\
        );

    \I__3658\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21004\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__21007\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__21004\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__20999\,
            I => \N__20995\
        );

    \I__3654\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20992\
        );

    \I__3653\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20989\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__20992\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__20989\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3650\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20980\
        );

    \I__3649\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20977\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__20980\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__20977\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__3645\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__20966\,
            I => \N__20963\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__20963\,
            I => \N_555\
        );

    \I__3642\ : SRMux
    port map (
            O => \N__20960\,
            I => \N__20956\
        );

    \I__3641\ : SRMux
    port map (
            O => \N__20959\,
            I => \N__20952\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20949\
        );

    \I__3639\ : SRMux
    port map (
            O => \N__20955\,
            I => \N__20946\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20942\
        );

    \I__3637\ : Span4Mux_s1_v
    port map (
            O => \N__20949\,
            I => \N__20937\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20937\
        );

    \I__3635\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20934\
        );

    \I__3634\ : Span4Mux_v
    port map (
            O => \N__20942\,
            I => \N__20931\
        );

    \I__3633\ : Span4Mux_h
    port map (
            O => \N__20937\,
            I => \N__20926\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__20934\,
            I => \N__20926\
        );

    \I__3631\ : Span4Mux_h
    port map (
            O => \N__20931\,
            I => \N__20921\
        );

    \I__3630\ : Span4Mux_v
    port map (
            O => \N__20926\,
            I => \N__20921\
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__20921\,
            I => \G_14\
        );

    \I__3628\ : InMux
    port map (
            O => \N__20918\,
            I => \N__20914\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__20917\,
            I => \N__20911\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20907\
        );

    \I__3625\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20902\
        );

    \I__3624\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20902\
        );

    \I__3623\ : Span4Mux_h
    port map (
            O => \N__20907\,
            I => \N__20897\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__20902\,
            I => \N__20897\
        );

    \I__3621\ : Sp12to4
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__3620\ : Span12Mux_v
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__3619\ : Odrv12
    port map (
            O => \N__20891\,
            I => \N_662\
        );

    \I__3618\ : InMux
    port map (
            O => \N__20888\,
            I => \POWERLED.un3_count_off_1_cry_6\
        );

    \I__3617\ : InMux
    port map (
            O => \N__20885\,
            I => \POWERLED.un3_count_off_1_cry_7\
        );

    \I__3616\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__20876\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__3613\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20867\
        );

    \I__3612\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20867\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__20864\,
            I => \POWERLED.count_off_1_9\
        );

    \I__3609\ : InMux
    port map (
            O => \N__20861\,
            I => \bfn_7_4_0_\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__3607\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20851\
        );

    \I__3606\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20848\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__20851\,
            I => \N__20845\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__20848\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__20845\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3602\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20834\
        );

    \I__3601\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20834\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__20831\,
            I => \POWERLED.count_off_1_10\
        );

    \I__3598\ : InMux
    port map (
            O => \N__20828\,
            I => \POWERLED.un3_count_off_1_cry_9\
        );

    \I__3597\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20821\
        );

    \I__3596\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20818\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20815\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__20818\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__20815\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3592\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20804\
        );

    \I__3591\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20804\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__20801\,
            I => \POWERLED.count_off_1_11\
        );

    \I__3588\ : InMux
    port map (
            O => \N__20798\,
            I => \POWERLED.un3_count_off_1_cry_10\
        );

    \I__3587\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20791\
        );

    \I__3586\ : InMux
    port map (
            O => \N__20794\,
            I => \N__20788\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__20791\,
            I => \N__20785\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__20788\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__20785\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3582\ : InMux
    port map (
            O => \N__20780\,
            I => \POWERLED.un3_count_off_1_cry_11\
        );

    \I__3581\ : InMux
    port map (
            O => \N__20777\,
            I => \POWERLED.un3_count_off_1_cry_12\
        );

    \I__3580\ : InMux
    port map (
            O => \N__20774\,
            I => \POWERLED.un3_count_off_1_cry_13\
        );

    \I__3579\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__20768\,
            I => \POWERLED.count_off_0_10\
        );

    \I__3577\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__20762\,
            I => \POWERLED.count_off_0_11\
        );

    \I__3575\ : InMux
    port map (
            O => \N__20759\,
            I => \POWERLED.un3_count_off_1_cry_1_cZ0\
        );

    \I__3574\ : InMux
    port map (
            O => \N__20756\,
            I => \POWERLED.un3_count_off_1_cry_2\
        );

    \I__3573\ : InMux
    port map (
            O => \N__20753\,
            I => \POWERLED.un3_count_off_1_cry_3\
        );

    \I__3572\ : InMux
    port map (
            O => \N__20750\,
            I => \POWERLED.un3_count_off_1_cry_4\
        );

    \I__3571\ : InMux
    port map (
            O => \N__20747\,
            I => \POWERLED.un3_count_off_1_cry_5\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__20744\,
            I => \N__20739\
        );

    \I__3569\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20735\
        );

    \I__3568\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20730\
        );

    \I__3567\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20730\
        );

    \I__3566\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20727\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__20735\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__20730\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__20727\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__3561\ : InMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__20714\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__3559\ : InMux
    port map (
            O => \N__20711\,
            I => \N__20708\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__20708\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__3557\ : InMux
    port map (
            O => \N__20705\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__3556\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__20699\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__20696\,
            I => \N__20692\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__20695\,
            I => \N__20688\
        );

    \I__3552\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20681\
        );

    \I__3551\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20681\
        );

    \I__3550\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20681\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__20681\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__3547\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__20672\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__3545\ : InMux
    port map (
            O => \N__20669\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__20666\,
            I => \N__20663\
        );

    \I__3543\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__20660\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__3541\ : InMux
    port map (
            O => \N__20657\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__20654\,
            I => \N__20650\
        );

    \I__3539\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20642\
        );

    \I__3538\ : InMux
    port map (
            O => \N__20650\,
            I => \N__20642\
        );

    \I__3537\ : InMux
    port map (
            O => \N__20649\,
            I => \N__20639\
        );

    \I__3536\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20634\
        );

    \I__3535\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20634\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__20642\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__20639\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__20634\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__3531\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__20624\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__3529\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20618\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__20618\,
            I => \POWERLED.count_off_0_9\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__20615\,
            I => \POWERLED.count_offZ0Z_9_cascade_\
        );

    \I__3526\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__20609\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__3524\ : InMux
    port map (
            O => \N__20606\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__3523\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20600\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__20600\,
            I => \N__20596\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__20599\,
            I => \N__20592\
        );

    \I__3520\ : Span4Mux_s2_v
    port map (
            O => \N__20596\,
            I => \N__20588\
        );

    \I__3519\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20583\
        );

    \I__3518\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20583\
        );

    \I__3517\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20580\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__20588\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__20583\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__20580\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__20573\,
            I => \N__20570\
        );

    \I__3512\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__20567\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__3510\ : InMux
    port map (
            O => \N__20564\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__3509\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__20558\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__20555\,
            I => \N__20551\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__20554\,
            I => \N__20547\
        );

    \I__3505\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20540\
        );

    \I__3504\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20540\
        );

    \I__3503\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20540\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__20540\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__3501\ : InMux
    port map (
            O => \N__20537\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__3499\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__20528\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__3497\ : InMux
    port map (
            O => \N__20525\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__20522\,
            I => \POWERLED.mult1_un75_sum_s_8_cascade_\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__20519\,
            I => \N__20516\
        );

    \I__3494\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__20513\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__3492\ : InMux
    port map (
            O => \N__20510\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__20507\,
            I => \N__20504\
        );

    \I__3490\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20501\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__20501\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__3488\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__20495\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__3486\ : InMux
    port map (
            O => \N__20492\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__3485\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20486\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__20486\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__3482\ : InMux
    port map (
            O => \N__20480\,
            I => \N__20477\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__20477\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__3480\ : InMux
    port map (
            O => \N__20474\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__3479\ : InMux
    port map (
            O => \N__20471\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__3478\ : InMux
    port map (
            O => \N__20468\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__3477\ : InMux
    port map (
            O => \N__20465\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__20462\,
            I => \N__20458\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__20461\,
            I => \N__20454\
        );

    \I__3474\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20447\
        );

    \I__3473\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20447\
        );

    \I__3472\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20447\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__20447\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__3470\ : InMux
    port map (
            O => \N__20444\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__3469\ : InMux
    port map (
            O => \N__20441\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__20438\,
            I => \POWERLED.mult1_un68_sum_s_8_cascade_\
        );

    \I__3467\ : InMux
    port map (
            O => \N__20435\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__3465\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__20426\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__3463\ : InMux
    port map (
            O => \N__20423\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__3462\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__20414\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__3458\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__20402\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__3455\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__3453\ : Span4Mux_h
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__20390\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__3451\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__20381\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__3448\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__20375\,
            I => \N__20372\
        );

    \I__3446\ : Span4Mux_v
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__20369\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__3444\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__3442\ : Span4Mux_s3_v
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__20357\,
            I => \POWERLED.mult1_un61_sum_i_8\
        );

    \I__3440\ : InMux
    port map (
            O => \N__20354\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__3438\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__20345\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__3436\ : InMux
    port map (
            O => \N__20342\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__3435\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__20336\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__20333\,
            I => \N__20330\
        );

    \I__3432\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__20327\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__3430\ : InMux
    port map (
            O => \N__20324\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__3429\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__20318\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__3427\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__20312\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__3425\ : InMux
    port map (
            O => \N__20309\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__3424\ : InMux
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__20303\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__3422\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__20297\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__3420\ : InMux
    port map (
            O => \N__20294\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__3419\ : InMux
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__20288\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__3417\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__20282\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__3415\ : InMux
    port map (
            O => \N__20279\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__3414\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__20273\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__3412\ : InMux
    port map (
            O => \N__20270\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__3411\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20263\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__20266\,
            I => \N__20260\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__20263\,
            I => \N__20254\
        );

    \I__3408\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20247\
        );

    \I__3407\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20247\
        );

    \I__3406\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20247\
        );

    \I__3405\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20244\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__20254\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__20247\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__20244\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__20237\,
            I => \N__20232\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__20236\,
            I => \N__20229\
        );

    \I__3399\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20224\
        );

    \I__3398\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20221\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20216\
        );

    \I__3396\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20216\
        );

    \I__3395\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20213\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__20224\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__20221\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__20216\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__20213\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__20204\,
            I => \N__20200\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__20203\,
            I => \N__20197\
        );

    \I__3388\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20193\
        );

    \I__3387\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20188\
        );

    \I__3386\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20188\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__20193\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__20188\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__3382\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__20174\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__3379\ : InMux
    port map (
            O => \N__20171\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__3378\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__20165\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__3376\ : InMux
    port map (
            O => \N__20162\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__3374\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__20153\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__3372\ : InMux
    port map (
            O => \N__20150\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__3371\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__20144\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__3369\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20137\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__20140\,
            I => \N__20134\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N__20129\
        );

    \I__3366\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20124\
        );

    \I__3365\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20124\
        );

    \I__3364\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20121\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__20129\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__20124\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__20121\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3360\ : InMux
    port map (
            O => \N__20114\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__20111\,
            I => \N__20107\
        );

    \I__3358\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20099\
        );

    \I__3357\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20099\
        );

    \I__3356\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20099\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__20099\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__3353\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__20090\,
            I => \N__20087\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__20087\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__3350\ : InMux
    port map (
            O => \N__20084\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__3349\ : InMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__20078\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__3347\ : InMux
    port map (
            O => \N__20075\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__3346\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20068\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__20071\,
            I => \N__20064\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__20068\,
            I => \N__20059\
        );

    \I__3343\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20056\
        );

    \I__3342\ : InMux
    port map (
            O => \N__20064\,
            I => \N__20051\
        );

    \I__3341\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20051\
        );

    \I__3340\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20048\
        );

    \I__3339\ : Odrv12
    port map (
            O => \N__20059\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__20056\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__20051\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__20048\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__20039\,
            I => \N__20034\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__20038\,
            I => \N__20031\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__20037\,
            I => \N__20028\
        );

    \I__3332\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20025\
        );

    \I__3331\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20020\
        );

    \I__3330\ : InMux
    port map (
            O => \N__20028\,
            I => \N__20020\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__20025\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__20020\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__3327\ : InMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__20012\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__3325\ : InMux
    port map (
            O => \N__20009\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__3324\ : InMux
    port map (
            O => \N__20006\,
            I => \N__20003\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__20003\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__3321\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__19994\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__3319\ : InMux
    port map (
            O => \N__19991\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__3317\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__19982\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__3315\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__19976\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__3313\ : InMux
    port map (
            O => \N__19973\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__3312\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__19967\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__3309\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__19958\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__3307\ : InMux
    port map (
            O => \N__19955\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__3306\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__19949\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__3304\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__19943\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__3302\ : InMux
    port map (
            O => \N__19940\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__3301\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__19934\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__3299\ : InMux
    port map (
            O => \N__19931\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__3298\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__19925\,
            I => \N__19921\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__19924\,
            I => \N__19918\
        );

    \I__3295\ : Span4Mux_v
    port map (
            O => \N__19921\,
            I => \N__19913\
        );

    \I__3294\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19908\
        );

    \I__3293\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19908\
        );

    \I__3292\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19905\
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__19913\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__19908\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__19905\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__19898\,
            I => \POWERLED.mult1_un138_sum_s_8_cascade_\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__19895\,
            I => \N__19891\
        );

    \I__3286\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19883\
        );

    \I__3285\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19883\
        );

    \I__3284\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19883\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__19883\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__3282\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__19877\,
            I => \VPP_VDDQ.un1_count_2_1_axb_6\
        );

    \I__3280\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__19871\,
            I => \VPP_VDDQ.count_2_0_4\
        );

    \I__3278\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19862\
        );

    \I__3277\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19862\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__19862\,
            I => \VPP_VDDQ.count_2_1_4\
        );

    \I__3275\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__19856\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__3273\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19847\
        );

    \I__3272\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19847\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__19847\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__19844\,
            I => \VPP_VDDQ.count_2Z0Z_4_cascade_\
        );

    \I__3269\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19832\
        );

    \I__3268\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19832\
        );

    \I__3267\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19832\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__19832\,
            I => \VPP_VDDQ.count_2_1_6\
        );

    \I__3265\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__19820\,
            I => \VPP_VDDQ.un9_clk_100khz_0\
        );

    \I__3261\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__19814\,
            I => \VPP_VDDQ.count_2_0_2\
        );

    \I__3259\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19805\
        );

    \I__3258\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19805\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__19805\,
            I => \VPP_VDDQ.count_2_1_2\
        );

    \I__3256\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19789\
        );

    \I__3255\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19789\
        );

    \I__3254\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19789\
        );

    \I__3253\ : CEMux
    port map (
            O => \N__19799\,
            I => \N__19789\
        );

    \I__3252\ : CEMux
    port map (
            O => \N__19798\,
            I => \N__19786\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__19789\,
            I => \N__19767\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19767\
        );

    \I__3249\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19754\
        );

    \I__3248\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19754\
        );

    \I__3247\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19754\
        );

    \I__3246\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19754\
        );

    \I__3245\ : CEMux
    port map (
            O => \N__19781\,
            I => \N__19750\
        );

    \I__3244\ : CEMux
    port map (
            O => \N__19780\,
            I => \N__19747\
        );

    \I__3243\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19738\
        );

    \I__3242\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19738\
        );

    \I__3241\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19738\
        );

    \I__3240\ : CEMux
    port map (
            O => \N__19776\,
            I => \N__19738\
        );

    \I__3239\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19729\
        );

    \I__3238\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19729\
        );

    \I__3237\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19729\
        );

    \I__3236\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19729\
        );

    \I__3235\ : Span4Mux_h
    port map (
            O => \N__19767\,
            I => \N__19726\
        );

    \I__3234\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19717\
        );

    \I__3233\ : CEMux
    port map (
            O => \N__19765\,
            I => \N__19717\
        );

    \I__3232\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19717\
        );

    \I__3231\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19717\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__19754\,
            I => \N__19714\
        );

    \I__3229\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19711\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19706\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__19747\,
            I => \N__19706\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__19738\,
            I => \N__19701\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__19729\,
            I => \N__19701\
        );

    \I__3224\ : Span4Mux_s3_h
    port map (
            O => \N__19726\,
            I => \N__19694\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19694\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__19714\,
            I => \N__19694\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__19711\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__19706\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__19701\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__19694\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__3217\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__19682\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__3215\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__19673\,
            I => \N__19669\
        );

    \I__3212\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19666\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__19669\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__19666\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__3209\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19654\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__19657\,
            I => \N__19651\
        );

    \I__3206\ : Span12Mux_s8_h
    port map (
            O => \N__19654\,
            I => \N__19648\
        );

    \I__3205\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19645\
        );

    \I__3204\ : Odrv12
    port map (
            O => \N__19648\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__19645\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__19640\,
            I => \VPP_VDDQ.count_2Z0Z_2_cascade_\
        );

    \I__3201\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__19631\,
            I => \N__19627\
        );

    \I__3198\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19624\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__19627\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__19624\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__3195\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__3193\ : Span4Mux_h
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__19610\,
            I => \VPP_VDDQ.un9_clk_100khz_9\
        );

    \I__3191\ : InMux
    port map (
            O => \N__19607\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__3190\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19600\
        );

    \I__3189\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19597\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__19600\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__19597\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3186\ : InMux
    port map (
            O => \N__19592\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__3185\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19585\
        );

    \I__3184\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19582\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__19585\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__19582\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__3181\ : InMux
    port map (
            O => \N__19577\,
            I => \bfn_6_7_0_\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__19574\,
            I => \N__19570\
        );

    \I__3179\ : InMux
    port map (
            O => \N__19573\,
            I => \N__19567\
        );

    \I__3178\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19564\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__19567\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__19564\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__3175\ : InMux
    port map (
            O => \N__19559\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__3174\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19552\
        );

    \I__3173\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19549\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__19552\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__19549\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__3170\ : InMux
    port map (
            O => \N__19544\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__3168\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19534\
        );

    \I__3167\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19531\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__19534\,
            I => \N__19528\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__19531\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__3164\ : Odrv12
    port map (
            O => \N__19528\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__3163\ : InMux
    port map (
            O => \N__19523\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__3162\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19516\
        );

    \I__3161\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19513\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19510\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__19513\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__3158\ : Odrv12
    port map (
            O => \N__19510\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__3157\ : InMux
    port map (
            O => \N__19505\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__3156\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19498\
        );

    \I__3155\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19495\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__19498\,
            I => \N__19492\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__19495\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__3152\ : Odrv12
    port map (
            O => \N__19492\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__3151\ : InMux
    port map (
            O => \N__19487\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__3150\ : InMux
    port map (
            O => \N__19484\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__3149\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19477\
        );

    \I__3148\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__19474\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__3145\ : Odrv12
    port map (
            O => \N__19471\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__3144\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19462\
        );

    \I__3143\ : InMux
    port map (
            O => \N__19465\,
            I => \N__19459\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__19462\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__19459\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3140\ : InMux
    port map (
            O => \N__19454\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__3139\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19447\
        );

    \I__3138\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19444\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__19447\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__19444\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3135\ : InMux
    port map (
            O => \N__19439\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__3134\ : InMux
    port map (
            O => \N__19436\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__3133\ : InMux
    port map (
            O => \N__19433\,
            I => \bfn_6_6_0_\
        );

    \I__3132\ : InMux
    port map (
            O => \N__19430\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__3131\ : InMux
    port map (
            O => \N__19427\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__3130\ : InMux
    port map (
            O => \N__19424\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__3129\ : InMux
    port map (
            O => \N__19421\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__3128\ : InMux
    port map (
            O => \N__19418\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__19415\,
            I => \N__19411\
        );

    \I__3126\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19407\
        );

    \I__3125\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19404\
        );

    \I__3124\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19401\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__19407\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__19404\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__19401\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3120\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__19391\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__3118\ : InMux
    port map (
            O => \N__19388\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__3117\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19381\
        );

    \I__3116\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19378\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__19381\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__19378\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3113\ : InMux
    port map (
            O => \N__19373\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__3112\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19366\
        );

    \I__3111\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__19366\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__19363\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3108\ : InMux
    port map (
            O => \N__19358\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__3107\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19351\
        );

    \I__3106\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19348\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__19351\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__19348\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3103\ : InMux
    port map (
            O => \N__19343\,
            I => \bfn_6_5_0_\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__19340\,
            I => \N__19336\
        );

    \I__3101\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19333\
        );

    \I__3100\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19330\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__19333\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__19330\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3097\ : InMux
    port map (
            O => \N__19325\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__3096\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19318\
        );

    \I__3095\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19315\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__19318\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__19315\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3092\ : InMux
    port map (
            O => \N__19310\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__19307\,
            I => \N__19303\
        );

    \I__3090\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19300\
        );

    \I__3089\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19297\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__19300\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__19297\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3086\ : InMux
    port map (
            O => \N__19292\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__3085\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19285\
        );

    \I__3084\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19282\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19285\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__19282\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3081\ : InMux
    port map (
            O => \N__19277\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__3080\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19270\
        );

    \I__3079\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19267\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__19270\,
            I => \N__19264\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__19267\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__3076\ : Odrv4
    port map (
            O => \N__19264\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__3075\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19255\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__19258\,
            I => \N__19251\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__19255\,
            I => \N__19248\
        );

    \I__3072\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19243\
        );

    \I__3071\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19243\
        );

    \I__3070\ : Span4Mux_s0_v
    port map (
            O => \N__19248\,
            I => \N__19240\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__19243\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__19240\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19231\
        );

    \I__3066\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19228\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__19231\,
            I => \N__19225\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__19228\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__19225\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__3062\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__19217\,
            I => \HDA_STRAP.un4_count_9\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19202\
        );

    \I__3059\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19202\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__19212\,
            I => \N__19199\
        );

    \I__3057\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19186\
        );

    \I__3056\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19186\
        );

    \I__3055\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19186\
        );

    \I__3054\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19186\
        );

    \I__3053\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19186\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19183\
        );

    \I__3051\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19180\
        );

    \I__3050\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19175\
        );

    \I__3049\ : InMux
    port map (
            O => \N__19197\,
            I => \N__19175\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__19186\,
            I => \N__19170\
        );

    \I__3047\ : Span4Mux_v
    port map (
            O => \N__19183\,
            I => \N__19170\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__19180\,
            I => \HDA_STRAP.un4_count\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__19175\,
            I => \HDA_STRAP.un4_count\
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__19170\,
            I => \HDA_STRAP.un4_count\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__19163\,
            I => \N__19157\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__19162\,
            I => \N__19154\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__19161\,
            I => \N__19151\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__19160\,
            I => \N__19147\
        );

    \I__3039\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19141\
        );

    \I__3038\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19135\
        );

    \I__3037\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19135\
        );

    \I__3036\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19132\
        );

    \I__3035\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19127\
        );

    \I__3034\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19127\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__19145\,
            I => \N__19124\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__19144\,
            I => \N__19121\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__19141\,
            I => \N__19117\
        );

    \I__3030\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19114\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__19135\,
            I => \N__19111\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__19132\,
            I => \N__19106\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19106\
        );

    \I__3026\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19099\
        );

    \I__3025\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19099\
        );

    \I__3024\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19099\
        );

    \I__3023\ : Span4Mux_s1_v
    port map (
            O => \N__19117\,
            I => \N__19096\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__19114\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__3021\ : Odrv12
    port map (
            O => \N__19111\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__3020\ : Odrv12
    port map (
            O => \N__19106\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__19099\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__19096\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__3016\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__19079\,
            I => \HDA_STRAP.un1_count_1_cry_15_THRU_CO\
        );

    \I__3014\ : InMux
    port map (
            O => \N__19076\,
            I => \N__19071\
        );

    \I__3013\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19066\
        );

    \I__3012\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19066\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__19071\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__19066\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__3009\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19055\
        );

    \I__3008\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19052\
        );

    \I__3007\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19047\
        );

    \I__3006\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19047\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__19055\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__19052\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__19047\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__19040\,
            I => \N__19035\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__19039\,
            I => \N__19032\
        );

    \I__3000\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19029\
        );

    \I__2999\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19026\
        );

    \I__2998\ : InMux
    port map (
            O => \N__19032\,
            I => \N__19023\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__19029\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__19026\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__19023\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__19016\,
            I => \N__19011\
        );

    \I__2993\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19008\
        );

    \I__2992\ : InMux
    port map (
            O => \N__19014\,
            I => \N__19003\
        );

    \I__2991\ : InMux
    port map (
            O => \N__19011\,
            I => \N__19003\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__19008\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__19003\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2988\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__2986\ : Odrv12
    port map (
            O => \N__18992\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__2985\ : InMux
    port map (
            O => \N__18989\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__2984\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18981\
        );

    \I__2983\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18978\
        );

    \I__2982\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18975\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__18981\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__18978\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__18975\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2978\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__18965\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__2976\ : InMux
    port map (
            O => \N__18962\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__2975\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18954\
        );

    \I__2974\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18949\
        );

    \I__2973\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18949\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__18954\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__18949\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2970\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__18941\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__2968\ : InMux
    port map (
            O => \N__18938\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__2967\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18930\
        );

    \I__2966\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18925\
        );

    \I__2965\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18925\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__18930\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__18925\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2962\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__18917\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__2960\ : InMux
    port map (
            O => \N__18914\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__2959\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18906\
        );

    \I__2958\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18903\
        );

    \I__2957\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18900\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__18906\,
            I => \N__18895\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__18903\,
            I => \N__18895\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__18900\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__18895\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__2952\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18886\
        );

    \I__2951\ : InMux
    port map (
            O => \N__18889\,
            I => \N__18883\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__18886\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__18883\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__2947\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18870\
        );

    \I__2946\ : InMux
    port map (
            O => \N__18874\,
            I => \N__18867\
        );

    \I__2945\ : InMux
    port map (
            O => \N__18873\,
            I => \N__18864\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__18870\,
            I => \N__18861\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__18867\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__18864\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__2941\ : Odrv12
    port map (
            O => \N__18861\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__2940\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18850\
        );

    \I__2939\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18847\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__18850\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__18847\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__2936\ : InMux
    port map (
            O => \N__18842\,
            I => \N__18838\
        );

    \I__2935\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__18838\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__18835\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__2932\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18826\
        );

    \I__2931\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18823\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__18826\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__18823\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__2927\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18811\
        );

    \I__2926\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18808\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__18811\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__18808\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__2923\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18799\
        );

    \I__2922\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18796\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__18799\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__18796\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__2919\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18787\
        );

    \I__2918\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18784\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__18787\,
            I => \N__18778\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__18784\,
            I => \N__18778\
        );

    \I__2915\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18775\
        );

    \I__2914\ : Span4Mux_s1_v
    port map (
            O => \N__18778\,
            I => \N__18772\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__18775\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__18772\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__2911\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18762\
        );

    \I__2910\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18759\
        );

    \I__2909\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18756\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__18762\,
            I => \N__18753\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__18759\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__18756\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__18753\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__2904\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__18743\,
            I => \HDA_STRAP.un4_count_12\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \HDA_STRAP.un4_count_13_cascade_\
        );

    \I__2901\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__18734\,
            I => \HDA_STRAP.un4_count_10\
        );

    \I__2899\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18727\
        );

    \I__2898\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18724\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__18727\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__18724\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__2895\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18715\
        );

    \I__2894\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18712\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__18715\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__18712\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__18707\,
            I => \N__18703\
        );

    \I__2890\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__2889\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18697\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__18700\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__18697\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__2886\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18688\
        );

    \I__2885\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18685\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__18688\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__18685\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__2882\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__18677\,
            I => \HDA_STRAP.un4_count_11\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__2879\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__18668\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__2877\ : InMux
    port map (
            O => \N__18665\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__2876\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__18659\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__2874\ : InMux
    port map (
            O => \N__18656\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__2872\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__18647\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__2870\ : InMux
    port map (
            O => \N__18644\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__2869\ : InMux
    port map (
            O => \N__18641\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__18638\,
            I => \N__18633\
        );

    \I__2867\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18629\
        );

    \I__2866\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18624\
        );

    \I__2865\ : InMux
    port map (
            O => \N__18633\,
            I => \N__18624\
        );

    \I__2864\ : InMux
    port map (
            O => \N__18632\,
            I => \N__18621\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__18629\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__18624\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__18621\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__18614\,
            I => \POWERLED.mult1_un89_sum_s_8_cascade_\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__18611\,
            I => \N__18607\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__18610\,
            I => \N__18603\
        );

    \I__2857\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18596\
        );

    \I__2856\ : InMux
    port map (
            O => \N__18606\,
            I => \N__18596\
        );

    \I__2855\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18596\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__18596\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__2852\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__18587\,
            I => \POWERLED.mult1_un75_sum_i_8\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__18584\,
            I => \N__18580\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__18583\,
            I => \N__18576\
        );

    \I__2848\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18569\
        );

    \I__2847\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18569\
        );

    \I__2846\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18569\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__18569\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__2844\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__18560\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__2841\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__18554\,
            I => \POWERLED.mult1_un82_sum_i_8\
        );

    \I__2839\ : InMux
    port map (
            O => \N__18551\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__2837\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__18542\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__2835\ : InMux
    port map (
            O => \N__18539\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__2834\ : InMux
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__18533\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__2832\ : InMux
    port map (
            O => \N__18530\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__2830\ : InMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__18521\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__2828\ : InMux
    port map (
            O => \N__18518\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__2827\ : InMux
    port map (
            O => \N__18515\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__2826\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18505\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__18508\,
            I => \N__18501\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__18505\,
            I => \N__18496\
        );

    \I__2822\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18491\
        );

    \I__2821\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18491\
        );

    \I__2820\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18488\
        );

    \I__2819\ : InMux
    port map (
            O => \N__18499\,
            I => \N__18485\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__18496\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__18491\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__18488\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__18485\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2814\ : InMux
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__18473\,
            I => \POWERLED.mult1_un131_sum_i_8\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__2811\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__18464\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__2809\ : InMux
    port map (
            O => \N__18461\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__2808\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__18455\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__2806\ : InMux
    port map (
            O => \N__18452\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__2805\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__18446\,
            I => \POWERLED.mult1_un138_sum_i_8\
        );

    \I__2803\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__18440\,
            I => \POWERLED.un85_clk_100khz_1\
        );

    \I__2801\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__18431\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__18428\,
            I => \N__18424\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__18427\,
            I => \N__18420\
        );

    \I__2796\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18413\
        );

    \I__2795\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18413\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18413\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__18413\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__18410\,
            I => \N__18405\
        );

    \I__2791\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18401\
        );

    \I__2790\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18396\
        );

    \I__2789\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18396\
        );

    \I__2788\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18393\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__18401\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__18396\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__18393\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__2783\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__18377\,
            I => \POWERLED.mult1_un103_sum_i_8\
        );

    \I__2780\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18368\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__18373\,
            I => \N__18365\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__18372\,
            I => \N__18362\
        );

    \I__2777\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18358\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__18368\,
            I => \N__18355\
        );

    \I__2775\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18352\
        );

    \I__2774\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18347\
        );

    \I__2773\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18347\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__18358\,
            I => \N__18344\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__18355\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__18352\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__18347\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__18344\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2767\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__18332\,
            I => \POWERLED.mult1_un124_sum_i_8\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__2764\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18323\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__18323\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__2762\ : InMux
    port map (
            O => \N__18320\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__2761\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18314\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__18314\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__18311\,
            I => \N__18307\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__18310\,
            I => \N__18303\
        );

    \I__2757\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18296\
        );

    \I__2756\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18296\
        );

    \I__2755\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18296\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__18296\,
            I => \G_2150\
        );

    \I__2753\ : InMux
    port map (
            O => \N__18293\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__2752\ : InMux
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__18284\,
            I => \POWERLED.un85_clk_100khz_0\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__18275\,
            I => \POWERLED.un85_clk_100khz_2\
        );

    \I__2746\ : InMux
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18269\,
            I => \POWERLED.un85_clk_100khz_3\
        );

    \I__2744\ : InMux
    port map (
            O => \N__18266\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__18263\,
            I => \N__18258\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__18262\,
            I => \N__18255\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__18261\,
            I => \N__18252\
        );

    \I__2740\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18249\
        );

    \I__2739\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18244\
        );

    \I__2738\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18244\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__18249\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__18244\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18239\,
            I => \POWERLED.mult1_un145_sum_cry_2_c\
        );

    \I__2734\ : InMux
    port map (
            O => \N__18236\,
            I => \POWERLED.mult1_un145_sum_cry_3_c\
        );

    \I__2733\ : InMux
    port map (
            O => \N__18233\,
            I => \POWERLED.mult1_un145_sum_cry_4_c\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18230\,
            I => \POWERLED.mult1_un145_sum_cry_5_c\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18227\,
            I => \POWERLED.mult1_un145_sum_cry_6_c\
        );

    \I__2730\ : InMux
    port map (
            O => \N__18224\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__18221\,
            I => \POWERLED.mult1_un145_sum_s_8_cascade_\
        );

    \I__2728\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18214\
        );

    \I__2727\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18211\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18214\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__18211\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__2724\ : InMux
    port map (
            O => \N__18206\,
            I => \N__18186\
        );

    \I__2723\ : InMux
    port map (
            O => \N__18205\,
            I => \N__18186\
        );

    \I__2722\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18186\
        );

    \I__2721\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18179\
        );

    \I__2720\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18179\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18179\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18170\
        );

    \I__2717\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18170\
        );

    \I__2716\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18170\
        );

    \I__2715\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18170\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18161\
        );

    \I__2713\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18161\
        );

    \I__2712\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18161\
        );

    \I__2711\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18161\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__18186\,
            I => \N__18155\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__18179\,
            I => \N__18155\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18150\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__18161\,
            I => \N__18150\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__18160\,
            I => \N__18146\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__18155\,
            I => \N__18142\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__18150\,
            I => \N__18139\
        );

    \I__2703\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18132\
        );

    \I__2702\ : InMux
    port map (
            O => \N__18146\,
            I => \N__18132\
        );

    \I__2701\ : InMux
    port map (
            O => \N__18145\,
            I => \N__18132\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__18142\,
            I => \VPP_VDDQ.count_2_1_sqmuxa\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__18139\,
            I => \VPP_VDDQ.count_2_1_sqmuxa\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__18132\,
            I => \VPP_VDDQ.count_2_1_sqmuxa\
        );

    \I__2697\ : InMux
    port map (
            O => \N__18125\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__2696\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18118\
        );

    \I__2695\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18115\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__18118\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__18115\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\
        );

    \I__2692\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__18107\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__2690\ : InMux
    port map (
            O => \N__18104\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__2689\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__18098\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__2687\ : InMux
    port map (
            O => \N__18095\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__2686\ : InMux
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__18089\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__2684\ : InMux
    port map (
            O => \N__18086\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__2683\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__18080\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__2681\ : InMux
    port map (
            O => \N__18077\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__2680\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__18071\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__2678\ : InMux
    port map (
            O => \N__18068\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__2677\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__18062\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__2675\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__18053\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18044\
        );

    \I__2671\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18044\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__18044\,
            I => \N__18040\
        );

    \I__2669\ : InMux
    port map (
            O => \N__18043\,
            I => \N__18037\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__18040\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__18037\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__2666\ : InMux
    port map (
            O => \N__18032\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__2665\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18025\
        );

    \I__2664\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18022\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__18025\,
            I => \VPP_VDDQ.count_2_1_8\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__18022\,
            I => \VPP_VDDQ.count_2_1_8\
        );

    \I__2661\ : InMux
    port map (
            O => \N__18017\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__2660\ : InMux
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__18008\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__2657\ : InMux
    port map (
            O => \N__18005\,
            I => \N__17999\
        );

    \I__2656\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17999\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__17996\,
            I => \VPP_VDDQ.count_2_1_9\
        );

    \I__2653\ : InMux
    port map (
            O => \N__17993\,
            I => \bfn_5_9_0_\
        );

    \I__2652\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__17987\,
            I => \N__17983\
        );

    \I__2650\ : InMux
    port map (
            O => \N__17986\,
            I => \N__17980\
        );

    \I__2649\ : Odrv4
    port map (
            O => \N__17983\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__17980\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2647\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17971\
        );

    \I__2646\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17968\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__17971\,
            I => \N__17965\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__17968\,
            I => \VPP_VDDQ.count_2_1_10\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__17965\,
            I => \VPP_VDDQ.count_2_1_10\
        );

    \I__2642\ : InMux
    port map (
            O => \N__17960\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__2641\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17953\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__17956\,
            I => \N__17950\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__17953\,
            I => \N__17947\
        );

    \I__2638\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17944\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__17947\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__17944\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__2635\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17933\
        );

    \I__2634\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17933\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__17933\,
            I => \N__17930\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__17930\,
            I => \VPP_VDDQ.count_2_1_11\
        );

    \I__2631\ : InMux
    port map (
            O => \N__17927\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__2630\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17920\
        );

    \I__2629\ : InMux
    port map (
            O => \N__17923\,
            I => \N__17917\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__17920\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__17917\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2626\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17906\
        );

    \I__2625\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17906\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__17906\,
            I => \VPP_VDDQ.count_2_1_12\
        );

    \I__2623\ : InMux
    port map (
            O => \N__17903\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__17900\,
            I => \N__17896\
        );

    \I__2621\ : InMux
    port map (
            O => \N__17899\,
            I => \N__17893\
        );

    \I__2620\ : InMux
    port map (
            O => \N__17896\,
            I => \N__17890\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__17893\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__17890\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__2617\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17879\
        );

    \I__2616\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17879\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__17879\,
            I => \VPP_VDDQ.count_2_1_13\
        );

    \I__2614\ : InMux
    port map (
            O => \N__17876\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__2613\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17869\
        );

    \I__2612\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17866\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__17869\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__17866\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__2609\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17855\
        );

    \I__2608\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17855\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__17855\,
            I => \VPP_VDDQ.count_2_1_14\
        );

    \I__2606\ : InMux
    port map (
            O => \N__17852\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__2605\ : InMux
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__17843\,
            I => \VPP_VDDQ.count_2_0_5\
        );

    \I__2602\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__17834\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__2599\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__17825\,
            I => \VPP_VDDQ.count_2_0_10\
        );

    \I__2596\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17817\
        );

    \I__2595\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17810\
        );

    \I__2594\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17810\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__17817\,
            I => \N__17807\
        );

    \I__2592\ : InMux
    port map (
            O => \N__17816\,
            I => \N__17802\
        );

    \I__2591\ : InMux
    port map (
            O => \N__17815\,
            I => \N__17802\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__17810\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__17807\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__17802\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__2586\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__17789\,
            I => \N__17784\
        );

    \I__2584\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17779\
        );

    \I__2583\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17779\
        );

    \I__2582\ : Span4Mux_v
    port map (
            O => \N__17784\,
            I => \N__17776\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__17779\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__17776\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__2579\ : InMux
    port map (
            O => \N__17771\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__2578\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17764\
        );

    \I__2577\ : InMux
    port map (
            O => \N__17767\,
            I => \N__17761\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__17764\,
            I => \VPP_VDDQ.count_2_1_3\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__17761\,
            I => \VPP_VDDQ.count_2_1_3\
        );

    \I__2574\ : InMux
    port map (
            O => \N__17756\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__2573\ : InMux
    port map (
            O => \N__17753\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__2572\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17746\
        );

    \I__2571\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17743\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__17746\,
            I => \VPP_VDDQ.count_2_1_5\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__17743\,
            I => \VPP_VDDQ.count_2_1_5\
        );

    \I__2568\ : InMux
    port map (
            O => \N__17738\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__2567\ : InMux
    port map (
            O => \N__17735\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__2566\ : CEMux
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__2564\ : Span4Mux_h
    port map (
            O => \N__17726\,
            I => \N__17723\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__17723\,
            I => \RSMRST_PWRGD.N_92_1\
        );

    \I__2562\ : InMux
    port map (
            O => \N__17720\,
            I => \N__17717\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__17714\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__2559\ : InMux
    port map (
            O => \N__17711\,
            I => \HDA_STRAP.un1_count_1_cry_13\
        );

    \I__2558\ : InMux
    port map (
            O => \N__17708\,
            I => \HDA_STRAP.un1_count_1_cry_14\
        );

    \I__2557\ : InMux
    port map (
            O => \N__17705\,
            I => \bfn_5_3_0_\
        );

    \I__2556\ : InMux
    port map (
            O => \N__17702\,
            I => \HDA_STRAP.un1_count_1_cry_16\
        );

    \I__2555\ : InMux
    port map (
            O => \N__17699\,
            I => \HDA_STRAP.un1_count_1_cry_4\
        );

    \I__2554\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__17693\,
            I => \HDA_STRAP.un1_count_1_cry_5_THRU_CO\
        );

    \I__2552\ : InMux
    port map (
            O => \N__17690\,
            I => \HDA_STRAP.un1_count_1_cry_5\
        );

    \I__2551\ : InMux
    port map (
            O => \N__17687\,
            I => \HDA_STRAP.un1_count_1_cry_6\
        );

    \I__2550\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__17681\,
            I => \HDA_STRAP.un1_count_1_cry_7_THRU_CO\
        );

    \I__2548\ : InMux
    port map (
            O => \N__17678\,
            I => \bfn_5_2_0_\
        );

    \I__2547\ : InMux
    port map (
            O => \N__17675\,
            I => \HDA_STRAP.un1_count_1_cry_8\
        );

    \I__2546\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__17669\,
            I => \HDA_STRAP.un1_count_1_cry_9_THRU_CO\
        );

    \I__2544\ : InMux
    port map (
            O => \N__17666\,
            I => \HDA_STRAP.un1_count_1_cry_9\
        );

    \I__2543\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17660\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__17660\,
            I => \HDA_STRAP.un1_count_1_cry_10_THRU_CO\
        );

    \I__2541\ : InMux
    port map (
            O => \N__17657\,
            I => \HDA_STRAP.un1_count_1_cry_10\
        );

    \I__2540\ : InMux
    port map (
            O => \N__17654\,
            I => \HDA_STRAP.un1_count_1_cry_11\
        );

    \I__2539\ : InMux
    port map (
            O => \N__17651\,
            I => \HDA_STRAP.un1_count_1_cry_12\
        );

    \I__2538\ : InMux
    port map (
            O => \N__17648\,
            I => \N__17645\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__17645\,
            I => \N__17641\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__17644\,
            I => \N__17637\
        );

    \I__2535\ : Span4Mux_v
    port map (
            O => \N__17641\,
            I => \N__17634\
        );

    \I__2534\ : InMux
    port map (
            O => \N__17640\,
            I => \N__17631\
        );

    \I__2533\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17628\
        );

    \I__2532\ : Odrv4
    port map (
            O => \N__17634\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__17631\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__17628\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__2528\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17615\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__17615\,
            I => \POWERLED.N_5050_i\
        );

    \I__2526\ : InMux
    port map (
            O => \N__17612\,
            I => \bfn_4_16_0_\
        );

    \I__2525\ : InMux
    port map (
            O => \N__17609\,
            I => \N__17604\
        );

    \I__2524\ : InMux
    port map (
            O => \N__17608\,
            I => \N__17598\
        );

    \I__2523\ : InMux
    port map (
            O => \N__17607\,
            I => \N__17598\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__17604\,
            I => \N__17595\
        );

    \I__2521\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17592\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__17598\,
            I => \N__17589\
        );

    \I__2519\ : Span4Mux_v
    port map (
            O => \N__17595\,
            I => \N__17586\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__17592\,
            I => \N__17583\
        );

    \I__2517\ : Span4Mux_s3_h
    port map (
            O => \N__17589\,
            I => \N__17580\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__17586\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2515\ : Odrv12
    port map (
            O => \N__17583\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__17580\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__17570\,
            I => \POWERLED.mult1_un89_sum_i_8\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__2510\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__17561\,
            I => \POWERLED.mult1_un68_sum_i_8\
        );

    \I__2508\ : InMux
    port map (
            O => \N__17558\,
            I => \HDA_STRAP.un1_count_1_cry_0\
        );

    \I__2507\ : InMux
    port map (
            O => \N__17555\,
            I => \HDA_STRAP.un1_count_1_cry_1\
        );

    \I__2506\ : InMux
    port map (
            O => \N__17552\,
            I => \HDA_STRAP.un1_count_1_cry_2\
        );

    \I__2505\ : InMux
    port map (
            O => \N__17549\,
            I => \HDA_STRAP.un1_count_1_cry_3\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__2503\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__17537\,
            I => \POWERLED.mult1_un110_sum_i_8\
        );

    \I__2500\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__17531\,
            I => \N__17527\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__17530\,
            I => \N__17523\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__17527\,
            I => \N__17520\
        );

    \I__2496\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17517\
        );

    \I__2495\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17514\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__17520\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__17517\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__17514\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__2491\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17504\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__17504\,
            I => \POWERLED.N_5043_i\
        );

    \I__2489\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17498\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__17498\,
            I => \N__17494\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__17497\,
            I => \N__17490\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__17494\,
            I => \N__17487\
        );

    \I__2485\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17484\
        );

    \I__2484\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17481\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__17487\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__17484\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__17481\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__2480\ : InMux
    port map (
            O => \N__17474\,
            I => \N__17471\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__17471\,
            I => \POWERLED.N_5044_i\
        );

    \I__2478\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__17465\,
            I => \N__17461\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__17464\,
            I => \N__17458\
        );

    \I__2475\ : Span4Mux_s3_v
    port map (
            O => \N__17461\,
            I => \N__17455\
        );

    \I__2474\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17451\
        );

    \I__2473\ : Span4Mux_v
    port map (
            O => \N__17455\,
            I => \N__17448\
        );

    \I__2472\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17445\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__17451\,
            I => \N__17442\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__17448\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__17445\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__17442\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__2466\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__17423\,
            I => \POWERLED.mult1_un96_sum_i_8\
        );

    \I__2462\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17417\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__17417\,
            I => \POWERLED.N_5045_i\
        );

    \I__2460\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__17411\,
            I => \N__17407\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__17410\,
            I => \N__17404\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__17407\,
            I => \N__17400\
        );

    \I__2456\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17397\
        );

    \I__2455\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17394\
        );

    \I__2454\ : Span4Mux_h
    port map (
            O => \N__17400\,
            I => \N__17389\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__17397\,
            I => \N__17389\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__17394\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__17389\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__2449\ : InMux
    port map (
            O => \N__17381\,
            I => \N__17378\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__17378\,
            I => \POWERLED.N_5046_i\
        );

    \I__2447\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17368\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__17368\,
            I => \N__17361\
        );

    \I__2443\ : InMux
    port map (
            O => \N__17365\,
            I => \N__17358\
        );

    \I__2442\ : InMux
    port map (
            O => \N__17364\,
            I => \N__17355\
        );

    \I__2441\ : Span4Mux_h
    port map (
            O => \N__17361\,
            I => \N__17350\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__17358\,
            I => \N__17350\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__17355\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__17350\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__17345\,
            I => \N__17342\
        );

    \I__2436\ : InMux
    port map (
            O => \N__17342\,
            I => \N__17339\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__17339\,
            I => \N__17336\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__17336\,
            I => \POWERLED.N_5047_i\
        );

    \I__2433\ : InMux
    port map (
            O => \N__17333\,
            I => \N__17330\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__17330\,
            I => \N__17325\
        );

    \I__2431\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17322\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__17328\,
            I => \N__17319\
        );

    \I__2429\ : Span4Mux_v
    port map (
            O => \N__17325\,
            I => \N__17316\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__17322\,
            I => \N__17313\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17310\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__17316\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__17313\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__17310\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__2423\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__17300\,
            I => \POWERLED.N_5048_i\
        );

    \I__2421\ : InMux
    port map (
            O => \N__17297\,
            I => \N__17294\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__17294\,
            I => \N__17289\
        );

    \I__2419\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17286\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__17292\,
            I => \N__17283\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__17289\,
            I => \N__17280\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__17286\,
            I => \N__17277\
        );

    \I__2415\ : InMux
    port map (
            O => \N__17283\,
            I => \N__17274\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__17280\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__17277\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__17274\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2411\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__17264\,
            I => \POWERLED.N_5049_i\
        );

    \I__2409\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17258\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__17255\,
            I => \N__17248\
        );

    \I__2406\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17241\
        );

    \I__2405\ : InMux
    port map (
            O => \N__17253\,
            I => \N__17241\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17252\,
            I => \N__17241\
        );

    \I__2403\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17238\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__17248\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__17241\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__17238\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__2398\ : InMux
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__17225\,
            I => \POWERLED.un1_count_cry_0_i\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__17219\,
            I => \N__17215\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__17218\,
            I => \N__17211\
        );

    \I__2393\ : Span12Mux_s6_v
    port map (
            O => \N__17215\,
            I => \N__17208\
        );

    \I__2392\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17205\
        );

    \I__2391\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17202\
        );

    \I__2390\ : Odrv12
    port map (
            O => \N__17208\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__17205\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__17202\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__2386\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__17186\,
            I => \POWERLED.N_5036_i\
        );

    \I__2383\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__17180\,
            I => \N__17176\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__2380\ : Span4Mux_s3_v
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__2379\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17166\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__17170\,
            I => \N__17163\
        );

    \I__2377\ : InMux
    port map (
            O => \N__17169\,
            I => \N__17160\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__17166\,
            I => \N__17157\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__17163\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__17160\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__17157\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__17150\,
            I => \N__17147\
        );

    \I__2371\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17144\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__17144\,
            I => \POWERLED.N_5037_i\
        );

    \I__2369\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17137\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__17140\,
            I => \N__17134\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__2366\ : InMux
    port map (
            O => \N__17134\,
            I => \N__17127\
        );

    \I__2365\ : Span12Mux_s7_v
    port map (
            O => \N__17131\,
            I => \N__17124\
        );

    \I__2364\ : InMux
    port map (
            O => \N__17130\,
            I => \N__17121\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__17127\,
            I => \N__17118\
        );

    \I__2362\ : Odrv12
    port map (
            O => \N__17124\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__17121\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__17118\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__2358\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__17105\,
            I => \POWERLED.N_5038_i\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17099\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__17099\,
            I => \N__17095\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__17098\,
            I => \N__17091\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__17095\,
            I => \N__17088\
        );

    \I__2352\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17085\
        );

    \I__2351\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17082\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__17088\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__17085\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__17082\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__17075\,
            I => \N__17072\
        );

    \I__2346\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17069\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__17069\,
            I => \POWERLED.N_5039_i\
        );

    \I__2344\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__17063\,
            I => \N__17060\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__17060\,
            I => \N__17055\
        );

    \I__2341\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17052\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__17058\,
            I => \N__17049\
        );

    \I__2339\ : Span4Mux_h
    port map (
            O => \N__17055\,
            I => \N__17046\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__17052\,
            I => \N__17043\
        );

    \I__2337\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17040\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__17046\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__17043\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__17040\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__17033\,
            I => \N__17030\
        );

    \I__2332\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17027\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__17027\,
            I => \POWERLED.N_5040_i\
        );

    \I__2330\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__17021\,
            I => \N__17016\
        );

    \I__2328\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17013\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__17019\,
            I => \N__17010\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__17016\,
            I => \N__17007\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__17013\,
            I => \N__17004\
        );

    \I__2324\ : InMux
    port map (
            O => \N__17010\,
            I => \N__17001\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__17007\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__17004\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__17001\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__2319\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__16985\,
            I => \POWERLED.N_5041_i\
        );

    \I__2316\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__16976\,
            I => \N__16971\
        );

    \I__2313\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16968\
        );

    \I__2312\ : InMux
    port map (
            O => \N__16974\,
            I => \N__16965\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__16971\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__16968\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__16965\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__2308\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__2306\ : Odrv12
    port map (
            O => \N__16952\,
            I => \POWERLED.mult1_un117_sum_i_8\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__16949\,
            I => \N__16946\
        );

    \I__2304\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__16943\,
            I => \POWERLED.N_5042_i\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__16940\,
            I => \POWERLED.mult1_un110_sum_s_8_cascade_\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__2300\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__16931\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__2298\ : InMux
    port map (
            O => \N__16928\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__2297\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__16922\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__2295\ : InMux
    port map (
            O => \N__16919\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__2293\ : InMux
    port map (
            O => \N__16913\,
            I => \N__16910\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__16910\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__2291\ : InMux
    port map (
            O => \N__16907\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__2290\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__16901\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__2288\ : InMux
    port map (
            O => \N__16898\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__2286\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__16889\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__2284\ : InMux
    port map (
            O => \N__16886\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__2283\ : InMux
    port map (
            O => \N__16883\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \POWERLED.mult1_un103_sum_s_8_cascade_\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__16877\,
            I => \N__16873\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__16876\,
            I => \N__16869\
        );

    \I__2279\ : InMux
    port map (
            O => \N__16873\,
            I => \N__16862\
        );

    \I__2278\ : InMux
    port map (
            O => \N__16872\,
            I => \N__16862\
        );

    \I__2277\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16862\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__16862\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__16859\,
            I => \N__16855\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__16858\,
            I => \N__16851\
        );

    \I__2273\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16844\
        );

    \I__2272\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16844\
        );

    \I__2271\ : InMux
    port map (
            O => \N__16851\,
            I => \N__16844\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__16844\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__2268\ : InMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__16835\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__2266\ : InMux
    port map (
            O => \N__16832\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__2265\ : InMux
    port map (
            O => \N__16829\,
            I => \N__16826\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__16826\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__2263\ : InMux
    port map (
            O => \N__16823\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__2262\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__16817\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__2260\ : InMux
    port map (
            O => \N__16814\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__2259\ : InMux
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__16808\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__2257\ : InMux
    port map (
            O => \N__16805\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__2256\ : InMux
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__16799\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__2254\ : InMux
    port map (
            O => \N__16796\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__2253\ : InMux
    port map (
            O => \N__16793\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__16790\,
            I => \N__16786\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__16789\,
            I => \N__16783\
        );

    \I__2250\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16778\
        );

    \I__2249\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16773\
        );

    \I__2248\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16773\
        );

    \I__2247\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16770\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__16778\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__16773\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__16770\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2243\ : InMux
    port map (
            O => \N__16763\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__2242\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__16757\,
            I => \POWERLED.mult1_un124_sum_axb_7_l_fx\
        );

    \I__2240\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__16751\,
            I => \N__16747\
        );

    \I__2238\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16744\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__16747\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__16744\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__2235\ : InMux
    port map (
            O => \N__16739\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__16736\,
            I => \N__16733\
        );

    \I__2233\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__16730\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__2231\ : InMux
    port map (
            O => \N__16727\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__2230\ : InMux
    port map (
            O => \N__16724\,
            I => \N__16721\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__16721\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__2228\ : InMux
    port map (
            O => \N__16718\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__2226\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16706\
        );

    \I__2225\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16706\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__16706\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__2223\ : InMux
    port map (
            O => \N__16703\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__2222\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16697\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__16697\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__2220\ : InMux
    port map (
            O => \N__16694\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__2219\ : InMux
    port map (
            O => \N__16691\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__2218\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__16685\,
            I => \N__16679\
        );

    \I__2216\ : InMux
    port map (
            O => \N__16684\,
            I => \N__16674\
        );

    \I__2215\ : InMux
    port map (
            O => \N__16683\,
            I => \N__16674\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__16682\,
            I => \N__16671\
        );

    \I__2213\ : Span12Mux_s4_v
    port map (
            O => \N__16679\,
            I => \N__16665\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__16674\,
            I => \N__16662\
        );

    \I__2211\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16655\
        );

    \I__2210\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16655\
        );

    \I__2209\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16655\
        );

    \I__2208\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16652\
        );

    \I__2207\ : Odrv12
    port map (
            O => \N__16665\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__16662\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__16655\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__16652\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__2203\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__16640\,
            I => \N__16637\
        );

    \I__2201\ : Span4Mux_v
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__16634\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \N__16628\
        );

    \I__2198\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16625\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__2196\ : Odrv12
    port map (
            O => \N__16622\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__2195\ : InMux
    port map (
            O => \N__16619\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__2193\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__16610\,
            I => \N__16607\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__16607\,
            I => \POWERLED.mult1_un124_sum_axb_4_l_fx\
        );

    \I__2190\ : InMux
    port map (
            O => \N__16604\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__2189\ : InMux
    port map (
            O => \N__16601\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__2188\ : InMux
    port map (
            O => \N__16598\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__2187\ : InMux
    port map (
            O => \N__16595\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__2186\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__16589\,
            I => \VPP_VDDQ.count_2_0_12\
        );

    \I__2184\ : InMux
    port map (
            O => \N__16586\,
            I => \N__16583\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__16583\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__2182\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__16577\,
            I => \VPP_VDDQ.count_2_0_14\
        );

    \I__2180\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__16571\,
            I => \N__16561\
        );

    \I__2178\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16556\
        );

    \I__2177\ : InMux
    port map (
            O => \N__16569\,
            I => \N__16556\
        );

    \I__2176\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16551\
        );

    \I__2175\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16551\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16544\
        );

    \I__2173\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16544\
        );

    \I__2172\ : InMux
    port map (
            O => \N__16564\,
            I => \N__16544\
        );

    \I__2171\ : Span4Mux_h
    port map (
            O => \N__16561\,
            I => \N__16539\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__16556\,
            I => \N__16539\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__16551\,
            I => \POWERLED.N_2305_i\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__16544\,
            I => \POWERLED.N_2305_i\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__16539\,
            I => \POWERLED.N_2305_i\
        );

    \I__2166\ : InMux
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__2164\ : Span4Mux_h
    port map (
            O => \N__16526\,
            I => \N__16522\
        );

    \I__2163\ : InMux
    port map (
            O => \N__16525\,
            I => \N__16519\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__16522\,
            I => \N__16516\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__16519\,
            I => \POWERLED.N_660\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__16516\,
            I => \POWERLED.N_660\
        );

    \I__2159\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16508\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__16502\,
            I => \POWERLED.curr_state_1_0\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__16499\,
            I => \N__16496\
        );

    \I__2154\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16488\
        );

    \I__2153\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16485\
        );

    \I__2152\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16482\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16479\
        );

    \I__2150\ : InMux
    port map (
            O => \N__16492\,
            I => \N__16476\
        );

    \I__2149\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16473\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__16488\,
            I => \N__16470\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__16485\,
            I => \N__16458\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__16482\,
            I => \N__16455\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__16479\,
            I => \N__16452\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__16476\,
            I => \N__16449\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__16473\,
            I => \N__16446\
        );

    \I__2142\ : Glb2LocalMux
    port map (
            O => \N__16470\,
            I => \N__16415\
        );

    \I__2141\ : CEMux
    port map (
            O => \N__16469\,
            I => \N__16415\
        );

    \I__2140\ : CEMux
    port map (
            O => \N__16468\,
            I => \N__16415\
        );

    \I__2139\ : CEMux
    port map (
            O => \N__16467\,
            I => \N__16415\
        );

    \I__2138\ : CEMux
    port map (
            O => \N__16466\,
            I => \N__16415\
        );

    \I__2137\ : CEMux
    port map (
            O => \N__16465\,
            I => \N__16415\
        );

    \I__2136\ : CEMux
    port map (
            O => \N__16464\,
            I => \N__16415\
        );

    \I__2135\ : CEMux
    port map (
            O => \N__16463\,
            I => \N__16415\
        );

    \I__2134\ : CEMux
    port map (
            O => \N__16462\,
            I => \N__16415\
        );

    \I__2133\ : CEMux
    port map (
            O => \N__16461\,
            I => \N__16415\
        );

    \I__2132\ : Glb2LocalMux
    port map (
            O => \N__16458\,
            I => \N__16415\
        );

    \I__2131\ : Glb2LocalMux
    port map (
            O => \N__16455\,
            I => \N__16415\
        );

    \I__2130\ : Glb2LocalMux
    port map (
            O => \N__16452\,
            I => \N__16415\
        );

    \I__2129\ : Glb2LocalMux
    port map (
            O => \N__16449\,
            I => \N__16415\
        );

    \I__2128\ : Glb2LocalMux
    port map (
            O => \N__16446\,
            I => \N__16415\
        );

    \I__2127\ : GlobalMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__2126\ : gio2CtrlBuf
    port map (
            O => \N__16412\,
            I => \N_557_g\
        );

    \I__2125\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__16403\,
            I => \N__16397\
        );

    \I__2122\ : InMux
    port map (
            O => \N__16402\,
            I => \N__16390\
        );

    \I__2121\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16390\
        );

    \I__2120\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16390\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__16397\,
            I => \N_639\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__16390\,
            I => \N_639\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16381\
        );

    \I__2116\ : InMux
    port map (
            O => \N__16384\,
            I => \N__16377\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__16381\,
            I => \N__16374\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__16380\,
            I => \N__16371\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__16377\,
            I => \N__16364\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__16374\,
            I => \N__16361\
        );

    \I__2111\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16350\
        );

    \I__2110\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16350\
        );

    \I__2109\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16350\
        );

    \I__2108\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16350\
        );

    \I__2107\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16350\
        );

    \I__2106\ : Span4Mux_h
    port map (
            O => \N__16364\,
            I => \N__16347\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__16361\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__16350\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__16347\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__16340\,
            I => \N__16337\
        );

    \I__2101\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16334\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__16331\,
            I => \N__16326\
        );

    \I__2098\ : InMux
    port map (
            O => \N__16330\,
            I => \N__16321\
        );

    \I__2097\ : InMux
    port map (
            O => \N__16329\,
            I => \N__16321\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__16326\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__16321\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__16316\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_\
        );

    \I__2093\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16310\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__16310\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__16307\,
            I => \VPP_VDDQ.count_2Z0Z_9_cascade_\
        );

    \I__2090\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16301\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__16301\,
            I => \VPP_VDDQ.un9_clk_100khz_7\
        );

    \I__2088\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16292\
        );

    \I__2087\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16292\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__16292\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__2085\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16286\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__16286\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__2083\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16280\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__16280\,
            I => \N__16277\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__16277\,
            I => \VPP_VDDQ.un9_clk_100khz_10\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__16274\,
            I => \VPP_VDDQ.count_2_1_1_cascade_\
        );

    \I__2079\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16268\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__16268\,
            I => \N__16264\
        );

    \I__2077\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16261\
        );

    \I__2076\ : Span4Mux_v
    port map (
            O => \N__16264\,
            I => \N__16258\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__16261\,
            I => \N__16255\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__16258\,
            I => \N__16252\
        );

    \I__2073\ : IoSpan4Mux
    port map (
            O => \N__16255\,
            I => \N__16249\
        );

    \I__2072\ : Span4Mux_h
    port map (
            O => \N__16252\,
            I => \N__16246\
        );

    \I__2071\ : IoSpan4Mux
    port map (
            O => \N__16249\,
            I => \N__16243\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__16246\,
            I => slp_susn
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__16243\,
            I => slp_susn
        );

    \I__2068\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16235\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__16235\,
            I => \N__16232\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__16232\,
            I => \N__16229\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__16229\,
            I => v5a_ok
        );

    \I__2064\ : IoInMux
    port map (
            O => \N__16226\,
            I => \N__16222\
        );

    \I__2063\ : IoInMux
    port map (
            O => \N__16225\,
            I => \N__16218\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__16222\,
            I => \N__16215\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__16221\,
            I => \N__16212\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__16218\,
            I => \N__16209\
        );

    \I__2059\ : Span4Mux_s3_h
    port map (
            O => \N__16215\,
            I => \N__16206\
        );

    \I__2058\ : InMux
    port map (
            O => \N__16212\,
            I => \N__16203\
        );

    \I__2057\ : IoSpan4Mux
    port map (
            O => \N__16209\,
            I => \N__16200\
        );

    \I__2056\ : Sp12to4
    port map (
            O => \N__16206\,
            I => \N__16195\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__16203\,
            I => \N__16195\
        );

    \I__2054\ : IoSpan4Mux
    port map (
            O => \N__16200\,
            I => \N__16192\
        );

    \I__2053\ : Span12Mux_v
    port map (
            O => \N__16195\,
            I => \N__16189\
        );

    \I__2052\ : IoSpan4Mux
    port map (
            O => \N__16192\,
            I => \N__16186\
        );

    \I__2051\ : Odrv12
    port map (
            O => \N__16189\,
            I => v33a_ok
        );

    \I__2050\ : Odrv4
    port map (
            O => \N__16186\,
            I => v33a_ok
        );

    \I__2049\ : IoInMux
    port map (
            O => \N__16181\,
            I => \N__16178\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__16178\,
            I => \N__16174\
        );

    \I__2047\ : InMux
    port map (
            O => \N__16177\,
            I => \N__16171\
        );

    \I__2046\ : Span4Mux_s2_h
    port map (
            O => \N__16174\,
            I => \N__16168\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__16171\,
            I => \N__16165\
        );

    \I__2044\ : Sp12to4
    port map (
            O => \N__16168\,
            I => \N__16162\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__16165\,
            I => \N__16159\
        );

    \I__2042\ : Span12Mux_s11_v
    port map (
            O => \N__16162\,
            I => \N__16156\
        );

    \I__2041\ : Span4Mux_v
    port map (
            O => \N__16159\,
            I => \N__16153\
        );

    \I__2040\ : Odrv12
    port map (
            O => \N__16156\,
            I => v1p8a_ok
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__16153\,
            I => v1p8a_ok
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__16148\,
            I => \rsmrst_pwrgd_signal_cascade_\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__16145\,
            I => \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__16142\,
            I => \N__16138\
        );

    \I__2035\ : InMux
    port map (
            O => \N__16141\,
            I => \N__16135\
        );

    \I__2034\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16132\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__16135\,
            I => \N__16127\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__16132\,
            I => \N__16127\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__16124\,
            I => \N__16121\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__16121\,
            I => \RSMRST_PWRGD.N_264_i\
        );

    \I__2028\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16115\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__16115\,
            I => \VPP_VDDQ.un9_clk_100khz_1\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__16112\,
            I => \VPP_VDDQ.un9_clk_100khz_13_cascade_\
        );

    \I__2025\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16103\
        );

    \I__2024\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16103\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__16103\,
            I => \N__16099\
        );

    \I__2022\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16096\
        );

    \I__2021\ : Span4Mux_s3_h
    port map (
            O => \N__16099\,
            I => \N__16093\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__16096\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__16093\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__2018\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16084\
        );

    \I__2017\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16080\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__16084\,
            I => \N__16077\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__16083\,
            I => \N__16074\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__16080\,
            I => \N__16070\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__16077\,
            I => \N__16067\
        );

    \I__2012\ : InMux
    port map (
            O => \N__16074\,
            I => \N__16064\
        );

    \I__2011\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16061\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__16070\,
            I => \N__16058\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__16067\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__16064\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__16061\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__16058\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__16049\,
            I => \VPP_VDDQ.N_1_i_cascade_\
        );

    \I__2004\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16040\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16045\,
            I => \N__16040\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__16040\,
            I => \N__16037\
        );

    \I__2001\ : Span4Mux_s3_h
    port map (
            O => \N__16037\,
            I => \N__16034\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__16034\,
            I => \VPP_VDDQ.N_664\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__16031\,
            I => \VPP_VDDQ.count_2_1_sqmuxa_cascade_\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__16028\,
            I => \VPP_VDDQ.count_2_1_0_cascade_\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__16025\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__1996\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__16019\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__1994\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16013\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__16013\,
            I => \VPP_VDDQ.count_2_1_1\
        );

    \I__1992\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16004\
        );

    \I__1991\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16004\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__16004\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__1989\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__1987\ : Span4Mux_v
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__15992\,
            I => \N__15989\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__15989\,
            I => gpio_fpga_soc_1
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__15986\,
            I => \HDA_STRAP.m14_i_0_cascade_\
        );

    \I__1983\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15977\
        );

    \I__1982\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15977\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__15977\,
            I => \N__15974\
        );

    \I__1980\ : Span4Mux_v
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__15971\,
            I => \N__15966\
        );

    \I__1978\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15963\
        );

    \I__1977\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15960\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__15966\,
            I => \N_428\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__15963\,
            I => \N_428\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__15960\,
            I => \N_428\
        );

    \I__1973\ : InMux
    port map (
            O => \N__15953\,
            I => \N__15938\
        );

    \I__1972\ : InMux
    port map (
            O => \N__15952\,
            I => \N__15938\
        );

    \I__1971\ : InMux
    port map (
            O => \N__15951\,
            I => \N__15938\
        );

    \I__1970\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15938\
        );

    \I__1969\ : InMux
    port map (
            O => \N__15949\,
            I => \N__15938\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__15938\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1967\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15927\
        );

    \I__1966\ : InMux
    port map (
            O => \N__15934\,
            I => \N__15927\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__15933\,
            I => \N__15924\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__15932\,
            I => \N__15921\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__15927\,
            I => \N__15917\
        );

    \I__1962\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15910\
        );

    \I__1961\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15910\
        );

    \I__1960\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15910\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__15917\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__15910\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1957\ : InMux
    port map (
            O => \N__15905\,
            I => \N__15901\
        );

    \I__1956\ : InMux
    port map (
            O => \N__15904\,
            I => \N__15898\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__15901\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__15898\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1953\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15890\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__15890\,
            I => \HDA_STRAP.HDA_SDO_ATP_3_0\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__15887\,
            I => \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_\
        );

    \I__1950\ : IoInMux
    port map (
            O => \N__15884\,
            I => \N__15881\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__15881\,
            I => \N__15878\
        );

    \I__1948\ : Span4Mux_s3_h
    port map (
            O => \N__15878\,
            I => \N__15875\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__15875\,
            I => \N__15872\
        );

    \I__1946\ : Odrv4
    port map (
            O => \N__15872\,
            I => hda_sdo_atp
        );

    \I__1945\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15866\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15863\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__15863\,
            I => \N__15859\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__15862\,
            I => \N__15856\
        );

    \I__1941\ : Span4Mux_h
    port map (
            O => \N__15859\,
            I => \N__15853\
        );

    \I__1940\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15850\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__15853\,
            I => \PCH_PWRGD.N_670\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__15850\,
            I => \PCH_PWRGD.N_670\
        );

    \I__1937\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15842\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__15842\,
            I => \N__15836\
        );

    \I__1935\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15828\
        );

    \I__1934\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15828\
        );

    \I__1933\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15828\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__15836\,
            I => \N__15825\
        );

    \I__1931\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15822\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__15828\,
            I => \PCH_PWRGD.N_2266_i\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__15825\,
            I => \PCH_PWRGD.N_2266_i\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__15822\,
            I => \PCH_PWRGD.N_2266_i\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__1926\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15809\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__15809\,
            I => \PCH_PWRGD.N_38_f0\
        );

    \I__1924\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15802\
        );

    \I__1923\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15799\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__15802\,
            I => \N__15793\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__15799\,
            I => \N__15793\
        );

    \I__1920\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15790\
        );

    \I__1919\ : Span12Mux_s6_v
    port map (
            O => \N__15793\,
            I => \N__15787\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__15790\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__15787\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__15782\,
            I => \PCH_PWRGD.N_38_f0_cascade_\
        );

    \I__1915\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15775\
        );

    \I__1914\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15772\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__15775\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__15772\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__15767\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__15764\,
            I => \HDA_STRAP.N_16_cascade_\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__15761\,
            I => \PCH_PWRGD.delayed_vccin_okZ0_cascade_\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__15758\,
            I => \N_428_cascade_\
        );

    \I__1907\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15749\
        );

    \I__1906\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15749\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__15749\,
            I => \POWERLED.count_1_5\
        );

    \I__1904\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__15743\,
            I => \POWERLED.count_0_5\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__1901\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15731\
        );

    \I__1900\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15731\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__15731\,
            I => \POWERLED.count_1_14\
        );

    \I__1898\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15725\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__15725\,
            I => \POWERLED.count_0_14\
        );

    \I__1896\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15716\
        );

    \I__1895\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15716\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__15716\,
            I => \POWERLED.count_1_6\
        );

    \I__1893\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15710\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__15710\,
            I => \POWERLED.count_0_6\
        );

    \I__1891\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15703\
        );

    \I__1890\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15700\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__15703\,
            I => \N__15697\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__15700\,
            I => \POWERLED.count_1_10\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__15697\,
            I => \POWERLED.count_1_10\
        );

    \I__1886\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__1884\ : Span4Mux_s2_h
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__15683\,
            I => \POWERLED.count_0_10\
        );

    \I__1882\ : IoInMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__1880\ : Span4Mux_s1_h
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__15671\,
            I => v33a_enn
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__1877\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15659\
        );

    \I__1876\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15659\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__15659\,
            I => \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0\
        );

    \I__1874\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__15653\,
            I => \POWERLED.count_0_15\
        );

    \I__1872\ : InMux
    port map (
            O => \N__15650\,
            I => \N__15644\
        );

    \I__1871\ : InMux
    port map (
            O => \N__15649\,
            I => \N__15644\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__15644\,
            I => \POWERLED.count_1_7\
        );

    \I__1869\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__15638\,
            I => \POWERLED.count_0_7\
        );

    \I__1867\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15629\
        );

    \I__1866\ : InMux
    port map (
            O => \N__15634\,
            I => \N__15629\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__15629\,
            I => \POWERLED.count_1_8\
        );

    \I__1864\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15623\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__15623\,
            I => \POWERLED.count_0_8\
        );

    \I__1862\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15614\
        );

    \I__1861\ : InMux
    port map (
            O => \N__15619\,
            I => \N__15614\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__15614\,
            I => \POWERLED.count_1_9\
        );

    \I__1859\ : InMux
    port map (
            O => \N__15611\,
            I => \N__15608\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__15608\,
            I => \POWERLED.count_0_9\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__15605\,
            I => \N__15602\
        );

    \I__1856\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15596\
        );

    \I__1855\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15596\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__15596\,
            I => \POWERLED.count_1_13\
        );

    \I__1853\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15590\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__15590\,
            I => \POWERLED.count_0_13\
        );

    \I__1851\ : SRMux
    port map (
            O => \N__15587\,
            I => \N__15584\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__15584\,
            I => \N__15581\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__15581\,
            I => \N__15578\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__15578\,
            I => \POWERLED.pwm_out_1_sqmuxa\
        );

    \I__1847\ : InMux
    port map (
            O => \N__15575\,
            I => \N__15572\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__15572\,
            I => \POWERLED.un79_clk_100khzlt6\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__15569\,
            I => \POWERLED.un79_clk_100khzlto15_5_cascade_\
        );

    \I__1844\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__15563\,
            I => \POWERLED.un79_clk_100khzlto15_4\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__15560\,
            I => \POWERLED.un79_clk_100khzlto15_7_cascade_\
        );

    \I__1841\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__15554\,
            I => \N__15549\
        );

    \I__1839\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15546\
        );

    \I__1838\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15543\
        );

    \I__1837\ : Span4Mux_s1_h
    port map (
            O => \N__15549\,
            I => \N__15538\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__15546\,
            I => \N__15538\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__15543\,
            I => \POWERLED.un79_clk_100khz\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__15538\,
            I => \POWERLED.un79_clk_100khz\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__15533\,
            I => \POWERLED.un79_clk_100khz_cascade_\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__15530\,
            I => \N__15527\
        );

    \I__1831\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15524\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__15524\,
            I => \N__15521\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__15521\,
            I => \POWERLED.g0_2_1\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__15518\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__15515\,
            I => \VPP_VDDQ.N_60_cascade_\
        );

    \I__1826\ : SRMux
    port map (
            O => \N__15512\,
            I => \N__15509\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__15509\,
            I => \N__15506\
        );

    \I__1824\ : Span4Mux_s2_h
    port map (
            O => \N__15506\,
            I => \N__15503\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__15503\,
            I => \VPP_VDDQ.N_60_i\
        );

    \I__1822\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15493\
        );

    \I__1821\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15493\
        );

    \I__1820\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15490\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__15493\,
            I => \VPP_VDDQ.N_60\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__15490\,
            I => \VPP_VDDQ.N_60\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__15485\,
            I => \N__15481\
        );

    \I__1816\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15476\
        );

    \I__1815\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15476\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__15476\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__1813\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15467\
        );

    \I__1812\ : InMux
    port map (
            O => \N__15472\,
            I => \N__15467\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__15467\,
            I => \VPP_VDDQ.delayed_vddq_ok_en\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__15464\,
            I => \VPP_VDDQ_delayed_vddq_ok_cascade_\
        );

    \I__1809\ : IoInMux
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__1807\ : Span4Mux_s0_v
    port map (
            O => \N__15455\,
            I => \N__15452\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__15449\,
            I => \N__15446\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__15446\,
            I => vccst_pwrgd
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__15443\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_\
        );

    \I__1802\ : IoInMux
    port map (
            O => \N__15440\,
            I => \N__15436\
        );

    \I__1801\ : IoInMux
    port map (
            O => \N__15439\,
            I => \N__15433\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__15436\,
            I => \N__15430\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__15433\,
            I => \N__15427\
        );

    \I__1798\ : Span4Mux_s1_h
    port map (
            O => \N__15430\,
            I => \N__15424\
        );

    \I__1797\ : Span12Mux_s10_h
    port map (
            O => \N__15427\,
            I => \N__15421\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__15424\,
            I => \N__15418\
        );

    \I__1795\ : Odrv12
    port map (
            O => \N__15421\,
            I => pch_pwrok
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__15418\,
            I => pch_pwrok
        );

    \I__1793\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15410\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__15410\,
            I => \PCH_PWRGD.curr_state_7_0\
        );

    \I__1791\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15403\
        );

    \I__1790\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__15403\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__15400\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__15395\,
            I => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__1786\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15383\
        );

    \I__1785\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15383\
        );

    \I__1784\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15383\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__15383\,
            I => \PCH_PWRGD.N_655\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__15380\,
            I => \N__15376\
        );

    \I__1781\ : InMux
    port map (
            O => \N__15379\,
            I => \N__15370\
        );

    \I__1780\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15361\
        );

    \I__1779\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15361\
        );

    \I__1778\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15361\
        );

    \I__1777\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15361\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__15370\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__15361\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15340\
        );

    \I__1773\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15340\
        );

    \I__1772\ : InMux
    port map (
            O => \N__15354\,
            I => \N__15340\
        );

    \I__1771\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15340\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__15352\,
            I => \N__15337\
        );

    \I__1769\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15331\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__15350\,
            I => \N__15325\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__15349\,
            I => \N__15320\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15316\
        );

    \I__1765\ : InMux
    port map (
            O => \N__15337\,
            I => \N__15307\
        );

    \I__1764\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15307\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15307\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15307\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15331\,
            I => \N__15304\
        );

    \I__1760\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15299\
        );

    \I__1759\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15299\
        );

    \I__1758\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15296\
        );

    \I__1757\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15285\
        );

    \I__1756\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15285\
        );

    \I__1755\ : InMux
    port map (
            O => \N__15323\,
            I => \N__15285\
        );

    \I__1754\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15285\
        );

    \I__1753\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15285\
        );

    \I__1752\ : Span4Mux_s1_h
    port map (
            O => \N__15316\,
            I => \N__15280\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__15307\,
            I => \N__15280\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__15304\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__15299\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__15296\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__15285\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__15280\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__15269\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa_cascade_\
        );

    \I__1744\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15263\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__15263\,
            I => \PCH_PWRGD.curr_state_0_0\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__15260\,
            I => \VPP_VDDQ.N_53_cascade_\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\
        );

    \I__1740\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15251\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__15251\,
            I => \VPP_VDDQ.curr_state_2_0_1\
        );

    \I__1738\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15245\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__15245\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__15242\,
            I => \VPP_VDDQ.m4_0_0_cascade_\
        );

    \I__1735\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__15236\,
            I => \PCH_PWRGD.count_1_i_a2_2_0\
        );

    \I__1733\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15230\,
            I => \N__15225\
        );

    \I__1731\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15220\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15228\,
            I => \N__15220\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__15225\,
            I => \PCH_PWRGD.count_1_i_a2_11_0\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__15220\,
            I => \PCH_PWRGD.count_1_i_a2_11_0\
        );

    \I__1727\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15209\
        );

    \I__1726\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15209\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__15209\,
            I => \PCH_PWRGD.count_rst\
        );

    \I__1724\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__15203\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__1722\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15191\
        );

    \I__1721\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15191\
        );

    \I__1720\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15191\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__15191\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__1718\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15182\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15182\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__15182\,
            I => \PCH_PWRGD.count_0_13\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__15179\,
            I => \N__15175\
        );

    \I__1714\ : InMux
    port map (
            O => \N__15178\,
            I => \N__15171\
        );

    \I__1713\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15168\
        );

    \I__1712\ : InMux
    port map (
            O => \N__15174\,
            I => \N__15165\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__15171\,
            I => \N__15162\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__15168\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__15165\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__15162\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1707\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15152\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__15152\,
            I => \N__15148\
        );

    \I__1705\ : InMux
    port map (
            O => \N__15151\,
            I => \N__15145\
        );

    \I__1704\ : Odrv12
    port map (
            O => \N__15148\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__15145\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__1702\ : CEMux
    port map (
            O => \N__15140\,
            I => \N__15133\
        );

    \I__1701\ : CEMux
    port map (
            O => \N__15139\,
            I => \N__15127\
        );

    \I__1700\ : CEMux
    port map (
            O => \N__15138\,
            I => \N__15124\
        );

    \I__1699\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15119\
        );

    \I__1698\ : CEMux
    port map (
            O => \N__15136\,
            I => \N__15119\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__15133\,
            I => \N__15116\
        );

    \I__1696\ : CEMux
    port map (
            O => \N__15132\,
            I => \N__15113\
        );

    \I__1695\ : InMux
    port map (
            O => \N__15131\,
            I => \N__15108\
        );

    \I__1694\ : CEMux
    port map (
            O => \N__15130\,
            I => \N__15108\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__15127\,
            I => \N__15103\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__15124\,
            I => \N__15103\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__15119\,
            I => \N__15095\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__15116\,
            I => \N__15090\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__15113\,
            I => \N__15090\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__15108\,
            I => \N__15085\
        );

    \I__1687\ : Span4Mux_s3_v
    port map (
            O => \N__15103\,
            I => \N__15082\
        );

    \I__1686\ : InMux
    port map (
            O => \N__15102\,
            I => \N__15073\
        );

    \I__1685\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15073\
        );

    \I__1684\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15073\
        );

    \I__1683\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15073\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__15098\,
            I => \N__15061\
        );

    \I__1681\ : Span4Mux_h
    port map (
            O => \N__15095\,
            I => \N__15056\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__15090\,
            I => \N__15056\
        );

    \I__1679\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15048\
        );

    \I__1678\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15048\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__15085\,
            I => \N__15041\
        );

    \I__1676\ : Span4Mux_s1_h
    port map (
            O => \N__15082\,
            I => \N__15041\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__15073\,
            I => \N__15041\
        );

    \I__1674\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15036\
        );

    \I__1673\ : CEMux
    port map (
            O => \N__15071\,
            I => \N__15036\
        );

    \I__1672\ : CEMux
    port map (
            O => \N__15070\,
            I => \N__15033\
        );

    \I__1671\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15026\
        );

    \I__1670\ : InMux
    port map (
            O => \N__15068\,
            I => \N__15026\
        );

    \I__1669\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15026\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15066\,
            I => \N__15019\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15065\,
            I => \N__15019\
        );

    \I__1666\ : InMux
    port map (
            O => \N__15064\,
            I => \N__15019\
        );

    \I__1665\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15013\
        );

    \I__1664\ : Span4Mux_s0_h
    port map (
            O => \N__15056\,
            I => \N__15010\
        );

    \I__1663\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15003\
        );

    \I__1662\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15003\
        );

    \I__1661\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15003\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__15048\,
            I => \N__14998\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__15041\,
            I => \N__14998\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__15036\,
            I => \N__14989\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__15033\,
            I => \N__14989\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__15026\,
            I => \N__14989\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__15019\,
            I => \N__14989\
        );

    \I__1654\ : InMux
    port map (
            O => \N__15018\,
            I => \N__14984\
        );

    \I__1653\ : InMux
    port map (
            O => \N__15017\,
            I => \N__14984\
        );

    \I__1652\ : InMux
    port map (
            O => \N__15016\,
            I => \N__14981\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__15013\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__15010\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__15003\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__14998\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__1647\ : Odrv12
    port map (
            O => \N__14989\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__14984\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__14981\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__1644\ : SRMux
    port map (
            O => \N__14966\,
            I => \N__14962\
        );

    \I__1643\ : SRMux
    port map (
            O => \N__14965\,
            I => \N__14954\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__14962\,
            I => \N__14951\
        );

    \I__1641\ : SRMux
    port map (
            O => \N__14961\,
            I => \N__14948\
        );

    \I__1640\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14945\
        );

    \I__1639\ : SRMux
    port map (
            O => \N__14959\,
            I => \N__14942\
        );

    \I__1638\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14918\
        );

    \I__1637\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14918\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__14954\,
            I => \N__14913\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__14951\,
            I => \N__14908\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__14948\,
            I => \N__14908\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__14945\,
            I => \N__14903\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__14942\,
            I => \N__14903\
        );

    \I__1631\ : SRMux
    port map (
            O => \N__14941\,
            I => \N__14900\
        );

    \I__1630\ : InMux
    port map (
            O => \N__14940\,
            I => \N__14897\
        );

    \I__1629\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14894\
        );

    \I__1628\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14885\
        );

    \I__1627\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14885\
        );

    \I__1626\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14885\
        );

    \I__1625\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14885\
        );

    \I__1624\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14876\
        );

    \I__1623\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14876\
        );

    \I__1622\ : InMux
    port map (
            O => \N__14932\,
            I => \N__14876\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14931\,
            I => \N__14876\
        );

    \I__1620\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14871\
        );

    \I__1619\ : SRMux
    port map (
            O => \N__14929\,
            I => \N__14871\
        );

    \I__1618\ : InMux
    port map (
            O => \N__14928\,
            I => \N__14864\
        );

    \I__1617\ : InMux
    port map (
            O => \N__14927\,
            I => \N__14864\
        );

    \I__1616\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14864\
        );

    \I__1615\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14857\
        );

    \I__1614\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14857\
        );

    \I__1613\ : InMux
    port map (
            O => \N__14923\,
            I => \N__14857\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__14918\,
            I => \N__14854\
        );

    \I__1611\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14851\
        );

    \I__1610\ : SRMux
    port map (
            O => \N__14916\,
            I => \N__14841\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__14913\,
            I => \N__14836\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__14908\,
            I => \N__14836\
        );

    \I__1607\ : Span4Mux_h
    port map (
            O => \N__14903\,
            I => \N__14833\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__14900\,
            I => \N__14822\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__14897\,
            I => \N__14822\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__14894\,
            I => \N__14822\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__14885\,
            I => \N__14822\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__14876\,
            I => \N__14822\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__14871\,
            I => \N__14811\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__14864\,
            I => \N__14811\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__14857\,
            I => \N__14811\
        );

    \I__1598\ : Span4Mux_h
    port map (
            O => \N__14854\,
            I => \N__14811\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__14851\,
            I => \N__14811\
        );

    \I__1596\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14800\
        );

    \I__1595\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14800\
        );

    \I__1594\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14800\
        );

    \I__1593\ : InMux
    port map (
            O => \N__14847\,
            I => \N__14800\
        );

    \I__1592\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14800\
        );

    \I__1591\ : SRMux
    port map (
            O => \N__14845\,
            I => \N__14795\
        );

    \I__1590\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14795\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__14841\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__14836\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__14833\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__14822\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__14811\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__14800\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__14795\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__14780\,
            I => \PCH_PWRGD.N_2266_i_cascade_\
        );

    \I__1581\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14774\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__14774\,
            I => \PCH_PWRGD.curr_state_0_1\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__14771\,
            I => \PCH_PWRGD.m6_i_i_a2_cascade_\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__14768\,
            I => \PCH_PWRGD.count_rst_14_cascade_\
        );

    \I__1577\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14762\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14762\,
            I => \PCH_PWRGD.count_rst_7\
        );

    \I__1575\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14753\
        );

    \I__1574\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14753\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__14753\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__14750\,
            I => \N__14745\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__14749\,
            I => \N__14742\
        );

    \I__1570\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14739\
        );

    \I__1569\ : InMux
    port map (
            O => \N__14745\,
            I => \N__14735\
        );

    \I__1568\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14732\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__14739\,
            I => \N__14729\
        );

    \I__1566\ : InMux
    port map (
            O => \N__14738\,
            I => \N__14726\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__14735\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__14732\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__14729\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__14726\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1561\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14714\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__14714\,
            I => \PCH_PWRGD.count_1_i_a2_6_0\
        );

    \I__1559\ : InMux
    port map (
            O => \N__14711\,
            I => \N__14708\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__14705\,
            I => \PCH_PWRGD.count_1_i_a2_4_0\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \PCH_PWRGD.count_1_i_a2_5_0_cascade_\
        );

    \I__1555\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14696\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__14696\,
            I => \N__14693\
        );

    \I__1553\ : Span4Mux_h
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__14690\,
            I => \PCH_PWRGD.count_1_i_a2_3_0\
        );

    \I__1551\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14683\
        );

    \I__1550\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14680\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__14683\,
            I => \PCH_PWRGD.count_1_i_a2_12_0\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__14680\,
            I => \PCH_PWRGD.count_1_i_a2_12_0\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \N__14671\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__14674\,
            I => \N__14664\
        );

    \I__1545\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14661\
        );

    \I__1544\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14658\
        );

    \I__1543\ : InMux
    port map (
            O => \N__14669\,
            I => \N__14653\
        );

    \I__1542\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14653\
        );

    \I__1541\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14650\
        );

    \I__1540\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14647\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__14661\,
            I => \N__14640\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__14658\,
            I => \N__14640\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__14653\,
            I => \N__14640\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__14650\,
            I => \N__14637\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__14647\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__14640\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__14637\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__14630\,
            I => \PCH_PWRGD.count_1_i_a2_12_0_cascade_\
        );

    \I__1531\ : InMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__14624\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__1529\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__14615\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__14612\,
            I => \PCH_PWRGD.countZ0Z_15_cascade_\
        );

    \I__1525\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14606\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__14606\,
            I => \PCH_PWRGD.un2_count_1_axb_13\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__1522\ : InMux
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__14597\,
            I => \N__14593\
        );

    \I__1520\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14590\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__14593\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__14590\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1517\ : InMux
    port map (
            O => \N__14585\,
            I => \N__14581\
        );

    \I__1516\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14578\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__14581\,
            I => \N__14573\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__14578\,
            I => \N__14573\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__14573\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1512\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14567\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__14567\,
            I => \PCH_PWRGD.count_1_i_a2_1_0\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__14564\,
            I => \PCH_PWRGD.count_1_i_a2_0_0_cascade_\
        );

    \I__1509\ : InMux
    port map (
            O => \N__14561\,
            I => \N__14558\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__14558\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__14555\,
            I => \PCH_PWRGD.count_rst_9_cascade_\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__14552\,
            I => \N__14549\
        );

    \I__1505\ : InMux
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__14546\,
            I => \N__14543\
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__14543\,
            I => \PCH_PWRGD.un2_count_1_axb_10\
        );

    \I__1502\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14536\
        );

    \I__1501\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__14536\,
            I => \N__14530\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__14533\,
            I => \N__14527\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__14530\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__14527\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__14522\,
            I => \PCH_PWRGD.N_386_cascade_\
        );

    \I__1495\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__14516\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__14513\,
            I => \PCH_PWRGD.count_rst_3_cascade_\
        );

    \I__1492\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14504\
        );

    \I__1491\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14501\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__14508\,
            I => \N__14498\
        );

    \I__1489\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14495\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__14504\,
            I => \N__14490\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__14501\,
            I => \N__14490\
        );

    \I__1486\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14487\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__14495\,
            I => \N__14482\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__14490\,
            I => \N__14482\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__14487\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__14482\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__14477\,
            I => \PCH_PWRGD.count_rst_7_cascade_\
        );

    \I__1480\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14470\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14467\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__14470\,
            I => \PCH_PWRGD.un2_count_1_axb_7\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__14467\,
            I => \PCH_PWRGD.un2_count_1_axb_7\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__14462\,
            I => \N__14458\
        );

    \I__1475\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14455\
        );

    \I__1474\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14452\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__14455\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__14452\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__14447\,
            I => \PCH_PWRGD.un2_count_1_axb_7_cascade_\
        );

    \I__1470\ : InMux
    port map (
            O => \N__14444\,
            I => \N__14440\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14443\,
            I => \N__14437\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__14440\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__14437\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1466\ : InMux
    port map (
            O => \N__14432\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__1465\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14425\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14422\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__14425\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__14422\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1461\ : InMux
    port map (
            O => \N__14417\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__1460\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14410\
        );

    \I__1459\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14407\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__14410\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__14407\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1456\ : InMux
    port map (
            O => \N__14402\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__1455\ : InMux
    port map (
            O => \N__14399\,
            I => \bfn_2_3_0_\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__14396\,
            I => \N__14393\
        );

    \I__1453\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14389\
        );

    \I__1452\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14386\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__14386\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__14383\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1448\ : InMux
    port map (
            O => \N__14378\,
            I => \N__14375\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__14375\,
            I => \PCH_PWRGD.count_0_12\
        );

    \I__1446\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14366\
        );

    \I__1445\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14366\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__14366\,
            I => \N__14363\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__14363\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__1442\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14356\
        );

    \I__1441\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14353\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__14356\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__14353\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__1438\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14344\
        );

    \I__1437\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14341\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__14344\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__14341\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14336\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__1433\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14329\
        );

    \I__1432\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14326\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__14329\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__14326\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1429\ : InMux
    port map (
            O => \N__14321\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__14318\,
            I => \N__14315\
        );

    \I__1427\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14311\
        );

    \I__1426\ : InMux
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__14311\,
            I => \N__14305\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__14308\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__14305\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1422\ : InMux
    port map (
            O => \N__14300\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__1421\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14293\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14290\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__14293\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__14290\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1417\ : InMux
    port map (
            O => \N__14285\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__1416\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14278\
        );

    \I__1415\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14275\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__14278\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__14275\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1412\ : InMux
    port map (
            O => \N__14270\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__1411\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14263\
        );

    \I__1410\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14260\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__14263\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__14260\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1407\ : InMux
    port map (
            O => \N__14255\,
            I => \bfn_2_2_0_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14248\
        );

    \I__1405\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14245\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__14248\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__14245\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1402\ : InMux
    port map (
            O => \N__14240\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__1401\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14233\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14230\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__14233\,
            I => \N__14227\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__14230\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__14227\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1396\ : InMux
    port map (
            O => \N__14222\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__1395\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14215\
        );

    \I__1394\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14212\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__14215\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__14212\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14207\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__14204\,
            I => \POWERLED.N_660_cascade_\
        );

    \I__1389\ : InMux
    port map (
            O => \N__14201\,
            I => \N__14177\
        );

    \I__1388\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14177\
        );

    \I__1387\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14177\
        );

    \I__1386\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14168\
        );

    \I__1385\ : InMux
    port map (
            O => \N__14197\,
            I => \N__14168\
        );

    \I__1384\ : InMux
    port map (
            O => \N__14196\,
            I => \N__14168\
        );

    \I__1383\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14168\
        );

    \I__1382\ : InMux
    port map (
            O => \N__14194\,
            I => \N__14159\
        );

    \I__1381\ : InMux
    port map (
            O => \N__14193\,
            I => \N__14159\
        );

    \I__1380\ : InMux
    port map (
            O => \N__14192\,
            I => \N__14159\
        );

    \I__1379\ : InMux
    port map (
            O => \N__14191\,
            I => \N__14159\
        );

    \I__1378\ : InMux
    port map (
            O => \N__14190\,
            I => \N__14150\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14189\,
            I => \N__14150\
        );

    \I__1376\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14150\
        );

    \I__1375\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14150\
        );

    \I__1374\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14143\
        );

    \I__1373\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14143\
        );

    \I__1372\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14143\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__14177\,
            I => \N__14140\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__14168\,
            I => \N__14137\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__14159\,
            I => \N__14134\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__14150\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__14143\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__14140\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__14137\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1364\ : Odrv12
    port map (
            O => \N__14134\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1363\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14120\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__14120\,
            I => \POWERLED.pwm_out_1_sqmuxa_0\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__14117\,
            I => \POWERLED.pwm_out_en_cascade_\
        );

    \I__1360\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14110\
        );

    \I__1359\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14107\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__14110\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__14107\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__1356\ : IoInMux
    port map (
            O => \N__14102\,
            I => \N__14099\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__14099\,
            I => \N__14096\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__14096\,
            I => pwrbtn_led
        );

    \I__1353\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14090\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__1351\ : Span4Mux_s3_v
    port map (
            O => \N__14087\,
            I => \N__14084\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__14084\,
            I => vpp_ok
        );

    \I__1349\ : IoInMux
    port map (
            O => \N__14081\,
            I => \N__14078\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__14078\,
            I => \N__14075\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__14075\,
            I => vddq_en
        );

    \I__1346\ : InMux
    port map (
            O => \N__14072\,
            I => \N__14068\
        );

    \I__1345\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__14068\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__14065\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1342\ : InMux
    port map (
            O => \N__14060\,
            I => \N__14056\
        );

    \I__1341\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14053\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__14056\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__14053\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1338\ : InMux
    port map (
            O => \N__14048\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__14045\,
            I => \N__14041\
        );

    \I__1336\ : InMux
    port map (
            O => \N__14044\,
            I => \N__14038\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__14038\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__14035\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1332\ : InMux
    port map (
            O => \N__14030\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__1331\ : InMux
    port map (
            O => \N__14027\,
            I => \POWERLED.un1_count_cry_11\
        );

    \I__1330\ : InMux
    port map (
            O => \N__14024\,
            I => \POWERLED.un1_count_cry_12\
        );

    \I__1329\ : InMux
    port map (
            O => \N__14021\,
            I => \POWERLED.un1_count_cry_13\
        );

    \I__1328\ : InMux
    port map (
            O => \N__14018\,
            I => \POWERLED.un1_count_cry_14\
        );

    \I__1327\ : InMux
    port map (
            O => \N__14015\,
            I => \N__14011\
        );

    \I__1326\ : InMux
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__14011\,
            I => \N__14005\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__14008\,
            I => \POWERLED.count_1_12\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__14005\,
            I => \POWERLED.count_1_12\
        );

    \I__1322\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13997\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__1320\ : Odrv12
    port map (
            O => \N__13994\,
            I => \POWERLED.count_0_12\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__13991\,
            I => \POWERLED.N_437_cascade_\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \POWERLED.N_2305_i_cascade_\
        );

    \I__1317\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13979\
        );

    \I__1316\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13979\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__13979\,
            I => \N__13976\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__13976\,
            I => \POWERLED.count_1_3\
        );

    \I__1313\ : InMux
    port map (
            O => \N__13973\,
            I => \POWERLED.un1_count_cry_2_cZ0\
        );

    \I__1312\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13964\
        );

    \I__1311\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13964\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__13964\,
            I => \POWERLED.count_1_4\
        );

    \I__1309\ : InMux
    port map (
            O => \N__13961\,
            I => \POWERLED.un1_count_cry_3_cZ0\
        );

    \I__1308\ : InMux
    port map (
            O => \N__13958\,
            I => \POWERLED.un1_count_cry_4_cZ0\
        );

    \I__1307\ : InMux
    port map (
            O => \N__13955\,
            I => \POWERLED.un1_count_cry_5\
        );

    \I__1306\ : InMux
    port map (
            O => \N__13952\,
            I => \POWERLED.un1_count_cry_6\
        );

    \I__1305\ : InMux
    port map (
            O => \N__13949\,
            I => \POWERLED.un1_count_cry_7\
        );

    \I__1304\ : InMux
    port map (
            O => \N__13946\,
            I => \bfn_1_12_0_\
        );

    \I__1303\ : InMux
    port map (
            O => \N__13943\,
            I => \POWERLED.un1_count_cry_9\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__13940\,
            I => \N__13937\
        );

    \I__1301\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13931\
        );

    \I__1300\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13931\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__13928\,
            I => \POWERLED.count_1_11\
        );

    \I__1297\ : InMux
    port map (
            O => \N__13925\,
            I => \POWERLED.un1_count_cry_10\
        );

    \I__1296\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__13919\,
            I => \POWERLED.count_0_0\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__13916\,
            I => \POWERLED.count_1_0_cascade_\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__13913\,
            I => \POWERLED.countZ0Z_0_cascade_\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__13910\,
            I => \POWERLED.count_1_1_cascade_\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__13907\,
            I => \POWERLED.countZ0Z_1_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__13901\,
            I => \POWERLED.count_0_1\
        );

    \I__1288\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__13895\,
            I => \POWERLED.count_0_4\
        );

    \I__1286\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13886\
        );

    \I__1285\ : InMux
    port map (
            O => \N__13891\,
            I => \N__13886\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__13883\,
            I => \POWERLED.count_1_2\
        );

    \I__1282\ : InMux
    port map (
            O => \N__13880\,
            I => \POWERLED.un1_count_cry_1\
        );

    \I__1281\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__13874\,
            I => \POWERLED.count_0_2\
        );

    \I__1279\ : IoInMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__13868\,
            I => \G_12\
        );

    \I__1277\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__13862\,
            I => \POWERLED.count_0_11\
        );

    \I__1275\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__13856\,
            I => \POWERLED.count_0_3\
        );

    \I__1273\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13850\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__13850\,
            I => \PCH_PWRGD.count_0_6\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__13847\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_\
        );

    \I__1270\ : InMux
    port map (
            O => \N__13844\,
            I => \N__13838\
        );

    \I__1269\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13838\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__13838\,
            I => \N__13835\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__13835\,
            I => \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__13832\,
            I => \PCH_PWRGD.un2_count_1_axb_1_cascade_\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__13829\,
            I => \PCH_PWRGD.N_2284_i_cascade_\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__13826\,
            I => \PCH_PWRGD.N_655_cascade_\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__13823\,
            I => \PCH_PWRGD.count_0_sqmuxa_cascade_\
        );

    \I__1262\ : InMux
    port map (
            O => \N__13820\,
            I => \N__13816\
        );

    \I__1261\ : InMux
    port map (
            O => \N__13819\,
            I => \N__13813\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__13816\,
            I => \N__13810\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__13813\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__13810\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__1257\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13799\
        );

    \I__1256\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13799\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__13799\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__13796\,
            I => \N__13793\
        );

    \I__1253\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13787\
        );

    \I__1252\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13787\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__13787\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__1250\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13780\
        );

    \I__1249\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13777\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__13780\,
            I => vr_ready_vccin
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__13777\,
            I => vr_ready_vccin
        );

    \I__1246\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13769\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__13769\,
            I => \PCH_PWRGD.N_2284_i\
        );

    \I__1244\ : InMux
    port map (
            O => \N__13766\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__1243\ : InMux
    port map (
            O => \N__13763\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__1242\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13757\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__13757\,
            I => \N__13754\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__13754\,
            I => \PCH_PWRGD.un2_count_1_axb_2\
        );

    \I__1239\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13744\
        );

    \I__1238\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13744\
        );

    \I__1237\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13741\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13738\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__13741\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__13738\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__1233\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13729\
        );

    \I__1232\ : InMux
    port map (
            O => \N__13732\,
            I => \N__13726\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__13729\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__13726\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__1229\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13718\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__13718\,
            I => \PCH_PWRGD.count_0_14\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__13715\,
            I => \N__13711\
        );

    \I__1226\ : InMux
    port map (
            O => \N__13714\,
            I => \N__13706\
        );

    \I__1225\ : InMux
    port map (
            O => \N__13711\,
            I => \N__13706\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__13706\,
            I => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\
        );

    \I__1223\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13697\
        );

    \I__1222\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13697\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__13697\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__1220\ : InMux
    port map (
            O => \N__13694\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__1219\ : InMux
    port map (
            O => \N__13691\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__1218\ : InMux
    port map (
            O => \N__13688\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__1217\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13680\
        );

    \I__1216\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13677\
        );

    \I__1215\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13674\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__13680\,
            I => \N__13671\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__13677\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__13674\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__13671\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__13664\,
            I => \N__13660\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__13663\,
            I => \N__13657\
        );

    \I__1208\ : InMux
    port map (
            O => \N__13660\,
            I => \N__13654\
        );

    \I__1207\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13651\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__13654\,
            I => \N__13646\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__13651\,
            I => \N__13646\
        );

    \I__1204\ : Span4Mux_s2_v
    port map (
            O => \N__13646\,
            I => \N__13643\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__13643\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1202\ : InMux
    port map (
            O => \N__13640\,
            I => \PCH_PWRGD.un2_count_1_cry_7\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__13637\,
            I => \N__13634\
        );

    \I__1200\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13630\
        );

    \I__1199\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13627\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__13630\,
            I => \N__13624\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__13627\,
            I => \N__13621\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__13624\,
            I => \PCH_PWRGD.un2_count_1_axb_9\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__13621\,
            I => \PCH_PWRGD.un2_count_1_axb_9\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13610\
        );

    \I__1193\ : InMux
    port map (
            O => \N__13615\,
            I => \N__13610\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__13610\,
            I => \N__13607\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__13607\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1190\ : InMux
    port map (
            O => \N__13604\,
            I => \bfn_1_6_0_\
        );

    \I__1189\ : InMux
    port map (
            O => \N__13601\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__1188\ : InMux
    port map (
            O => \N__13598\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__1187\ : InMux
    port map (
            O => \N__13595\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__1186\ : InMux
    port map (
            O => \N__13592\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__13589\,
            I => \PCH_PWRGD.un2_count_1_axb_4_cascade_\
        );

    \I__1184\ : InMux
    port map (
            O => \N__13586\,
            I => \N__13583\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__13583\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__1182\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13577\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__13577\,
            I => \PCH_PWRGD.count_rst_10\
        );

    \I__1180\ : InMux
    port map (
            O => \N__13574\,
            I => \N__13568\
        );

    \I__1179\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13568\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__13568\,
            I => \N__13565\
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__13565\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__13562\,
            I => \PCH_PWRGD.count_rst_10_cascade_\
        );

    \I__1175\ : InMux
    port map (
            O => \N__13559\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \I__1174\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13548\
        );

    \I__1173\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13548\
        );

    \I__1172\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13545\
        );

    \I__1171\ : InMux
    port map (
            O => \N__13553\,
            I => \N__13542\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__13548\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__13545\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__13542\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__13535\,
            I => \N__13531\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__13534\,
            I => \N__13528\
        );

    \I__1165\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13523\
        );

    \I__1164\ : InMux
    port map (
            O => \N__13528\,
            I => \N__13523\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__13523\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__1162\ : InMux
    port map (
            O => \N__13520\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__1161\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13513\
        );

    \I__1160\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13510\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__13513\,
            I => \PCH_PWRGD.un2_count_1_axb_4\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__13510\,
            I => \PCH_PWRGD.un2_count_1_axb_4\
        );

    \I__1157\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13499\
        );

    \I__1156\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13499\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__13499\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__1154\ : InMux
    port map (
            O => \N__13496\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__13493\,
            I => \PCH_PWRGD.count_rst_5_cascade_\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \PCH_PWRGD.un2_count_1_axb_9_cascade_\
        );

    \I__1151\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__13484\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__13481\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__1148\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13472\
        );

    \I__1147\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13472\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__13472\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__13469\,
            I => \PCH_PWRGD.countZ0Z_8_cascade_\
        );

    \I__1144\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__13463\,
            I => \PCH_PWRGD.count_rst_5\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__13460\,
            I => \PCH_PWRGD.count_rst_11_cascade_\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__13457\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10_cascade_\
        );

    \I__1140\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__13451\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__13448\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__13442\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12\
        );

    \I__1135\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__13436\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un3_count_off_1_cry_8\,
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_6_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_16_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_15_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_cry_8\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_5_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_1_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_7\,
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_15\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_2_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_1_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_7_15_0_\
        );

    \N_92_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__13871\,
            GLOBALBUFFEROUTPUT => \N_92_g\
        );

    \N_557_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32674\,
            GLOBALBUFFEROUTPUT => \N_557_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI4MLK1_1_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14251\,
            in1 => \N__14332\,
            in2 => \N__14045\,
            in3 => \N__14059\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIST215_10_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13454\,
            in1 => \N__13439\,
            in2 => \N__13457\,
            in3 => \N__13445\,
            lcout => \N_662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIMVQE1_3_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21173\,
            in1 => \N__14347\,
            in2 => \N__14318\,
            in3 => \N__14296\,
            lcout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIVSS4_11_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14443\,
            in2 => \_gnd_net_\,
            in3 => \N__14218\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI6CM11_10_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14237\,
            in1 => \N__14266\,
            in2 => \N__13448\,
            in3 => \N__14281\,
            lcout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14428\,
            in1 => \N__14413\,
            in2 => \N__14396\,
            in3 => \N__14071\,
            lcout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_8_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__15351\,
            in1 => \N__14940\,
            in2 => \N__13664\,
            in3 => \N__13683\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32317\,
            ce => \N__15138\,
            sr => \N__14941\
        );

    \PCH_PWRGD.count_11_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__14937\,
            in1 => \N__15355\,
            in2 => \N__14508\,
            in3 => \N__14539\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32355\,
            ce => \N__15132\,
            sr => \N__14965\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__14936\,
            in1 => \N__13615\,
            in2 => \N__13637\,
            in3 => \N__15354\,
            lcout => \PCH_PWRGD.count_rst_5\,
            ltout => \PCH_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI27DA2_9_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15068\,
            in1 => \_gnd_net_\,
            in2 => \N__13493\,
            in3 => \N__13477\,
            lcout => \PCH_PWRGD.un2_count_1_axb_9\,
            ltout => \PCH_PWRGD.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_9_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__14938\,
            in1 => \N__15356\,
            in2 => \N__13490\,
            in3 => \N__13616\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32355\,
            ce => \N__15132\,
            sr => \N__14965\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__15353\,
            in1 => \N__14935\,
            in2 => \N__13663\,
            in3 => \N__13684\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQOP84_8_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13487\,
            in2 => \N__13481\,
            in3 => \N__15067\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => \PCH_PWRGD.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI27DA2_0_9_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__15069\,
            in1 => \N__13478\,
            in2 => \N__13469\,
            in3 => \N__13466\,
            lcout => \PCH_PWRGD.count_1_i_a2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__13556\,
            in1 => \N__15319\,
            in2 => \N__13534\,
            in3 => \N__14931\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15064\,
            in1 => \_gnd_net_\,
            in2 => \N__13460\,
            in3 => \N__13586\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIT1DA2_4_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13573\,
            in1 => \N__15065\,
            in2 => \_gnd_net_\,
            in3 => \N__13580\,
            lcout => \PCH_PWRGD.un2_count_1_axb_4\,
            ltout => \PCH_PWRGD.un2_count_1_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__15324\,
            in1 => \N__14960\,
            in2 => \N__13589\,
            in3 => \N__13505\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32335\,
            ce => \N__15070\,
            sr => \N__14966\
        );

    \PCH_PWRGD.count_3_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__13555\,
            in1 => \N__15323\,
            in2 => \N__13535\,
            in3 => \N__14934\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32335\,
            ce => \N__15070\,
            sr => \N__14966\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__14932\,
            in1 => \N__13517\,
            in2 => \N__15349\,
            in3 => \N__13504\,
            lcout => \PCH_PWRGD.count_rst_10\,
            ltout => \PCH_PWRGD.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIT1DA2_0_4_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__13574\,
            in1 => \N__15066\,
            in2 => \N__13562\,
            in3 => \N__13554\,
            lcout => \PCH_PWRGD.count_1_i_a2_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_5_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__14933\,
            in1 => \N__14748\,
            in2 => \N__15350\,
            in3 => \N__14360\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32335\,
            ce => \N__15070\,
            sr => \N__14966\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13820\,
            in2 => \N__14674\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14917\,
            in1 => \N__13760\,
            in2 => \_gnd_net_\,
            in3 => \N__13559\,
            lcout => \PCH_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13553\,
            in2 => \_gnd_net_\,
            in3 => \N__13520\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13516\,
            in2 => \_gnd_net_\,
            in3 => \N__13496\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14738\,
            in2 => \_gnd_net_\,
            in3 => \N__13694\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14603\,
            in3 => \N__13691\,
            lcout => \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14473\,
            in2 => \_gnd_net_\,
            in3 => \N__13688\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13685\,
            in2 => \_gnd_net_\,
            in3 => \N__13640\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13633\,
            in2 => \_gnd_net_\,
            in3 => \N__13604\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__14926\,
            in1 => \_gnd_net_\,
            in2 => \N__14552\,
            in3 => \N__13601\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14510\,
            in2 => \_gnd_net_\,
            in3 => \N__13598\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14927\,
            in1 => \N__14584\,
            in2 => \_gnd_net_\,
            in3 => \N__13595\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNI523P1_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14939\,
            in1 => \N__14609\,
            in2 => \_gnd_net_\,
            in3 => \N__13592\,
            lcout => \PCH_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13702\,
            in2 => \_gnd_net_\,
            in3 => \N__13766\,
            lcout => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__14621\,
            in1 => \N__14928\,
            in2 => \_gnd_net_\,
            in3 => \N__13763\,
            lcout => \PCH_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIE6J84_0_2_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010011"
        )
    port map (
            in0 => \N__13749\,
            in1 => \N__13733\,
            in2 => \N__15098\,
            in3 => \N__13703\,
            lcout => \PCH_PWRGD.count_1_i_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_6_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__13843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14849\,
            lcout => \PCH_PWRGD.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32401\,
            ce => \N__15140\,
            sr => \N__14916\
        );

    \PCH_PWRGD.count_RNIE6J84_2_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13732\,
            in1 => \N__15017\,
            in2 => \_gnd_net_\,
            in3 => \N__13750\,
            lcout => \PCH_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_2_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13751\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32401\,
            ce => \N__15140\,
            sr => \N__14916\
        );

    \PCH_PWRGD.count_14_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__14848\,
            in1 => \N__13714\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32401\,
            ce => \N__15140\,
            sr => \N__14916\
        );

    \PCH_PWRGD.count_RNIKP0C4_14_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__15018\,
            in1 => \N__13721\,
            in2 => \N__13715\,
            in3 => \N__14847\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNISDK72_0_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000000"
        )
    port map (
            in0 => \N__15407\,
            in1 => \N__14846\,
            in2 => \N__15862\,
            in3 => \N__32675\,
            lcout => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\,
            ltout => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIMIN84_6_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__14850\,
            in1 => \N__13853\,
            in2 => \N__13847\,
            in3 => \N__13844\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQUCA2_1_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13792\,
            in1 => \N__15016\,
            in2 => \_gnd_net_\,
            in3 => \N__13805\,
            lcout => \PCH_PWRGD.un2_count_1_axb_1\,
            ltout => \PCH_PWRGD.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIRP9H1_1_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14668\,
            in2 => \N__13832\,
            in3 => \N__14844\,
            lcout => \PCH_PWRGD.count_rst_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15379\,
            lcout => \PCH_PWRGD.N_2284_i\,
            ltout => \PCH_PWRGD.N_2284_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIDKSB1_0_1_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13783\,
            in2 => \N__13829\,
            in3 => \N__29609\,
            lcout => \PCH_PWRGD.N_655\,
            ltout => \PCH_PWRGD.N_655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15835\,
            in2 => \N__13826\,
            in3 => \N__25739\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => \PCH_PWRGD.count_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_1_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14669\,
            in2 => \N__13823\,
            in3 => \N__13819\,
            lcout => \PCH_PWRGD.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32431\,
            ce => \N__15071\,
            sr => \N__14845\
        );

    \PCH_PWRGD.count_RNIQUCA2_0_1_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__15072\,
            in1 => \N__13804\,
            in2 => \N__13796\,
            in3 => \N__14509\,
            lcout => \PCH_PWRGD.count_1_i_a2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__13784\,
            in1 => \N__13772\,
            in2 => \_gnd_net_\,
            in3 => \N__29610\,
            lcout => \PCH_PWRGD.N_670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIAKSS_2_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25734\,
            in1 => \N__13877\,
            in2 => \_gnd_net_\,
            in3 => \N__13891\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32436\,
            ce => \N__16464\,
            sr => \_gnd_net_\
        );

    \POWERLED.G_12_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25738\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22549\,
            lcout => \G_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIALHT_11_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13865\,
            in1 => \N__25736\,
            in2 => \_gnd_net_\,
            in3 => \N__13936\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_11_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13940\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32436\,
            ce => \N__16464\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICNTS_3_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13859\,
            in1 => \N__25735\,
            in2 => \_gnd_net_\,
            in3 => \N__13984\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_3_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13985\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32436\,
            ce => \N__16464\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICOIT_12_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14000\,
            in1 => \N__25737\,
            in2 => \_gnd_net_\,
            in3 => \N__14015\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIEQUS_4_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25747\,
            in1 => \N__13898\,
            in2 => \_gnd_net_\,
            in3 => \N__13969\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17252\,
            lcout => \POWERLED.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32460\,
            ce => \N__16463\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIE5D5_0_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14191\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNITFSJ_0_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13922\,
            in2 => \N__13916\,
            in3 => \N__25745\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => \POWERLED.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIE5D5_1_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__17214\,
            in1 => \_gnd_net_\,
            in2 => \N__13913\,
            in3 => \N__14192\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUGSJ_1_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13904\,
            in2 => \N__13910\,
            in3 => \N__25746\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => \POWERLED.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__17253\,
            in1 => \_gnd_net_\,
            in2 => \N__13907\,
            in3 => \N__14194\,
            lcout => \POWERLED.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32460\,
            ce => \N__16463\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_4_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13970\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32460\,
            ce => \N__16463\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17251\,
            in2 => \N__17218\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \POWERLED.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14195\,
            in1 => \_gnd_net_\,
            in2 => \N__17179\,
            in3 => \N__13880\,
            lcout => \POWERLED.count_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_1\,
            carryout => \POWERLED.un1_count_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_2_c_RNIQ9EE_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14199\,
            in1 => \_gnd_net_\,
            in2 => \N__17140\,
            in3 => \N__13973\,
            lcout => \POWERLED.count_1_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_2_cZ0\,
            carryout => \POWERLED.un1_count_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_3_c_RNIRBFE_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14196\,
            in1 => \_gnd_net_\,
            in2 => \N__17098\,
            in3 => \N__13961\,
            lcout => \POWERLED.count_1_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_3_cZ0\,
            carryout => \POWERLED.un1_count_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNISDGE_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14200\,
            in1 => \_gnd_net_\,
            in2 => \N__17058\,
            in3 => \N__13958\,
            lcout => \POWERLED.count_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_4_cZ0\,
            carryout => \POWERLED.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNITFHE_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14197\,
            in1 => \_gnd_net_\,
            in2 => \N__17019\,
            in3 => \N__13955\,
            lcout => \POWERLED.count_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_5\,
            carryout => \POWERLED.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__14201\,
            in1 => \N__16974\,
            in2 => \_gnd_net_\,
            in3 => \N__13952\,
            lcout => \POWERLED.count_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_6\,
            carryout => \POWERLED.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14198\,
            in1 => \_gnd_net_\,
            in2 => \N__17530\,
            in3 => \N__13949\,
            lcout => \POWERLED.count_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_7\,
            carryout => \POWERLED.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14184\,
            in1 => \_gnd_net_\,
            in2 => \N__17497\,
            in3 => \N__13946\,
            lcout => \POWERLED.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \POWERLED.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14187\,
            in1 => \_gnd_net_\,
            in2 => \N__17464\,
            in3 => \N__13943\,
            lcout => \POWERLED.count_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_9\,
            carryout => \POWERLED.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14185\,
            in1 => \_gnd_net_\,
            in2 => \N__17410\,
            in3 => \N__13925\,
            lcout => \POWERLED.count_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_10\,
            carryout => \POWERLED.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14188\,
            in1 => \_gnd_net_\,
            in2 => \N__17371\,
            in3 => \N__14027\,
            lcout => \POWERLED.count_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_11\,
            carryout => \POWERLED.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14186\,
            in1 => \_gnd_net_\,
            in2 => \N__17328\,
            in3 => \N__14024\,
            lcout => \POWERLED.count_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_12\,
            carryout => \POWERLED.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_13_c_RNICO0D_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__14189\,
            in1 => \_gnd_net_\,
            in2 => \N__17292\,
            in3 => \N__14021\,
            lcout => \POWERLED.count_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_13\,
            carryout => \POWERLED.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__17640\,
            in1 => \N__14190\,
            in2 => \_gnd_net_\,
            in3 => \N__14018\,
            lcout => \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_12_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14014\,
            lcout => \POWERLED.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32469\,
            ce => \N__16469\,
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIE5D5_0_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__16565\,
            in1 => \_gnd_net_\,
            in2 => \N__25744\,
            in3 => \N__15557\,
            lcout => \POWERLED.pwm_out_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011000000"
        )
    port map (
            in0 => \N__17608\,
            in1 => \N__14113\,
            in2 => \N__15530\,
            in3 => \N__16564\,
            lcout => \POWERLED.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32470\,
            ce => 'H',
            sr => \N__15587\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__16566\,
            in1 => \N__16525\,
            in2 => \_gnd_net_\,
            in3 => \N__17607\,
            lcout => OPEN,
            ltout => \POWERLED.N_437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNICO541_0_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16511\,
            in2 => \N__13991\,
            in3 => \N__25697\,
            lcout => \POWERLED.N_2305_i\,
            ltout => \POWERLED.N_2305_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI_0_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__15553\,
            in1 => \_gnd_net_\,
            in2 => \N__13988\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_660\,
            ltout => \POWERLED.N_660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIE5D5_0_0_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14204\,
            in3 => \N__25698\,
            lcout => \POWERLED.count_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNIPOMA1_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__17609\,
            in1 => \N__14123\,
            in2 => \N__16499\,
            in3 => \N__16568\,
            lcout => OPEN,
            ltout => \POWERLED.pwm_out_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNIKIDQ1_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16567\,
            in1 => \_gnd_net_\,
            in2 => \N__14117\,
            in3 => \N__14114\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__33131\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14093\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25426\,
            in1 => \N__14072\,
            in2 => \N__16142\,
            in3 => \N__16141\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_1_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25411\,
            in1 => \N__14060\,
            in2 => \_gnd_net_\,
            in3 => \N__14048\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25427\,
            in1 => \N__14044\,
            in2 => \_gnd_net_\,
            in3 => \N__14030\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_3_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25412\,
            in1 => \N__14348\,
            in2 => \_gnd_net_\,
            in3 => \N__14336\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_4_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25428\,
            in1 => \N__14333\,
            in2 => \_gnd_net_\,
            in3 => \N__14321\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25413\,
            in1 => \N__14314\,
            in2 => \_gnd_net_\,
            in3 => \N__14300\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_6_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25429\,
            in1 => \N__14297\,
            in2 => \_gnd_net_\,
            in3 => \N__14285\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25414\,
            in1 => \N__14282\,
            in2 => \_gnd_net_\,
            in3 => \N__14270\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__32235\,
            ce => 'H',
            sr => \N__20960\
        );

    \RSMRST_PWRGD.count_8_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25425\,
            in1 => \N__14267\,
            in2 => \_gnd_net_\,
            in3 => \N__14255\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__32316\,
            ce => 'H',
            sr => \N__20955\
        );

    \RSMRST_PWRGD.count_9_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25410\,
            in1 => \N__14252\,
            in2 => \_gnd_net_\,
            in3 => \N__14240\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__32316\,
            ce => 'H',
            sr => \N__20955\
        );

    \RSMRST_PWRGD.count_10_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25422\,
            in1 => \N__14236\,
            in2 => \_gnd_net_\,
            in3 => \N__14222\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__32316\,
            ce => 'H',
            sr => \N__20955\
        );

    \RSMRST_PWRGD.count_11_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25408\,
            in1 => \N__14219\,
            in2 => \_gnd_net_\,
            in3 => \N__14207\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__32316\,
            ce => 'H',
            sr => \N__20955\
        );

    \RSMRST_PWRGD.count_12_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25423\,
            in1 => \N__14444\,
            in2 => \_gnd_net_\,
            in3 => \N__14432\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__32316\,
            ce => 'H',
            sr => \N__20955\
        );

    \RSMRST_PWRGD.count_13_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25409\,
            in1 => \N__14429\,
            in2 => \_gnd_net_\,
            in3 => \N__14417\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__32316\,
            ce => 'H',
            sr => \N__20955\
        );

    \RSMRST_PWRGD.count_14_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25424\,
            in1 => \N__14414\,
            in2 => \_gnd_net_\,
            in3 => \N__14402\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__32316\,
            ce => 'H',
            sr => \N__20955\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25193\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14392\,
            in2 => \_gnd_net_\,
            in3 => \N__14399\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32354\,
            ce => \N__17732\,
            sr => \N__20959\
        );

    \PCH_PWRGD.count_12_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14372\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32318\,
            ce => \N__15139\,
            sr => \N__14959\
        );

    \PCH_PWRGD.count_RNIGJUB4_12_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14378\,
            in1 => \N__15101\,
            in2 => \_gnd_net_\,
            in3 => \N__14371\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__14359\,
            in1 => \N__15328\,
            in2 => \N__14750\,
            in3 => \N__14957\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIKFM84_5_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14561\,
            in2 => \N__14555\,
            in3 => \N__15099\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15100\,
            in1 => \N__15155\,
            in2 => \_gnd_net_\,
            in3 => \N__15178\,
            lcout => \PCH_PWRGD.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIPCK99_0_1_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__14667\,
            in1 => \N__14686\,
            in2 => \_gnd_net_\,
            in3 => \N__15233\,
            lcout => \PCH_PWRGD.N_386\,
            ltout => \PCH_PWRGD.N_386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__14540\,
            in1 => \N__14507\,
            in2 => \N__14522\,
            in3 => \N__14958\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIEGTB4_11_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__14519\,
            in1 => \_gnd_net_\,
            in2 => \N__14513\,
            in3 => \N__15102\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__15329\,
            in1 => \N__14474\,
            in2 => \N__14462\,
            in3 => \N__14923\,
            lcout => \PCH_PWRGD.count_rst_7\,
            ltout => \PCH_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI05DA2_7_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14758\,
            in2 => \N__14477\,
            in3 => \N__15088\,
            lcout => \PCH_PWRGD.un2_count_1_axb_7\,
            ltout => \PCH_PWRGD.un2_count_1_axb_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_7_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__15330\,
            in1 => \N__14461\,
            in2 => \N__14447\,
            in3 => \N__14925\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32356\,
            ce => \N__15136\,
            sr => \N__14929\
        );

    \PCH_PWRGD.count_RNIK6UQA_1_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__14687\,
            in1 => \N__14930\,
            in2 => \N__14675\,
            in3 => \N__15228\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNID4B5D_0_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15137\,
            in1 => \_gnd_net_\,
            in2 => \N__14768\,
            in3 => \N__14627\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI05DA2_0_7_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__14765\,
            in1 => \N__14759\,
            in2 => \N__14749\,
            in3 => \N__15089\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIPCK99_1_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14717\,
            in1 => \N__14711\,
            in2 => \N__14702\,
            in3 => \N__14699\,
            lcout => \PCH_PWRGD.count_1_i_a2_12_0\,
            ltout => \PCH_PWRGD.count_1_i_a2_12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__14924\,
            in1 => \N__14670\,
            in2 => \N__14630\,
            in3 => \N__15229\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32356\,
            ce => \N__15136\,
            sr => \N__14929\
        );

    \PCH_PWRGD.count_RNIMS1C4_15_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15215\,
            in1 => \N__15206\,
            in2 => \_gnd_net_\,
            in3 => \N__15055\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => \PCH_PWRGD.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIIMVB4_0_13_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__15200\,
            in1 => \N__15188\,
            in2 => \N__14612\,
            in3 => \N__15131\,
            lcout => \PCH_PWRGD.count_1_i_a2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIIMVB4_13_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15187\,
            in1 => \N__15053\,
            in2 => \_gnd_net_\,
            in3 => \N__15198\,
            lcout => \PCH_PWRGD.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI58BH4_0_10_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000010011"
        )
    port map (
            in0 => \N__15054\,
            in1 => \N__14596\,
            in2 => \N__15179\,
            in3 => \N__15151\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI55U5D_2_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14585\,
            in1 => \N__14570\,
            in2 => \N__14564\,
            in3 => \N__15239\,
            lcout => \PCH_PWRGD.count_1_i_a2_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_15_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15214\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32411\,
            ce => \N__15130\,
            sr => \N__14961\
        );

    \PCH_PWRGD.count_13_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15199\,
            lcout => \PCH_PWRGD.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32411\,
            ce => \N__15130\,
            sr => \N__14961\
        );

    \PCH_PWRGD.count_10_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15174\,
            lcout => \PCH_PWRGD.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32411\,
            ce => \N__15130\,
            sr => \N__14961\
        );

    \PCH_PWRGD.curr_state_1_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__15840\,
            in1 => \N__15391\,
            in2 => \N__15352\,
            in3 => \N__15375\,
            lcout => \PCH_PWRGD.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32402\,
            ce => \N__16462\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15406\,
            lcout => \PCH_PWRGD.N_2266_i\,
            ltout => \PCH_PWRGD.N_2266_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__15335\,
            in1 => \N__15798\,
            in2 => \N__14780\,
            in3 => \N__15373\,
            lcout => \PCH_PWRGD.curr_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__15392\,
            in1 => \N__15334\,
            in2 => \N__15380\,
            in3 => \N__15841\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.m6_i_i_a2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIC58V1_1_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14777\,
            in2 => \N__14771\,
            in3 => \N__25732\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25733\,
            in1 => \N__15266\,
            in2 => \_gnd_net_\,
            in3 => \N__15413\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15395\,
            in3 => \N__15390\,
            lcout => \PCH_PWRGD.curr_state_0_sqmuxa\,
            ltout => \PCH_PWRGD.curr_state_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__15374\,
            in1 => \N__15336\,
            in2 => \N__15269\,
            in3 => \N__15839\,
            lcout => \PCH_PWRGD.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32402\,
            ce => \N__16462\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__16369\,
            in1 => \N__16329\,
            in2 => \N__22334\,
            in3 => \N__16046\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32430\,
            ce => \N__16465\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__16401\,
            in1 => \N__16108\,
            in2 => \N__16083\,
            in3 => \N__16367\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__25741\,
            in1 => \_gnd_net_\,
            in2 => \N__15260\,
            in3 => \N__15254\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__16400\,
            in1 => \N__16109\,
            in2 => \N__15257\,
            in3 => \N__16370\,
            lcout => \VPP_VDDQ.curr_state_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32430\,
            ce => \N__16465\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__22330\,
            in1 => \N__16330\,
            in2 => \N__16380\,
            in3 => \N__16045\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.m4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15248\,
            in2 => \N__15242\,
            in3 => \N__25740\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__25742\,
            in1 => \_gnd_net_\,
            in2 => \N__15518\,
            in3 => \N__16402\,
            lcout => \VPP_VDDQ.N_60\,
            ltout => \VPP_VDDQ.N_60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNINI731_0_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__16493\,
            in1 => \N__16368\,
            in2 => \N__15515\,
            in3 => \N__22331\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNO_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15498\,
            lcout => \VPP_VDDQ.N_60_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__15472\,
            in1 => \N__22323\,
            in2 => \N__15485\,
            in3 => \N__15499\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32435\,
            ce => 'H',
            sr => \N__15512\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__15500\,
            in1 => \N__15484\,
            in2 => \N__22333\,
            in3 => \N__15473\,
            lcout => OPEN,
            ltout => \VPP_VDDQ_delayed_vddq_ok_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_PWRGD_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__15983\,
            in1 => \_gnd_net_\,
            in2 => \N__15464\,
            in3 => \_gnd_net_\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16073\,
            lcout => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_a2_0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15443\,
            in3 => \N__22322\,
            lcout => \N_639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15982\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI1Q9V_10_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15692\,
            in1 => \N__25743\,
            in2 => \_gnd_net_\,
            in3 => \N__15707\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25756\,
            in1 => \N__16570\,
            in2 => \_gnd_net_\,
            in3 => \N__15552\,
            lcout => \POWERLED.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_2_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17169\,
            in1 => \N__17094\,
            in2 => \_gnd_net_\,
            in3 => \N__17130\,
            lcout => \POWERLED.un79_clk_100khzlt6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_7_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17493\,
            in1 => \N__17526\,
            in2 => \_gnd_net_\,
            in3 => \N__16975\,
            lcout => \POWERLED.un79_clk_100khzlto15_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_15_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17364\,
            in1 => \N__17329\,
            in2 => \N__17644\,
            in3 => \N__17293\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_5_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__15575\,
            in1 => \N__17020\,
            in2 => \N__15569\,
            in3 => \N__17059\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_10_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15566\,
            in1 => \N__17454\,
            in2 => \N__15560\,
            in3 => \N__17403\,
            lcout => \POWERLED.un79_clk_100khz\,
            ltout => \POWERLED.un79_clk_100khz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101111111"
        )
    port map (
            in0 => \N__25757\,
            in1 => \N__16494\,
            in2 => \N__15533\,
            in3 => \N__16569\,
            lcout => \POWERLED.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNII1MT_15_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15656\,
            in1 => \N__25755\,
            in2 => \_gnd_net_\,
            in3 => \N__15664\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_15_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15668\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32459\,
            ce => \N__16466\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIK32T_7_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15641\,
            in1 => \N__25752\,
            in2 => \_gnd_net_\,
            in3 => \N__15649\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_7_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32459\,
            ce => \N__16466\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIM63T_8_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15626\,
            in1 => \N__25753\,
            in2 => \_gnd_net_\,
            in3 => \N__15634\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_8_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32459\,
            ce => \N__16466\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIO94T_9_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15611\,
            in1 => \N__25754\,
            in2 => \_gnd_net_\,
            in3 => \N__15619\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_9_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32459\,
            ce => \N__16466\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIERJT_13_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15593\,
            in1 => \N__25750\,
            in2 => \_gnd_net_\,
            in3 => \N__15601\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_13_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15605\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32468\,
            ce => \N__16468\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGTVS_5_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15746\,
            in1 => \N__25748\,
            in2 => \_gnd_net_\,
            in3 => \N__15754\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_5_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15755\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32468\,
            ce => \N__16468\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGUKT_14_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15728\,
            in1 => \N__25751\,
            in2 => \_gnd_net_\,
            in3 => \N__15736\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_14_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15740\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32468\,
            ce => \N__16468\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNII01T_6_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15713\,
            in1 => \N__25749\,
            in2 => \_gnd_net_\,
            in3 => \N__15721\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_6_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32468\,
            ce => \N__16468\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18512\,
            lcout => \POWERLED.mult1_un96_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_10_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15706\,
            lcout => \POWERLED.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32467\,
            ce => \N__16467\,
            sr => \_gnd_net_\
        );

    \SLP_SUSn_RNIN4K9_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => v33a_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__17696\,
            in1 => \N__18874\,
            in2 => \N__19162\,
            in3 => \N__19211\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32166\,
            ce => \N__25310\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__19209\,
            in1 => \N__18909\,
            in2 => \N__19145\,
            in3 => \N__17684\,
            lcout => \HDA_STRAP.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32166\,
            ce => \N__25310\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__17672\,
            in1 => \N__18766\,
            in2 => \N__19161\,
            in3 => \N__19210\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32166\,
            ce => \N__25310\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__19208\,
            in1 => \N__18783\,
            in2 => \N__19144\,
            in3 => \N__17663\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32166\,
            ce => \N__25310\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_2_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19120\,
            in2 => \_gnd_net_\,
            in3 => \N__19207\,
            lcout => OPEN,
            ltout => \HDA_STRAP.N_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__15893\,
            in1 => \N__15905\,
            in2 => \N__15764\,
            in3 => \N__15970\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32166\,
            ce => \N__25310\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__15805\,
            in1 => \N__15778\,
            in2 => \N__15815\,
            in3 => \N__16492\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.delayed_vccin_okZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15761\,
            in3 => \N__29617\,
            lcout => \N_428\,
            ltout => \N_428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111000101010"
        )
    port map (
            in0 => \N__15953\,
            in1 => \N__15934\,
            in2 => \N__15758\,
            in3 => \N__19214\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32126\,
            ce => \N__25308\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIH91A_0_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15949\,
            in2 => \_gnd_net_\,
            in3 => \N__15920\,
            lcout => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_0_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001010010"
        )
    port map (
            in0 => \N__15951\,
            in1 => \N__16001\,
            in2 => \N__15933\,
            in3 => \N__19213\,
            lcout => OPEN,
            ltout => \HDA_STRAP.m14_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111001"
        )
    port map (
            in0 => \N__15935\,
            in1 => \N__15952\,
            in2 => \N__15986\,
            in3 => \N__15969\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32126\,
            ce => \N__25308\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIRV1F_2_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__15950\,
            in1 => \_gnd_net_\,
            in2 => \N__15932\,
            in3 => \N__15904\,
            lcout => \HDA_STRAP.HDA_SDO_ATP_3_0\,
            ltout => \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15887\,
            in3 => \_gnd_net_\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32126\,
            ce => \N__25308\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_0_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15869\,
            in2 => \_gnd_net_\,
            in3 => \N__15845\,
            lcout => \PCH_PWRGD.N_38_f0\,
            ltout => \PCH_PWRGD.N_38_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__15779\,
            in1 => \N__15806\,
            in2 => \N__15782\,
            in3 => \N__16495\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111010011001"
        )
    port map (
            in0 => \N__23311\,
            in1 => \N__33144\,
            in2 => \N__23267\,
            in3 => \N__25403\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001111000010"
        )
    port map (
            in0 => \N__33145\,
            in1 => \N__23312\,
            in2 => \N__15767\,
            in3 => \N__23345\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21509\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16688\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21668\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIM9AN_1_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19764\,
            in1 => \N__16009\,
            in2 => \_gnd_net_\,
            in3 => \N__16016\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_1_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__16102\,
            in1 => \N__16087\,
            in2 => \_gnd_net_\,
            in3 => \N__16385\,
            lcout => \VPP_VDDQ.count_2_1_sqmuxa\,
            ltout => \VPP_VDDQ.count_2_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__17821\,
            in1 => \_gnd_net_\,
            in2 => \N__16031\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIL8AN_0_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16022\,
            in2 => \N__16028\,
            in3 => \N__19763\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16025\,
            in3 => \N__18149\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32282\,
            ce => \N__19765\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__17816\,
            in1 => \_gnd_net_\,
            in2 => \N__18160\,
            in3 => \N__17787\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32282\,
            ce => \N__19765\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__17788\,
            in1 => \N__18145\,
            in2 => \_gnd_net_\,
            in3 => \N__17815\,
            lcout => \VPP_VDDQ.count_2_1_1\,
            ltout => \VPP_VDDQ.count_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010001"
        )
    port map (
            in0 => \N__16010\,
            in1 => \N__17820\,
            in2 => \N__16274\,
            in3 => \N__19766\,
            lcout => \VPP_VDDQ.un9_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16271\,
            in1 => \N__16238\,
            in2 => \N__16221\,
            in3 => \N__16177\,
            lcout => rsmrst_pwrgd_signal,
            ltout => \rsmrst_pwrgd_signal_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21197\,
            in2 => \N__16148\,
            in3 => \N__21168\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__21198\,
            in1 => \_gnd_net_\,
            in2 => \N__16145\,
            in3 => \N__20918\,
            lcout => \RSMRST_PWRGD_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32299\,
            ce => \N__25314\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__26804\,
            in1 => \N__21196\,
            in2 => \_gnd_net_\,
            in3 => \N__21167\,
            lcout => \RSMRST_PWRGD.N_264_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFQNU_1_7_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__17990\,
            in1 => \N__16304\,
            in2 => \N__17956\,
            in3 => \N__16283\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI0JCD2_1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19829\,
            in1 => \N__16118\,
            in2 => \N__16112\,
            in3 => \N__19619\,
            lcout => \VPP_VDDQ.N_1_i\,
            ltout => \VPP_VDDQ.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__16088\,
            in1 => \_gnd_net_\,
            in2 => \N__16049\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.N_664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18004\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32284\,
            ce => \N__19776\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__16409\,
            in1 => \N__16384\,
            in2 => \N__16340\,
            in3 => \N__16491\,
            lcout => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFQNU_7_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18050\,
            in2 => \N__16316\,
            in3 => \N__16297\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJ0QU_9_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18005\,
            in1 => \N__16313\,
            in2 => \_gnd_net_\,
            in3 => \N__19779\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => \VPP_VDDQ.count_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__19778\,
            in1 => \N__18049\,
            in2 => \N__16307\,
            in3 => \N__16298\,
            lcout => \VPP_VDDQ.un9_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18043\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32284\,
            ce => \N__19776\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI52L41_11_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19777\,
            in1 => \N__16289\,
            in2 => \_gnd_net_\,
            in3 => \N__17939\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32284\,
            ce => \N__19776\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_15_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17872\,
            in1 => \N__17923\,
            in2 => \N__17900\,
            in3 => \N__18217\,
            lcout => \VPP_VDDQ.un9_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI75M41_12_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17912\,
            in1 => \N__16592\,
            in2 => \_gnd_net_\,
            in3 => \N__19800\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17911\,
            lcout => \VPP_VDDQ.count_2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32397\,
            ce => \N__19799\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI98N41_13_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17885\,
            in1 => \N__16586\,
            in2 => \_gnd_net_\,
            in3 => \N__19801\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17884\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32397\,
            ce => \N__19799\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIBBO41_14_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17861\,
            in1 => \N__16580\,
            in2 => \_gnd_net_\,
            in3 => \N__19802\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17860\,
            lcout => \VPP_VDDQ.count_2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32397\,
            ce => \N__19799\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIDEP41_15_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19753\,
            in1 => \N__18110\,
            in2 => \_gnd_net_\,
            in3 => \N__18121\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__17603\,
            in1 => \N__16574\,
            in2 => \_gnd_net_\,
            in3 => \N__16532\,
            lcout => \POWERLED.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32406\,
            ce => \N__16461\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI7EJU_3_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19772\,
            in1 => \N__17720\,
            in2 => \_gnd_net_\,
            in3 => \N__17767\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIBKLU_5_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17849\,
            in1 => \N__19773\,
            in2 => \_gnd_net_\,
            in3 => \N__17749\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIHTOU_8_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19774\,
            in1 => \N__17840\,
            in2 => \_gnd_net_\,
            in3 => \N__18029\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIS3FU_10_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17831\,
            in1 => \N__17974\,
            in2 => \_gnd_net_\,
            in3 => \N__19775\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16684\,
            in2 => \_gnd_net_\,
            in3 => \N__16754\,
            lcout => \POWERLED.mult1_un124_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16683\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21530\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16643\,
            in2 => \N__16631\,
            in3 => \N__16619\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16750\,
            in2 => \N__16616\,
            in3 => \N__16604\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16670\,
            in2 => \N__16736\,
            in3 => \N__16601\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16724\,
            in2 => \N__16682\,
            in3 => \N__16598\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18371\,
            in1 => \N__16760\,
            in2 => \N__16715\,
            in3 => \N__16595\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16700\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16763\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__16711\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16669\,
            lcout => \POWERLED.mult1_un124_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21502\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20378\,
            in2 => \N__16858\,
            in3 => \N__16739\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16854\,
            in2 => \N__16841\,
            in3 => \N__16727\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16829\,
            in2 => \N__16790\,
            in3 => \N__16718\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16820\,
            in2 => \N__16789\,
            in3 => \N__16703\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16668\,
            in1 => \N__16811\,
            in2 => \N__16859\,
            in3 => \N__16694\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16691\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16782\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21482\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20399\,
            in2 => \N__16876\,
            in3 => \N__16832\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16872\,
            in2 => \N__16937\,
            in3 => \N__16823\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16925\,
            in2 => \N__18410\,
            in3 => \N__16814\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18408\,
            in2 => \N__16916\,
            in3 => \N__16805\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16781\,
            in1 => \N__16904\,
            in2 => \N__16877\,
            in3 => \N__16796\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16895\,
            in3 => \N__16793\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => \POWERLED.mult1_un110_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16940\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un110_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21758\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18437\,
            in2 => \N__18427\,
            in3 => \N__16928\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18423\,
            in2 => \N__18329\,
            in3 => \N__16919\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18317\,
            in2 => \N__18508\,
            in3 => \N__16907\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18504\,
            in2 => \N__18548\,
            in3 => \N__16898\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18404\,
            in1 => \N__18536\,
            in2 => \N__18428\,
            in3 => \N__16886\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18527\,
            in3 => \N__16883\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => \POWERLED.mult1_un103_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16880\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17261\,
            in1 => \N__18290\,
            in2 => \N__17231\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17222\,
            in1 => \N__18443\,
            in2 => \N__17195\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5036_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_0\,
            carryout => \POWERLED.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18281\,
            in2 => \N__17150\,
            in3 => \N__17183\,
            lcout => \POWERLED.N_5037_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_1\,
            carryout => \POWERLED.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18272\,
            in2 => \N__17111\,
            in3 => \N__17141\,
            lcout => \POWERLED.N_5038_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_2\,
            carryout => \POWERLED.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18449\,
            in2 => \N__17075\,
            in3 => \N__17102\,
            lcout => \POWERLED.N_5039_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_3\,
            carryout => \POWERLED.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18476\,
            in2 => \N__17033\,
            in3 => \N__17066\,
            lcout => \POWERLED.N_5040_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_4\,
            carryout => \POWERLED.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17024\,
            in1 => \N__18335\,
            in2 => \N__16994\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5041_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_5\,
            carryout => \POWERLED.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16982\,
            in1 => \N__16958\,
            in2 => \N__16949\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5042_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_6\,
            carryout => \POWERLED.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17507\,
            in2 => \N__17546\,
            in3 => \N__17534\,
            lcout => \POWERLED.N_5043_i\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17474\,
            in2 => \N__18386\,
            in3 => \N__17501\,
            lcout => \POWERLED.N_5044_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_8\,
            carryout => \POWERLED.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17468\,
            in1 => \N__17420\,
            in2 => \N__17435\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5045_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_9\,
            carryout => \POWERLED.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17573\,
            in2 => \N__17384\,
            in3 => \N__17414\,
            lcout => \POWERLED.N_5046_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_10\,
            carryout => \POWERLED.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18557\,
            in2 => \N__17345\,
            in3 => \N__17375\,
            lcout => \POWERLED.N_5047_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_11\,
            carryout => \POWERLED.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17303\,
            in2 => \N__18593\,
            in3 => \N__17333\,
            lcout => \POWERLED.N_5048_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_12\,
            carryout => \POWERLED.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17297\,
            in1 => \N__17267\,
            in2 => \N__17567\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5049_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_13\,
            carryout => \POWERLED.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20366\,
            in2 => \N__17621\,
            in3 => \N__17648\,
            lcout => \POWERLED.N_5050_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_14\,
            carryout => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17612\,
            lcout => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18637\,
            lcout => \POWERLED.mult1_un89_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20603\,
            lcout => \POWERLED.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_0_c_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19259\,
            in2 => \N__19163\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_1_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19273\,
            in2 => \_gnd_net_\,
            in3 => \N__17558\,
            lcout => \HDA_STRAP.countZ0Z_1\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_0\,
            carryout => \HDA_STRAP.un1_count_1_cry_1\,
            clk => \N__32053\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18829\,
            in2 => \_gnd_net_\,
            in3 => \N__17555\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_1\,
            carryout => \HDA_STRAP.un1_count_1_cry_2\,
            clk => \N__32053\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18814\,
            in2 => \_gnd_net_\,
            in3 => \N__17552\,
            lcout => \HDA_STRAP.countZ0Z_3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_2\,
            carryout => \HDA_STRAP.un1_count_1_cry_3\,
            clk => \N__32053\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18842\,
            in2 => \_gnd_net_\,
            in3 => \N__17549\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_3\,
            carryout => \HDA_STRAP.un1_count_1_cry_4\,
            clk => \N__32053\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18803\,
            in2 => \_gnd_net_\,
            in3 => \N__17699\,
            lcout => \HDA_STRAP.countZ0Z_5\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_4\,
            carryout => \HDA_STRAP.un1_count_1_cry_5\,
            clk => \N__32053\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18873\,
            in2 => \_gnd_net_\,
            in3 => \N__17690\,
            lcout => \HDA_STRAP.un1_count_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_5\,
            carryout => \HDA_STRAP.un1_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18692\,
            in2 => \_gnd_net_\,
            in3 => \N__17687\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_6\,
            carryout => \HDA_STRAP.un1_count_1_cry_7\,
            clk => \N__32053\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18911\,
            in2 => \_gnd_net_\,
            in3 => \N__17678\,
            lcout => \HDA_STRAP.un1_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18731\,
            in2 => \_gnd_net_\,
            in3 => \N__17675\,
            lcout => \HDA_STRAP.countZ0Z_9\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_8\,
            carryout => \HDA_STRAP.un1_count_1_cry_9\,
            clk => \N__32220\,
            ce => \N__25315\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18765\,
            in2 => \_gnd_net_\,
            in3 => \N__17666\,
            lcout => \HDA_STRAP.un1_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_9\,
            carryout => \HDA_STRAP.un1_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18791\,
            in2 => \_gnd_net_\,
            in3 => \N__17657\,
            lcout => \HDA_STRAP.un1_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_10\,
            carryout => \HDA_STRAP.un1_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18719\,
            in2 => \_gnd_net_\,
            in3 => \N__17654\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_11\,
            carryout => \HDA_STRAP.un1_count_1_cry_12\,
            clk => \N__32220\,
            ce => \N__25315\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18706\,
            in2 => \_gnd_net_\,
            in3 => \N__17651\,
            lcout => \HDA_STRAP.countZ0Z_13\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_12\,
            carryout => \HDA_STRAP.un1_count_1_cry_13\,
            clk => \N__32220\,
            ce => \N__25315\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18890\,
            in2 => \_gnd_net_\,
            in3 => \N__17711\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_13\,
            carryout => \HDA_STRAP.un1_count_1_cry_14\,
            clk => \N__32220\,
            ce => \N__25315\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18854\,
            in2 => \_gnd_net_\,
            in3 => \N__17708\,
            lcout => \HDA_STRAP.countZ0Z_15\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_14\,
            carryout => \HDA_STRAP.un1_count_1_cry_15\,
            clk => \N__32220\,
            ce => \N__25315\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19076\,
            in2 => \_gnd_net_\,
            in3 => \N__17705\,
            lcout => \HDA_STRAP.un1_count_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__19140\,
            in1 => \N__19234\,
            in2 => \N__19212\,
            in3 => \N__17702\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32226\,
            ce => \N__25312\,
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__19059\,
            in1 => \_gnd_net_\,
            in2 => \N__22550\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22543\,
            in1 => \N__18920\,
            in2 => \_gnd_net_\,
            in3 => \N__18934\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__19014\,
            in1 => \N__18998\,
            in2 => \_gnd_net_\,
            in3 => \N__22547\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19321\,
            in1 => \N__19354\,
            in2 => \N__19340\,
            in3 => \N__19369\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18984\,
            in1 => \N__18957\,
            in2 => \N__19016\,
            in3 => \N__19058\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__19384\,
            in1 => \N__19410\,
            in2 => \N__19039\,
            in3 => \N__18933\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18944\,
            in1 => \N__18958\,
            in2 => \_gnd_net_\,
            in3 => \N__22548\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20945\,
            in2 => \_gnd_net_\,
            in3 => \N__25402\,
            lcout => \RSMRST_PWRGD.N_92_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19465\,
            in1 => \N__19288\,
            in2 => \N__19307\,
            in3 => \N__19450\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__19038\,
            in1 => \N__22538\,
            in2 => \_gnd_net_\,
            in3 => \N__19061\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18968\,
            in1 => \N__18986\,
            in2 => \_gnd_net_\,
            in3 => \N__22539\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22537\,
            in1 => \N__19394\,
            in2 => \_gnd_net_\,
            in3 => \N__19414\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19603\,
            in1 => \N__19555\,
            in2 => \N__19574\,
            in3 => \N__19588\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__26805\,
            in1 => \N__21195\,
            in2 => \_gnd_net_\,
            in3 => \N__21169\,
            lcout => \N_555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17768\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32283\,
            ce => \N__19780\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17750\,
            lcout => \VPP_VDDQ.count_2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32283\,
            ce => \N__19780\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18028\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32283\,
            ce => \N__19780\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17975\,
            lcout => \VPP_VDDQ.count_2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32283\,
            ce => \N__19780\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17822\,
            in2 => \N__17795\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18193\,
            in1 => \N__19685\,
            in2 => \_gnd_net_\,
            in3 => \N__17771\,
            lcout => \VPP_VDDQ.count_2_1_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18201\,
            in1 => \N__19630\,
            in2 => \_gnd_net_\,
            in3 => \N__17756\,
            lcout => \VPP_VDDQ.count_2_1_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18194\,
            in1 => \N__19859\,
            in2 => \_gnd_net_\,
            in3 => \N__17753\,
            lcout => \VPP_VDDQ.count_2_1_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18202\,
            in1 => \N__19672\,
            in2 => \_gnd_net_\,
            in3 => \N__17738\,
            lcout => \VPP_VDDQ.count_2_1_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIDNMU_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18195\,
            in1 => \N__19880\,
            in2 => \_gnd_net_\,
            in3 => \N__17735\,
            lcout => \VPP_VDDQ.count_2_1_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18203\,
            in1 => \N__18059\,
            in2 => \_gnd_net_\,
            in3 => \N__18032\,
            lcout => \VPP_VDDQ.count_2_1_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__18196\,
            in1 => \_gnd_net_\,
            in2 => \N__19657\,
            in3 => \N__18017\,
            lcout => \VPP_VDDQ.count_2_1_8\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18205\,
            in1 => \N__18014\,
            in2 => \_gnd_net_\,
            in3 => \N__17993\,
            lcout => \VPP_VDDQ.count_2_1_9\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18197\,
            in1 => \N__17986\,
            in2 => \_gnd_net_\,
            in3 => \N__17960\,
            lcout => \VPP_VDDQ.count_2_1_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18204\,
            in1 => \N__17957\,
            in2 => \_gnd_net_\,
            in3 => \N__17927\,
            lcout => \VPP_VDDQ.count_2_1_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18198\,
            in1 => \N__17924\,
            in2 => \_gnd_net_\,
            in3 => \N__17903\,
            lcout => \VPP_VDDQ.count_2_1_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18206\,
            in1 => \N__17899\,
            in2 => \_gnd_net_\,
            in3 => \N__17876\,
            lcout => \VPP_VDDQ.count_2_1_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18199\,
            in1 => \N__17873\,
            in2 => \_gnd_net_\,
            in3 => \N__17852\,
            lcout => \VPP_VDDQ.count_2_1_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__18218\,
            in1 => \N__18200\,
            in2 => \_gnd_net_\,
            in3 => \N__18125\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18122\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32350\,
            ce => \N__19781\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21551\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20387\,
            in2 => \N__18261\,
            in3 => \N__18104\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18101\,
            in2 => \N__18263\,
            in3 => \N__18095\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18092\,
            in2 => \N__18373\,
            in3 => \N__18086\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18083\,
            in2 => \N__18372\,
            in3 => \N__18077\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20062\,
            in1 => \N__18074\,
            in2 => \N__18262\,
            in3 => \N__18068\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18065\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18266\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18361\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21587\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19890\,
            in2 => \N__20183\,
            in3 => \N__18239\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2_c\,
            carryout => \POWERLED.mult1_un145_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20015\,
            in2 => \N__19895\,
            in3 => \N__18236\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3_c\,
            carryout => \POWERLED.mult1_un145_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19917\,
            in2 => \N__20000\,
            in3 => \N__18233\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4_c\,
            carryout => \POWERLED.mult1_un145_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19979\,
            in2 => \N__19924\,
            in3 => \N__18230\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5_c\,
            carryout => \POWERLED.mult1_un145_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20132\,
            in1 => \N__19894\,
            in2 => \N__19964\,
            in3 => \N__18227\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6_c\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18224\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => \POWERLED.mult1_un145_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18221\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26558\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22754\,
            in2 => \N__18310\,
            in3 => \N__20258\,
            lcout => \G_2150\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18306\,
            in2 => \N__20351\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20259\,
            in2 => \N__20333\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20315\,
            in2 => \N__20266\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20300\,
            in2 => \N__18311\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__20285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18293\,
            lcout => \POWERLED.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20235\,
            lcout => \POWERLED.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20141\,
            lcout => \POWERLED.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19928\,
            lcout => \POWERLED.mult1_un138_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20267\,
            lcout => \POWERLED.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21739\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18499\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18409\,
            lcout => \POWERLED.mult1_un103_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21740\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18566\,
            in2 => \N__18610\,
            in3 => \N__18320\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18606\,
            in2 => \N__18470\,
            in3 => \N__18551\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18458\,
            in2 => \N__18638\,
            in3 => \N__18539\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18636\,
            in2 => \N__18674\,
            in3 => \N__18530\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18500\,
            in1 => \N__18662\,
            in2 => \N__18611\,
            in3 => \N__18518\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18653\,
            in3 => \N__18515\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20072\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21715\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21788\,
            in2 => \N__18583\,
            in3 => \N__18461\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18579\,
            in2 => \N__20519\,
            in3 => \N__18452\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20498\,
            in2 => \N__20654\,
            in3 => \N__18665\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20653\,
            in2 => \N__20483\,
            in3 => \N__18656\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18632\,
            in1 => \N__20711\,
            in2 => \N__18584\,
            in3 => \N__18644\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20678\,
            in3 => \N__18641\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => \POWERLED.mult1_un89_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18614\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20743\,
            lcout => \POWERLED.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20647\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21716\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20648\,
            lcout => \POWERLED.mult1_un82_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21977\,
            lcout => \POWERLED.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31836\,
            ce => \N__23545\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22052\,
            lcout => \POWERLED.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31836\,
            ce => \N__23545\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDLB61_6_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__18910\,
            in1 => \N__18889\,
            in2 => \N__18878\,
            in3 => \N__18853\,
            lcout => \HDA_STRAP.un4_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI2L821_2_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18841\,
            in1 => \N__18830\,
            in2 => \N__18818\,
            in3 => \N__18802\,
            lcout => \HDA_STRAP.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIH7IR1_10_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18790\,
            in1 => \N__18767\,
            in2 => \_gnd_net_\,
            in3 => \N__19220\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB5IA5_2_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18746\,
            in1 => \N__18680\,
            in2 => \N__18740\,
            in3 => \N__18737\,
            lcout => \HDA_STRAP.un4_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIBJB61_7_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18730\,
            in1 => \N__18718\,
            in2 => \N__18707\,
            in3 => \N__18691\,
            lcout => \HDA_STRAP.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_0_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__19254\,
            in1 => \N__19150\,
            in2 => \N__19160\,
            in3 => \N__19198\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32225\,
            ce => \N__25313\,
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19502\,
            in1 => \N__19481\,
            in2 => \N__19541\,
            in3 => \N__19520\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI4CB61_17_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__19074\,
            in1 => \N__19274\,
            in2 => \N__19258\,
            in3 => \N__19235\,
            lcout => \HDA_STRAP.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__19197\,
            in1 => \N__19146\,
            in2 => \N__19085\,
            in3 => \N__19075\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32225\,
            ce => \N__25313\,
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19060\,
            in2 => \N__19040\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19015\,
            in2 => \_gnd_net_\,
            in3 => \N__18989\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18985\,
            in2 => \_gnd_net_\,
            in3 => \N__18962\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18959\,
            in2 => \_gnd_net_\,
            in3 => \N__18938\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18935\,
            in2 => \_gnd_net_\,
            in3 => \N__18914\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19415\,
            in3 => \N__19388\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19385\,
            in2 => \_gnd_net_\,
            in3 => \N__19373\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__32224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19370\,
            in2 => \_gnd_net_\,
            in3 => \N__19358\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__32224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19355\,
            in2 => \_gnd_net_\,
            in3 => \N__19343\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19339\,
            in2 => \_gnd_net_\,
            in3 => \N__19325\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19322\,
            in2 => \_gnd_net_\,
            in3 => \N__19310\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19306\,
            in2 => \_gnd_net_\,
            in3 => \N__19292\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19289\,
            in2 => \_gnd_net_\,
            in3 => \N__19277\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19466\,
            in2 => \_gnd_net_\,
            in3 => \N__19454\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19451\,
            in2 => \_gnd_net_\,
            in3 => \N__19439\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21035\,
            in2 => \_gnd_net_\,
            in3 => \N__19436\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__32227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21062\,
            in2 => \_gnd_net_\,
            in3 => \N__19433\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21049\,
            in2 => \_gnd_net_\,
            in3 => \N__19430\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21074\,
            in2 => \_gnd_net_\,
            in3 => \N__19427\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21011\,
            in2 => \_gnd_net_\,
            in3 => \N__19424\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20998\,
            in2 => \_gnd_net_\,
            in3 => \N__19421\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20984\,
            in2 => \_gnd_net_\,
            in3 => \N__19418\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21023\,
            in2 => \_gnd_net_\,
            in3 => \N__19607\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19604\,
            in2 => \_gnd_net_\,
            in3 => \N__19592\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__32180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19589\,
            in2 => \_gnd_net_\,
            in3 => \N__19577\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__32052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19573\,
            in2 => \_gnd_net_\,
            in3 => \N__19559\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__32052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19556\,
            in2 => \_gnd_net_\,
            in3 => \N__19544\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__32052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19537\,
            in2 => \_gnd_net_\,
            in3 => \N__19523\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__32052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19519\,
            in2 => \_gnd_net_\,
            in3 => \N__19505\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__32052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19501\,
            in2 => \_gnd_net_\,
            in3 => \N__19487\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__32052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19480\,
            in2 => \_gnd_net_\,
            in3 => \N__19484\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32206\,
            ce => \N__19798\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32206\,
            ce => \N__19798\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIREAN_6_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19852\,
            in1 => \N__19784\,
            in2 => \_gnd_net_\,
            in3 => \N__19839\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI9HKU_4_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19783\,
            in1 => \N__19874\,
            in2 => \_gnd_net_\,
            in3 => \N__19867\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => \VPP_VDDQ.count_2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIREAN_0_6_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__19853\,
            in1 => \N__19785\,
            in2 => \N__19844\,
            in3 => \N__19841\,
            lcout => \VPP_VDDQ.un9_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32206\,
            ce => \N__19798\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI5BIU_2_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19817\,
            in1 => \N__19810\,
            in2 => \_gnd_net_\,
            in3 => \N__19782\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => \VPP_VDDQ.count_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_2_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19679\,
            in1 => \N__19661\,
            in2 => \N__19640\,
            in3 => \N__19637\,
            lcout => \VPP_VDDQ.un9_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21569\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20420\,
            in2 => \N__20037\,
            in3 => \N__20009\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20006\,
            in2 => \N__20039\,
            in3 => \N__19991\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20063\,
            in2 => \N__19988\,
            in3 => \N__19973\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19970\,
            in2 => \N__20071\,
            in3 => \N__19955\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19916\,
            in1 => \N__19952\,
            in2 => \N__20038\,
            in3 => \N__19940\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19937\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19931\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => \POWERLED.mult1_un138_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19898\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_2_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32955\,
            in2 => \_gnd_net_\,
            in3 => \N__29442\,
            lcout => \POWERLED.N_613\,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20106\,
            in2 => \N__20411\,
            in3 => \N__20171\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20168\,
            in2 => \N__20111\,
            in3 => \N__20162\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20133\,
            in2 => \N__20159\,
            in3 => \N__20150\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20147\,
            in2 => \N__20140\,
            in3 => \N__20114\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20227\,
            in1 => \N__20110\,
            in2 => \N__20096\,
            in3 => \N__20084\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20075\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20067\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30929\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20196\,
            in2 => \N__22592\,
            in3 => \N__20342\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20339\,
            in2 => \N__20203\,
            in3 => \N__20324\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20321\,
            in2 => \N__20237\,
            in3 => \N__20309\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20306\,
            in2 => \N__20236\,
            in3 => \N__20294\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20257\,
            in1 => \N__20291\,
            in2 => \N__20204\,
            in3 => \N__20279\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20270\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20228\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21565\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21544\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21580\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21757\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21523\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21478\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21615\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21614\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21829\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21764\,
            in2 => \N__20461\,
            in3 => \N__20354\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20457\,
            in2 => \N__21431\,
            in3 => \N__20471\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21407\,
            in2 => \N__21626\,
            in3 => \N__20468\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21625\,
            in2 => \N__21389\,
            in3 => \N__20465\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20591\,
            in1 => \N__21365\,
            in2 => \N__20462\,
            in3 => \N__20444\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21344\,
            in2 => \_gnd_net_\,
            in3 => \N__20441\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => \POWERLED.mult1_un68_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20438\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21688\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21818\,
            in2 => \N__20554\,
            in3 => \N__20435\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20550\,
            in2 => \N__20432\,
            in3 => \N__20423\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20612\,
            in2 => \N__20599\,
            in3 => \N__20606\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20595\,
            in2 => \N__20573\,
            in3 => \N__20564\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20738\,
            in1 => \N__20561\,
            in2 => \N__20555\,
            in3 => \N__20537\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20534\,
            in3 => \N__20525\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => \POWERLED.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20522\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21806\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_16_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20627\,
            in2 => \N__20695\,
            in3 => \N__20510\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20691\,
            in2 => \N__20507\,
            in3 => \N__20492\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20489\,
            in2 => \N__20744\,
            in3 => \N__20474\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20742\,
            in2 => \N__20720\,
            in3 => \N__20705\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20649\,
            in1 => \N__20702\,
            in2 => \N__20696\,
            in3 => \N__20669\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20666\,
            in3 => \N__20657\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21692\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32045\,
            ce => \N__23546\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIN3TIG_9_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20621\,
            in1 => \N__23541\,
            in2 => \_gnd_net_\,
            in3 => \N__20872\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => \POWERLED.count_offZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_10_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20794\,
            in1 => \N__20854\,
            in2 => \N__20615\,
            in3 => \N__20824\,
            lcout => \POWERLED.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI0E2HG_10_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20771\,
            in1 => \N__20839\,
            in2 => \_gnd_net_\,
            in3 => \N__23542\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32045\,
            ce => \N__23546\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI9LFFG_11_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20765\,
            in1 => \N__20809\,
            in2 => \_gnd_net_\,
            in3 => \N__23543\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20810\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32045\,
            ce => \N__23546\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIBOGFG_12_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21083\,
            in1 => \N__21098\,
            in2 => \_gnd_net_\,
            in3 => \N__23544\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23396\,
            in2 => \N__22090\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNI5IAA7_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26130\,
            in1 => \N__21919\,
            in2 => \_gnd_net_\,
            in3 => \N__20759\,
            lcout => \POWERLED.count_off_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_1_cZ0\,
            carryout => \POWERLED.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23210\,
            in2 => \_gnd_net_\,
            in3 => \N__20756\,
            lcout => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_2\,
            carryout => \POWERLED.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23606\,
            in2 => \_gnd_net_\,
            in3 => \N__20753\,
            lcout => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_3\,
            carryout => \POWERLED.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_4_c_RNI8ODA7_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26126\,
            in1 => \N__21959\,
            in2 => \_gnd_net_\,
            in3 => \N__20750\,
            lcout => \POWERLED.count_off_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_4\,
            carryout => \POWERLED.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNI9QEA7_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26128\,
            in1 => \N__22036\,
            in2 => \_gnd_net_\,
            in3 => \N__20747\,
            lcout => \POWERLED.count_off_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_5\,
            carryout => \POWERLED.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNIASFA7_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26127\,
            in1 => \N__23191\,
            in2 => \_gnd_net_\,
            in3 => \N__20888\,
            lcout => \POWERLED.count_off_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_6\,
            carryout => \POWERLED.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_7_c_RNIBUGA7_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26129\,
            in1 => \N__23167\,
            in2 => \_gnd_net_\,
            in3 => \N__20885\,
            lcout => \POWERLED.count_off_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_7\,
            carryout => \POWERLED.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNIC0IA7_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26119\,
            in1 => \N__20882\,
            in2 => \_gnd_net_\,
            in3 => \N__20861\,
            lcout => \POWERLED.count_off_1_9\,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_9_c_RNID2JA7_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26122\,
            in1 => \_gnd_net_\,
            in2 => \N__20858\,
            in3 => \N__20828\,
            lcout => \POWERLED.count_off_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_9\,
            carryout => \POWERLED.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNIL8097_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26120\,
            in1 => \N__20825\,
            in2 => \_gnd_net_\,
            in3 => \N__20798\,
            lcout => \POWERLED.count_off_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_10\,
            carryout => \POWERLED.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_11_c_RNIMA197_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26123\,
            in1 => \N__20795\,
            in2 => \_gnd_net_\,
            in3 => \N__20780\,
            lcout => \POWERLED.count_off_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_11\,
            carryout => \POWERLED.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_12_c_RNINC297_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26121\,
            in1 => \N__22117\,
            in2 => \_gnd_net_\,
            in3 => \N__20777\,
            lcout => \POWERLED.count_off_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_12\,
            carryout => \POWERLED.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_13_c_RNIOE397_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26124\,
            in1 => \N__22105\,
            in2 => \_gnd_net_\,
            in3 => \N__20774\,
            lcout => \POWERLED.count_off_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_13\,
            carryout => \POWERLED.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_14_c_RNIPG497_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__22124\,
            in1 => \N__26125\,
            in2 => \_gnd_net_\,
            in3 => \N__21101\,
            lcout => \POWERLED.un3_count_off_1_cry_14_c_RNIPGZ0Z497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21097\,
            lcout => \POWERLED.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32046\,
            ce => \N__23537\,
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__25620\,
            in1 => \_gnd_net_\,
            in2 => \N__22524\,
            in3 => \_gnd_net_\,
            lcout => \clk_100Khz_signalkeep_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_en_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__29557\,
            in1 => \N__25619\,
            in2 => \N__30739\,
            in3 => \N__22504\,
            lcout => \POWERLED.func_state_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21073\,
            in1 => \N__21061\,
            in2 => \N__21050\,
            in3 => \N__21034\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21022\,
            in1 => \N__21010\,
            in2 => \N__20999\,
            in3 => \N__20983\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_14_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__21213\,
            in1 => \N__20910\,
            in2 => \N__20972\,
            in3 => \N__25399\,
            lcout => \G_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__26824\,
            in1 => \N__21216\,
            in2 => \N__20917\,
            in3 => \N__21152\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32179\,
            ce => \N__25311\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21148\,
            in1 => \N__26821\,
            in2 => \_gnd_net_\,
            in3 => \N__21217\,
            lcout => \RSMRSTn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32179\,
            ce => \N__25311\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__26822\,
            in1 => \N__21215\,
            in2 => \_gnd_net_\,
            in3 => \N__21151\,
            lcout => \RSMRSTn_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32179\,
            ce => \N__25311\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21149\,
            in1 => \N__26823\,
            in2 => \_gnd_net_\,
            in3 => \N__21218\,
            lcout => \RSMRSTn_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32179\,
            ce => \N__25311\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__26820\,
            in1 => \N__21214\,
            in2 => \_gnd_net_\,
            in3 => \N__21150\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32179\,
            ce => \N__25311\,
            sr => \_gnd_net_\
        );

    \POWERLED.N_430_i_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__26747\,
            in1 => \N__26367\,
            in2 => \N__27617\,
            in3 => \N__25658\,
            lcout => \POWERLED.N_430_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.VCCST_EN_i_0_o2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30575\,
            in2 => \_gnd_net_\,
            in3 => \N__29844\,
            lcout => \VCCST_EN_i_1\,
            ltout => \VCCST_EN_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21113\,
            in1 => \N__28813\,
            in2 => \N__21119\,
            in3 => \N__28590\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_o_N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__21107\,
            in1 => \N__25988\,
            in2 => \N__21116\,
            in3 => \N__23738\,
            lcout => \POWERLED.un1_func_state25_6_0_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_0_o2_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__30420\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26748\,
            lcout => \POWERLED.N_432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__30577\,
            in2 => \N__26756\,
            in3 => \N__30421\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__30576\,
            in1 => \N__27574\,
            in2 => \N__30422\,
            in3 => \N__26235\,
            lcout => \POWERLED.func_state_RNIBVNSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI78D82_1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__22426\,
            in1 => \N__21257\,
            in2 => \N__30074\,
            in3 => \N__25655\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_ss0_i_0_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3H2K3_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__28814\,
            in1 => \N__21251\,
            in2 => \N__21260\,
            in3 => \N__25874\,
            lcout => \POWERLED.N_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_215_i_0_o2_0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__30388\,
            in1 => \N__30722\,
            in2 => \N__27663\,
            in3 => \N__26752\,
            lcout => \POWERLED.N_423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMJ6IF_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__21241\,
            in1 => \N__33067\,
            in2 => \N__21230\,
            in3 => \N__22396\,
            lcout => \func_state_RNIMJ6IF_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_1_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__30389\,
            in1 => \N__30723\,
            in2 => \N__27664\,
            in3 => \N__28815\,
            lcout => \POWERLED.N_673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIP4521_0_1_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__25656\,
            in1 => \N__27640\,
            in2 => \N__26383\,
            in3 => \N__30022\,
            lcout => \POWERLED.N_542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_0_a2_5_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__26753\,
            in1 => \N__25657\,
            in2 => \N__27665\,
            in3 => \N__26371\,
            lcout => \POWERLED.N_671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__21229\,
            in1 => \N__33068\,
            in2 => \N__21245\,
            in3 => \N__22397\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_11_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011001100"
        )
    port map (
            in0 => \N__29862\,
            in1 => \N__30266\,
            in2 => \N__29742\,
            in3 => \N__24703\,
            lcout => OPEN,
            ltout => \POWERLED.N_512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5TUF2_11_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24704\,
            in1 => \N__27452\,
            in2 => \N__21302\,
            in3 => \N__30014\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_39_and_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRUFD6_11_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__32629\,
            in1 => \N__32812\,
            in2 => \N__21299\,
            in3 => \N__21296\,
            lcout => \POWERLED.dutycycle_en_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_10_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101010"
        )
    port map (
            in0 => \N__27878\,
            in1 => \N__33086\,
            in2 => \N__24815\,
            in3 => \N__27834\,
            lcout => \POWERLED.N_508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_11_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__24702\,
            in1 => \N__33085\,
            in2 => \N__27892\,
            in3 => \N__27833\,
            lcout => \POWERLED.N_514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5TUF2_10_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__24813\,
            in1 => \N__30073\,
            in2 => \N__27461\,
            in3 => \N__23801\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_33_and_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRUFD6_10_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__21290\,
            in1 => \N__32630\,
            in2 => \N__21284\,
            in3 => \N__32813\,
            lcout => \POWERLED.dutycycle_en_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJTQIG_7_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21266\,
            in1 => \N__23520\,
            in2 => \_gnd_net_\,
            in3 => \N__21280\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32322\,
            ce => \N__23538\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIL0SIG_8_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21320\,
            in1 => \N__23521\,
            in2 => \_gnd_net_\,
            in3 => \N__21331\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21332\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32322\,
            ce => \N__23538\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000101"
        )
    port map (
            in0 => \N__22812\,
            in1 => \_gnd_net_\,
            in2 => \N__22790\,
            in3 => \N__21853\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22813\,
            in2 => \N__21857\,
            in3 => \N__22789\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22811\,
            lcout => \POWERLED.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21658\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21596\,
            in3 => \N__21314\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22871\,
            in2 => \N__22853\,
            in3 => \N__21311\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25182\,
            in2 => \N__22709\,
            in3 => \N__21308\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25194\,
            in2 => \N__22688\,
            in3 => \N__21305\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22632\,
            in1 => \N__22667\,
            in2 => \N__21455\,
            in3 => \N__21461\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21458\,
            lcout => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__22665\,
            in1 => \N__22666\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21779\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21446\,
            in2 => \N__22615\,
            in3 => \N__21419\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22611\,
            in2 => \N__21416\,
            in3 => \N__21398\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21395\,
            in2 => \N__22637\,
            in3 => \N__21377\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22636\,
            in2 => \N__21374\,
            in3 => \N__21353\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21616\,
            in1 => \N__21350\,
            in2 => \N__22616\,
            in3 => \N__21335\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21638\,
            in3 => \N__21629\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22744\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_53_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26548\,
            in2 => \N__31028\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_53_axb_0\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22844\,
            in2 => \N__26557\,
            in3 => \N__21554\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32949\,
            in2 => \N__22826\,
            in3 => \N__21533\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_1\,
            carryout => \POWERLED.un1_dutycycle_53_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32858\,
            in2 => \N__32957\,
            in3 => \N__21512\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_2\,
            carryout => \POWERLED.un1_dutycycle_53_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31169\,
            in2 => \N__31186\,
            in3 => \N__21485\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_3\,
            carryout => \POWERLED.un1_dutycycle_53_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31321\,
            in2 => \N__22835\,
            in3 => \N__21464\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_4\,
            carryout => \POWERLED.un1_dutycycle_53_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31314\,
            in2 => \N__22976\,
            in3 => \N__21743\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_5\,
            carryout => \POWERLED.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22988\,
            in2 => \N__24809\,
            in3 => \N__21719\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_6\,
            carryout => \POWERLED.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24701\,
            in2 => \N__24203\,
            in3 => \N__21698\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26973\,
            in2 => \N__22952\,
            in3 => \N__21695\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_8\,
            carryout => \POWERLED.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24093\,
            in2 => \N__22898\,
            in3 => \N__21677\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_9\,
            carryout => \POWERLED.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27747\,
            in2 => \N__24254\,
            in3 => \N__21674\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_10\,
            carryout => \POWERLED.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27506\,
            in2 => \N__23063\,
            in3 => \N__21671\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_11\,
            carryout => \POWERLED.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24094\,
            in2 => \N__24278\,
            in3 => \N__21644\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_12\,
            carryout => \POWERLED.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23030\,
            in2 => \N__27763\,
            in3 => \N__21641\,
            lcout => \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_13\,
            carryout => \POWERLED.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21812\,
            in2 => \N__27519\,
            in3 => \N__21866\,
            lcout => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_14\,
            carryout => \POWERLED.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27510\,
            in2 => \N__21839\,
            in3 => \N__21863\,
            lcout => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21860\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27746\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23096\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21830\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_15_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27745\,
            in1 => \N__27511\,
            in2 => \_gnd_net_\,
            in3 => \N__23095\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21802\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI12AS_8_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__30602\,
            in1 => \N__24441\,
            in2 => \_gnd_net_\,
            in3 => \N__29894\,
            lcout => \POWERLED.N_599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21778\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI99TE_13_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__21878\,
            in1 => \N__30550\,
            in2 => \_gnd_net_\,
            in3 => \N__27677\,
            lcout => OPEN,
            ltout => \POWERLED.N_598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIAB7B1_13_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__27236\,
            in1 => \N__24115\,
            in2 => \N__21893\,
            in3 => \N__27836\,
            lcout => OPEN,
            ltout => \POWERLED.N_450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI35P35_13_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__22352\,
            in1 => \N__32843\,
            in2 => \N__21890\,
            in3 => \N__32673\,
            lcout => \POWERLED.dutycycle_en_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_8_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__27235\,
            in1 => \N__21887\,
            in2 => \N__24623\,
            in3 => \N__27835\,
            lcout => OPEN,
            ltout => \POWERLED.N_449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRT5H5_8_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__22351\,
            in1 => \N__32842\,
            in2 => \N__21881\,
            in3 => \N__32672\,
            lcout => \POWERLED.dutycycle_RNIRT5H5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_13_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24114\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_2376_i\,
            ltout => \POWERLED.N_2376_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_12_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24443\,
            in1 => \N__24875\,
            in2 => \N__21872\,
            in3 => \N__23036\,
            lcout => \POWERLED.N_612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIG4L3G_0_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21950\,
            in1 => \N__21944\,
            in2 => \_gnd_net_\,
            in3 => \N__23483\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => \POWERLED.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_1_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21869\,
            in3 => \N__23392\,
            lcout => \POWERLED.count_off_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIFNOIG_5_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21989\,
            in1 => \N__21970\,
            in2 => \_gnd_net_\,
            in3 => \N__23485\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => \POWERLED.count_offZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_1_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21920\,
            in1 => \N__22037\,
            in2 => \N__21953\,
            in3 => \N__23391\,
            lcout => \POWERLED.un34_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__26132\,
            in1 => \_gnd_net_\,
            in2 => \N__22091\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32265\,
            ce => \N__23518\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIEAAR6_0_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22085\,
            in2 => \_gnd_net_\,
            in3 => \N__26131\,
            lcout => \POWERLED.count_off_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21928\,
            lcout => \POWERLED.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32265\,
            ce => \N__23518\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI9ELIG_2_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__23484\,
            in1 => \N__21938\,
            in2 => \N__21932\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22138\,
            lcout => \POWERLED.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32279\,
            ce => \N__23489\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDRHFG_13_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21899\,
            in1 => \N__21907\,
            in2 => \_gnd_net_\,
            in3 => \N__23487\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21908\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32279\,
            ce => \N__23489\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIFUIFG_14_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22145\,
            in1 => \N__22153\,
            in2 => \_gnd_net_\,
            in3 => \N__23488\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22154\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32279\,
            ce => \N__23489\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIH1KFG_15_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22139\,
            in1 => \N__22130\,
            in2 => \_gnd_net_\,
            in3 => \N__23490\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => \POWERLED.count_offZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_15_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22118\,
            in1 => \N__22106\,
            in2 => \N__22094\,
            in3 => \N__22089\,
            lcout => \POWERLED.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHQPIG_6_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22064\,
            in1 => \N__23486\,
            in2 => \_gnd_net_\,
            in3 => \N__22048\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22025\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22013\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22001\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22229\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22214\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22205\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22196\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22181\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22166\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_0_0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__30736\,
            in1 => \N__30414\,
            in2 => \N__22252\,
            in3 => \N__28847\,
            lcout => OPEN,
            ltout => \POWERLED.N_673_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIE48E2_1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__22160\,
            in1 => \N__23657\,
            in2 => \N__22163\,
            in3 => \N__30075\,
            lcout => \POWERLED.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_11_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__30737\,
            in1 => \N__30415\,
            in2 => \N__22253\,
            in3 => \N__26745\,
            lcout => \POWERLED.N_423_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23656\,
            in2 => \_gnd_net_\,
            in3 => \N__22521\,
            lcout => \clk_100Khz_signalkeep_3_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__30738\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30416\,
            lcout => \N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__23678\,
            in1 => \N__22271\,
            in2 => \N__33084\,
            in3 => \N__22265\,
            lcout => \POWERLED.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28832\,
            in2 => \_gnd_net_\,
            in3 => \N__30049\,
            lcout => \POWERLED.N_633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_5_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29231\,
            lcout => \POWERLED.un1_dutycycle_164_0_a3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27151\,
            in3 => \N__30412\,
            lcout => v5s_enn,
            ltout => \v5s_enn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_19_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__30727\,
            in1 => \N__25578\,
            in2 => \N__22274\,
            in3 => \N__22503\,
            lcout => \POWERLED.func_state_en_0_0\,
            ltout => \POWERLED.func_state_en_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6BR4J_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__22264\,
            in1 => \N__33063\,
            in2 => \N__22256\,
            in3 => \N__23677\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_m1_e_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__30413\,
            in1 => \_gnd_net_\,
            in2 => \N__22251\,
            in3 => \N__30735\,
            lcout => \POWERLED.dutycycle_N_3_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_rep1_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__25579\,
            in1 => \N__22522\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \clk_100Khz_signalkeep_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIU8AB2_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__22388\,
            in1 => \N__32768\,
            in2 => \N__25873\,
            in3 => \N__26280\,
            lcout => \POWERLED.func_state_1_m0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI7LSV8_0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__31590\,
            in1 => \N__26240\,
            in2 => \N__32667\,
            in3 => \N__22358\,
            lcout => \POWERLED.func_state_RNI7LSV8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5SKJ1_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110010"
        )
    port map (
            in0 => \N__29654\,
            in1 => \N__29558\,
            in2 => \N__29743\,
            in3 => \N__28925\,
            lcout => \POWERLED.func_state_RNI5SKJ1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25864\,
            in2 => \_gnd_net_\,
            in3 => \N__29980\,
            lcout => \POWERLED.N_617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22332\,
            in2 => \_gnd_net_\,
            in3 => \N__33077\,
            lcout => \N_626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26425\,
            lcout => \func_state_RNI_2_0\,
            ltout => \func_state_RNI_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29981\,
            in1 => \_gnd_net_\,
            in2 => \N__22283\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_215_i_0_o2_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__26746\,
            in1 => \N__26366\,
            in2 => \N__27582\,
            in3 => \N__25577\,
            lcout => \POWERLED.N_430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQHVM3_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22442\,
            in2 => \N__26015\,
            in3 => \N__22280\,
            lcout => \POWERLED.func_state_1_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30705\,
            in1 => \N__28791\,
            in2 => \N__30409\,
            in3 => \N__30012\,
            lcout => \POWERLED.dutycycle_1_0_iv_i_0_a2_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__27625\,
            in1 => \N__30708\,
            in2 => \_gnd_net_\,
            in3 => \N__30387\,
            lcout => \POWERLED.N_443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_0_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30706\,
            in1 => \N__28790\,
            in2 => \N__30410\,
            in3 => \N__27624\,
            lcout => \POWERLED.N_540_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIP4521_1_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111111"
        )
    port map (
            in0 => \N__30013\,
            in1 => \N__22436\,
            in2 => \N__23831\,
            in3 => \N__29267\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m2s2_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNINDFD3_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__32744\,
            in1 => \N__22430\,
            in2 => \N__22415\,
            in3 => \N__26276\,
            lcout => \POWERLED.N_74\,
            ltout => \POWERLED.N_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI4TUGC_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011101111"
        )
    port map (
            in0 => \N__22373\,
            in1 => \N__22412\,
            in2 => \N__22406\,
            in3 => \N__22403\,
            lcout => \POWERLED.func_state_1_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIGCDO1_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__30707\,
            in1 => \N__22387\,
            in2 => \N__30411\,
            in3 => \N__26275\,
            lcout => \POWERLED.N_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIFBNT_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__26029\,
            in1 => \_gnd_net_\,
            in2 => \N__23885\,
            in3 => \N__27861\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_i_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__26742\,
            in1 => \N__22367\,
            in2 => \N__22361\,
            in3 => \N__25582\,
            lcout => \POWERLED.N_71\,
            ltout => \POWERLED.N_71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVSVI5_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__22574\,
            in1 => \N__22558\,
            in2 => \N__22598\,
            in3 => \N__32626\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => \POWERLED.dutycycleZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22595\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32913\,
            in2 => \_gnd_net_\,
            in3 => \N__30018\,
            lcout => OPEN,
            ltout => \POWERLED.N_426_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIIASA2_2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111111"
        )
    port map (
            in0 => \N__29572\,
            in1 => \N__32783\,
            in2 => \N__22577\,
            in3 => \N__29489\,
            lcout => \POWERLED.dutycycle_eena_1\,
            ltout => \POWERLED.dutycycle_eena_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__22568\,
            in1 => \N__22559\,
            in2 => \N__22562\,
            in3 => \N__32627\,
            lcout => \POWERLED.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32450\,
            ce => 'H',
            sr => \N__31754\
        );

    \POWERLED.G_141_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25581\,
            in2 => \_gnd_net_\,
            in3 => \N__22523\,
            lcout => \G_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_7_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__22460\,
            in1 => \N__26771\,
            in2 => \N__32628\,
            in3 => \N__22454\,
            lcout => \POWERLED.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32412\,
            ce => 'H',
            sr => \N__31731\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23861\,
            in1 => \N__27234\,
            in2 => \N__30721\,
            in3 => \N__27623\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0\,
            ltout => \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNICSH47_7_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__32575\,
            in1 => \N__22453\,
            in2 => \N__22445\,
            in3 => \N__26770\,
            lcout => \POWERLED.dutycycleZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_5_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__30672\,
            in1 => \N__30288\,
            in2 => \_gnd_net_\,
            in3 => \N__27621\,
            lcout => \POWERLED.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_2_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27622\,
            in1 => \N__30671\,
            in2 => \N__30314\,
            in3 => \N__28816\,
            lcout => \POWERLED.func_state_RNIBVNS_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22721\,
            in3 => \N__22712\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22763\,
            in3 => \N__22700\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25195\,
            in2 => \N__22697\,
            in3 => \N__22679\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25183\,
            in2 => \N__22676\,
            in3 => \N__22652\,
            lcout => \POWERLED.mult1_un47_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_5\,
            carryout => \POWERLED.mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22649\,
            in3 => \N__22640\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => \POWERLED.mult1_un54_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22619\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__22869\,
            in1 => \N__22870\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__26552\,
            in1 => \N__30925\,
            in2 => \_gnd_net_\,
            in3 => \N__31400\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__31401\,
            in1 => \_gnd_net_\,
            in2 => \N__27098\,
            in3 => \N__31013\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNIZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_8_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__31298\,
            in1 => \N__31406\,
            in2 => \N__22838\,
            in3 => \N__24607\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011000110"
        )
    port map (
            in0 => \N__30926\,
            in1 => \N__31297\,
            in2 => \N__31430\,
            in3 => \N__32953\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31014\,
            in1 => \N__31405\,
            in2 => \_gnd_net_\,
            in3 => \N__27073\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22817\,
            in3 => \N__22785\,
            lcout => \POWERLED.mult1_un47_sum_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30927\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_7_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__27074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30144\,
            lcout => \POWERLED.N_510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRPVQ5_13_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__24062\,
            in1 => \N__22915\,
            in2 => \N__22934\,
            in3 => \N__31566\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31567\,
            in1 => \N__24061\,
            in2 => \N__22919\,
            in3 => \N__22930\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32466\,
            ce => 'H',
            sr => \N__31721\
        );

    \POWERLED.dutycycle_9_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__23849\,
            in1 => \N__27248\,
            in2 => \N__22889\,
            in3 => \N__31568\,
            lcout => \POWERLED.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32466\,
            ce => 'H',
            sr => \N__31721\
        );

    \POWERLED.dutycycle_RNI_1_10_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24796\,
            lcout => \POWERLED.un1_dutycycle_53_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_8_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27345\,
            in2 => \N__24618\,
            in3 => \N__24860\,
            lcout => \POWERLED.un1_dutycycle_53_40_0\,
            ltout => \POWERLED.un1_dutycycle_53_40_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_13_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111100"
        )
    port map (
            in0 => \N__24111\,
            in1 => \N__22907\,
            in2 => \N__22901\,
            in3 => \N__24473\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITR8L6_9_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__23848\,
            in1 => \N__27247\,
            in2 => \N__22888\,
            in3 => \N__31565\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => \POWERLED.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_8_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__27065\,
            in1 => \_gnd_net_\,
            in2 => \N__22874\,
            in3 => \N__24599\,
            lcout => \POWERLED.un1_dutycycle_53_31_a5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_8_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001000"
        )
    port map (
            in0 => \N__31020\,
            in1 => \N__31425\,
            in2 => \N__27106\,
            in3 => \N__24604\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_8\,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__27341\,
            in1 => \_gnd_net_\,
            in2 => \N__22994\,
            in3 => \N__31149\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNIZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_7_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__27096\,
            in1 => \N__31148\,
            in2 => \N__22991\,
            in3 => \N__24794\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_5_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27342\,
            in1 => \N__31150\,
            in2 => \N__31322\,
            in3 => \N__22982\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24425\,
            in1 => \N__31424\,
            in2 => \_gnd_net_\,
            in3 => \N__27340\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_31_a4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_6_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011011"
        )
    port map (
            in0 => \N__31147\,
            in1 => \N__22958\,
            in2 => \N__22967\,
            in3 => \N__22964\,
            lcout => \POWERLED.un1_dutycycle_53_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_8_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31019\,
            in1 => \N__31423\,
            in2 => \N__27105\,
            in3 => \N__24603\,
            lcout => \POWERLED.un1_dutycycle_53_31_a0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__27343\,
            in1 => \N__26963\,
            in2 => \N__24368\,
            in3 => \N__24608\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITTAN6_14_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__22942\,
            in1 => \N__27913\,
            in2 => \N__23960\,
            in3 => \N__31583\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__31585\,
            in1 => \N__23956\,
            in2 => \N__27917\,
            in3 => \N__22943\,
            lcout => \POWERLED.dutycycleZ1Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32472\,
            ce => 'H',
            sr => \N__31781\
        );

    \POWERLED.dutycycle_15_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__27962\,
            in1 => \N__31586\,
            in2 => \N__23054\,
            in3 => \N__23935\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32472\,
            ce => 'H',
            sr => \N__31781\
        );

    \POWERLED.dutycycle_RNI_12_8_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__24866\,
            in1 => \N__24332\,
            in2 => \N__24542\,
            in3 => \N__24472\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_12Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__27512\,
            in1 => \N__26952\,
            in2 => \N__23066\,
            in3 => \N__24677\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIV0CN6_15_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__31584\,
            in1 => \N__23050\,
            in2 => \N__23936\,
            in3 => \N__27961\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => \POWERLED.dutycycleZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_15_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23042\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_2381_i\,
            ltout => \POWERLED.N_2381_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_14_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24678\,
            in1 => \N__27754\,
            in2 => \N__23039\,
            in3 => \N__29335\,
            lcout => \POWERLED.un2_count_clk_17_0_0_a2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__23009\,
            in1 => \N__23020\,
            in2 => \N__31592\,
            in3 => \N__24137\,
            lcout => \POWERLED.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32479\,
            ce => 'H',
            sr => \N__31750\
        );

    \POWERLED.dutycycle_RNI_13_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001011010"
        )
    port map (
            in0 => \N__24113\,
            in1 => \N__27755\,
            in2 => \N__23108\,
            in3 => \N__24449\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFDK47_11_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__24136\,
            in1 => \N__31575\,
            in2 => \N__23021\,
            in3 => \N__23008\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => \POWERLED.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_11_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23114\,
            in3 => \N__24767\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_12_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__24348\,
            in1 => \N__26978\,
            in2 => \N__23111\,
            in3 => \N__24442\,
            lcout => \POWERLED.un1_dutycycle_53_2_1\,
            ltout => \POWERLED.un1_dutycycle_53_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_13_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__24112\,
            in1 => \N__24349\,
            in2 => \N__23099\,
            in3 => \N__24364\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24980\,
            in1 => \N__25052\,
            in2 => \N__25523\,
            in3 => \N__25070\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23078\,
            in1 => \N__23084\,
            in2 => \N__23087\,
            in3 => \N__23072\,
            lcout => \VPP_VDDQ_un6_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24998\,
            in1 => \N__25016\,
            in2 => \N__24962\,
            in3 => \N__25034\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__25544\,
            in1 => \N__24509\,
            in2 => \N__25499\,
            in3 => \N__24941\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25223\,
            in1 => \N__25454\,
            in2 => \N__25103\,
            in3 => \N__25475\,
            lcout => \VPP_VDDQ.un6_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIMTB22_0_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__23339\,
            in1 => \N__23289\,
            in2 => \_gnd_net_\,
            in3 => \N__23251\,
            lcout => \VPP_VDDQ.N_64_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000111010"
        )
    port map (
            in0 => \N__23254\,
            in1 => \N__23360\,
            in2 => \N__23302\,
            in3 => \N__23341\,
            lcout => \VPP_VDDQ_curr_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32280\,
            ce => \N__25316\,
            sr => \_gnd_net_\
        );

    \POWERLED.G_30_0_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__23252\,
            in1 => \N__23338\,
            in2 => \N__23301\,
            in3 => \N__25400\,
            lcout => OPEN,
            ltout => \POWERLED.G_30Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_30_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__23297\,
            in1 => \N__23253\,
            in2 => \N__23363\,
            in3 => \N__23359\,
            lcout => \G_30\,
            ltout => \G_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23348\,
            in3 => \N__25401\,
            lcout => \VPP_VDDQ.N_92_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__23340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23296\,
            lcout => \VPP_VDDQ_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32280\,
            ce => \N__25316\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23224\,
            lcout => \POWERLED.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32269\,
            ce => \N__23519\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIBHMIG_3_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23234\,
            in1 => \N__23511\,
            in2 => \N__23228\,
            in3 => \N__26097\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => \POWERLED.count_offZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_3_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23198\,
            in1 => \N__23602\,
            in2 => \N__23174\,
            in3 => \N__23171\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_10_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23144\,
            in1 => \N__23138\,
            in2 => \N__23126\,
            in3 => \N__23123\,
            lcout => \POWERLED.count_off_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDKNIG_4_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__26098\,
            in1 => \N__23570\,
            in2 => \N__23539\,
            in3 => \N__23588\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23587\,
            in2 => \_gnd_net_\,
            in3 => \N__26101\,
            lcout => \POWERLED.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32269\,
            ce => \N__23519\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23563\,
            lcout => \POWERLED.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32269\,
            ce => \N__23519\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIH5L3G_1_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__23564\,
            in1 => \N__23552\,
            in2 => \N__23540\,
            in3 => \N__26096\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S3n_RNI5DLR_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111111111"
        )
    port map (
            in0 => \N__30354\,
            in1 => \N__30734\,
            in2 => \_gnd_net_\,
            in3 => \N__28850\,
            lcout => OPEN,
            ltout => \N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNI8TRB2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011110010"
        )
    port map (
            in0 => \N__26734\,
            in1 => \N__26342\,
            in2 => \N__23372\,
            in3 => \N__23655\,
            lcout => OPEN,
            ltout => \N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep2_RNIDD505_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110011"
        )
    port map (
            in0 => \N__29893\,
            in1 => \N__23627\,
            in2 => \N__23369\,
            in3 => \N__30118\,
            lcout => \POWERLED_g2_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_5_1_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__30733\,
            in1 => \N__30353\,
            in2 => \N__26754\,
            in3 => \N__27177\,
            lcout => OPEN,
            ltout => \POWERLED.g0_5Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIA2VR1_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__25580\,
            in1 => \N__25866\,
            in2 => \N__23366\,
            in3 => \N__28849\,
            lcout => OPEN,
            ltout => \POWERLED.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIUKM0G_1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000111011"
        )
    port map (
            in0 => \N__23699\,
            in1 => \N__23693\,
            in2 => \N__23681\,
            in3 => \N__23663\,
            lcout => \POWERLED.func_state_1_m2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIGN2N5_1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__23669\,
            in1 => \N__25867\,
            in2 => \N__23639\,
            in3 => \N__23786\,
            lcout => \POWERLED.func_state_1_m2_N_3_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_17_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__26735\,
            in1 => \N__23654\,
            in2 => \N__26365\,
            in3 => \N__27176\,
            lcout => \POWERLED.N_671_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S3n_RNI5DLR_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30352\,
            in2 => \N__26239\,
            in3 => \N__30732\,
            lcout => OPEN,
            ltout => \G_7_i_a4_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep1_RNI75Q52_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__27172\,
            in1 => \N__26285\,
            in2 => \N__23630\,
            in3 => \N__26349\,
            lcout => \RSMRST_PWRGD.G_7_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPGQN2_4_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28133\,
            in2 => \_gnd_net_\,
            in3 => \N__28112\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_0_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26231\,
            lcout => \POWERLED.N_533\,
            ltout => \POWERLED.N_533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI98AF2_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23612\,
            in2 => \N__23621\,
            in3 => \N__27171\,
            lcout => \POWERLED.un1_clk_100khz_51_and_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIA70J1_1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__23618\,
            in1 => \N__29655\,
            in2 => \N__30377\,
            in3 => \N__29726\,
            lcout => \POWERLED.un1_clk_100khz_51_and_i_3_0_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOI5P1_0_5_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__23747\,
            in1 => \N__29423\,
            in2 => \N__25969\,
            in3 => \N__25934\,
            lcout => \POWERLED.un1_dutycycle_172_m3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25865\,
            in2 => \_gnd_net_\,
            in3 => \N__30115\,
            lcout => \POWERLED.func_state_RNI_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI1TUN2_7_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29099\,
            in1 => \N__23720\,
            in2 => \_gnd_net_\,
            in3 => \N__28264\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => \POWERLED.count_clkZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__30116\,
            in1 => \N__23728\,
            in2 => \N__23741\,
            in3 => \N__28624\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPGQN2_7_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23729\,
            in1 => \N__28300\,
            in2 => \N__28628\,
            in3 => \N__26281\,
            lcout => \POWERLED.N_490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_7_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32385\,
            ce => \N__29117\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_5_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__31308\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30117\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIV0AS_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000101"
        )
    port map (
            in0 => \N__29536\,
            in1 => \N__23819\,
            in2 => \N__23714\,
            in3 => \N__29408\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_52_and_i_0_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIGV3L6_5_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__23711\,
            in1 => \N__23774\,
            in2 => \N__23702\,
            in3 => \N__29537\,
            lcout => OPEN,
            ltout => \POWERLED.N_448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIS28SB_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__23768\,
            in1 => \N__32740\,
            in2 => \N__23789\,
            in3 => \N__32593\,
            lcout => \POWERLED.func_state_RNIS28SBZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__30696\,
            in1 => \N__27173\,
            in2 => \N__30347\,
            in3 => \N__26230\,
            lcout => \POWERLED.N_656_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__31589\,
            in1 => \N__28801\,
            in2 => \_gnd_net_\,
            in3 => \N__31306\,
            lcout => OPEN,
            ltout => \POWERLED.N_133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQAA33_0_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23815\,
            in1 => \_gnd_net_\,
            in2 => \N__23777\,
            in3 => \N__23756\,
            lcout => \POWERLED.un1_dutycycle_172_m4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIO5723_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111111"
        )
    port map (
            in0 => \N__29699\,
            in1 => \N__29573\,
            in2 => \N__29668\,
            in3 => \N__32745\,
            lcout => \POWERLED.dutycycle_eena_14_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30318\,
            in1 => \N__30709\,
            in2 => \N__32956\,
            in3 => \N__27174\,
            lcout => OPEN,
            ltout => \POWERLED.N_488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQAA33_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__25946\,
            in1 => \N__26627\,
            in2 => \N__23759\,
            in3 => \N__31305\,
            lcout => \POWERLED.un1_dutycycle_172_m2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_0_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__28800\,
            in1 => \N__30061\,
            in2 => \N__30346\,
            in3 => \N__28923\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_30_and_i_0_0_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIV0AS_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__28924\,
            in1 => \_gnd_net_\,
            in2 => \N__23750\,
            in3 => \N__27175\,
            lcout => \POWERLED.N_91_1_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_5_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31145\,
            in1 => \N__29355\,
            in2 => \N__31307\,
            in3 => \N__30781\,
            lcout => \POWERLED.func_state_1_m2s2_i_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_8_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27227\,
            lcout => \POWERLED.func_state_RNI_8Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_6_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29274\,
            lcout => \POWERLED.N_435_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI02AS_0_1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30694\,
            in1 => \N__28841\,
            in2 => \N__27185\,
            in3 => \N__27228\,
            lcout => \POWERLED.count_off_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30928\,
            in1 => \N__29275\,
            in2 => \N__29230\,
            in3 => \N__26553\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_96_0_a3_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__26623\,
            in1 => \N__31024\,
            in2 => \N__23822\,
            in3 => \N__31432\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30695\,
            in2 => \_gnd_net_\,
            in3 => \N__26755\,
            lcout => \POWERLED.N_251\,
            ltout => \POWERLED.N_251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_10_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000100010"
        )
    port map (
            in0 => \N__30317\,
            in1 => \N__24793\,
            in2 => \N__23804\,
            in3 => \N__29892\,
            lcout => \POWERLED.N_506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26547\,
            in3 => \N__30905\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__26578\,
            in1 => \N__24029\,
            in2 => \N__30924\,
            in3 => \N__23792\,
            lcout => \POWERLED.g0_i_m2_rn_1_0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24010\,
            in2 => \N__32940\,
            in3 => \N__23876\,
            lcout => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31018\,
            in2 => \N__24036\,
            in3 => \N__23873\,
            lcout => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31431\,
            in2 => \N__24042\,
            in3 => \N__23870\,
            lcout => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31310\,
            in2 => \N__24038\,
            in3 => \N__23867\,
            lcout => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_4\,
            carryout => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24014\,
            in2 => \N__31146\,
            in3 => \N__23864\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27075\,
            in2 => \N__24037\,
            in3 => \N__23855\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24619\,
            in2 => \N__24044\,
            in3 => \N__23852\,
            lcout => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27354\,
            in2 => \N__24039\,
            in3 => \N__23837\,
            lcout => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_8\,
            carryout => \POWERLED.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24022\,
            in2 => \N__24814\,
            in3 => \N__23834\,
            lcout => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_9\,
            carryout => \POWERLED.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24705\,
            in2 => \N__24040\,
            in3 => \N__24122\,
            lcout => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_10\,
            carryout => \POWERLED.un1_dutycycle_94_cry_11_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24021\,
            in2 => \N__26977\,
            in3 => \N__24119\,
            lcout => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_11_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24116\,
            in2 => \N__24041\,
            in3 => \N__24047\,
            lcout => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_12\,
            carryout => \POWERLED.un1_dutycycle_94_cry_13_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27770\,
            in2 => \N__24043\,
            in3 => \N__23942\,
            lcout => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_13_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__27524\,
            in1 => \_gnd_net_\,
            in2 => \N__29294\,
            in3 => \N__23939\,
            lcout => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.VCCST_EN_i_1_i_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27672\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30666\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIP1UT_4_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101010101"
        )
    port map (
            in0 => \N__24222\,
            in1 => \N__31564\,
            in2 => \N__23900\,
            in3 => \N__32607\,
            lcout => \POWERLED.dutycycle_RNIP1UTZ0Z_4\,
            ltout => \POWERLED.dutycycle_RNIP1UTZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIDH8E6_4_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001101"
        )
    port map (
            in0 => \N__32834\,
            in1 => \N__24223\,
            in2 => \N__23888\,
            in3 => \N__24239\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => \POWERLED.dutycycleZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31122\,
            in2 => \N__24242\,
            in3 => \N__27355\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIF86R3_4_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27932\,
            in1 => \N__26900\,
            in2 => \N__27457\,
            in3 => \N__29812\,
            lcout => \POWERLED.dutycycle_RNIF86R3Z0Z_4\,
            ltout => \POWERLED.dutycycle_RNIF86R3Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101000110011"
        )
    port map (
            in0 => \N__24224\,
            in1 => \N__24233\,
            in2 => \N__24227\,
            in3 => \N__32835\,
            lcout => \POWERLED.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32419\,
            ce => 'H',
            sr => \N__31757\
        );

    \POWERLED.dutycycle_8_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__24164\,
            in1 => \N__24175\,
            in2 => \N__31563\,
            in3 => \N__24188\,
            lcout => \POWERLED.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32449\,
            ce => 'H',
            sr => \N__31771\
        );

    \POWERLED.dutycycle_RNI_3_8_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111010"
        )
    port map (
            in0 => \N__24606\,
            in1 => \_gnd_net_\,
            in2 => \N__27097\,
            in3 => \N__31144\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_31_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_11_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__24143\,
            in1 => \N__24706\,
            in2 => \N__24212\,
            in3 => \N__24209\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRNTO5_8_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__24187\,
            in1 => \N__31508\,
            in2 => \N__24179\,
            in3 => \N__24163\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => \POWERLED.dutycycleZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_8_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24149\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_10_8\,
            ltout => \POWERLED.dutycycle_RNI_10_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_8_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__24605\,
            in1 => \N__24320\,
            in2 => \N__24146\,
            in3 => \N__24326\,
            lcout => \POWERLED.un1_dutycycle_53_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_7_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111000000"
        )
    port map (
            in0 => \N__27364\,
            in1 => \N__31399\,
            in2 => \N__31154\,
            in3 => \N__27066\,
            lcout => \POWERLED.un1_dutycycle_53_9_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_3_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110100000"
        )
    port map (
            in0 => \N__31398\,
            in1 => \N__31023\,
            in2 => \N__27371\,
            in3 => \N__31140\,
            lcout => \POWERLED.un1_dutycycle_53_9_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__31580\,
            in1 => \N__24298\,
            in2 => \N__26996\,
            in3 => \N__24314\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32463\,
            ce => 'H',
            sr => \N__31767\
        );

    \POWERLED.dutycycle_RNIHGL47_12_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26992\,
            in1 => \N__24313\,
            in2 => \N__24299\,
            in3 => \N__31579\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => \POWERLED.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_12_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24284\,
            in3 => \N__24778\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_9_a0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_8_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__24427\,
            in1 => \N__24468\,
            in2 => \N__24281\,
            in3 => \N__24830\,
            lcout => \POWERLED.un1_dutycycle_53_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_14_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27743\,
            in2 => \_gnd_net_\,
            in3 => \N__24700\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_11_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_10_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111010010"
        )
    port map (
            in0 => \N__24777\,
            in1 => \N__24266\,
            in2 => \N__24260\,
            in3 => \N__24491\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_14_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24257\,
            in3 => \N__27744\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__27344\,
            in1 => \N__24426\,
            in2 => \N__24795\,
            in3 => \N__24467\,
            lcout => \POWERLED.un1_dutycycle_53_45_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__31151\,
            in1 => \N__31421\,
            in2 => \N__27375\,
            in3 => \N__27085\,
            lcout => \POWERLED.un1_dutycycle_53_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_8_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__31422\,
            in1 => \N__31152\,
            in2 => \N__27104\,
            in3 => \N__24612\,
            lcout => \POWERLED.un1_dutycycle_53_35_1\,
            ltout => \POWERLED.un1_dutycycle_53_35_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_7_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__27359\,
            in1 => \N__24485\,
            in2 => \N__24476\,
            in3 => \N__27089\,
            lcout => \POWERLED.un1_dutycycle_53_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_6_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__24386\,
            in1 => \N__24858\,
            in2 => \N__24353\,
            in3 => \N__24377\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_6_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__31153\,
            in1 => \_gnd_net_\,
            in2 => \N__27376\,
            in3 => \N__24434\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_6\,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_6_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24856\,
            in2 => \N__24380\,
            in3 => \N__24376\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_11_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__27360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24676\,
            lcout => \POWERLED.un1_dutycycle_53_50_a0_0\,
            ltout => \POWERLED.un1_dutycycle_53_50_a0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_11_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24857\,
            in2 => \N__24335\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_53_50_a0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__24919\,
            in1 => \N__24904\,
            in2 => \N__24890\,
            in3 => \N__31582\,
            lcout => \POWERLED.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32480\,
            ce => 'H',
            sr => \N__31780\
        );

    \POWERLED.dutycycle_RNI6P2N6_10_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__31581\,
            in1 => \N__24920\,
            in2 => \N__24908\,
            in3 => \N__24886\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => \POWERLED.dutycycleZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_12_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__27370\,
            in1 => \_gnd_net_\,
            in2 => \N__24878\,
            in3 => \N__26969\,
            lcout => \POWERLED.un2_count_clk_17_0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__24748\,
            in1 => \N__27368\,
            in2 => \_gnd_net_\,
            in3 => \N__24696\,
            lcout => \POWERLED.un1_dutycycle_53_50_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_12_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110101000"
        )
    port map (
            in0 => \N__24695\,
            in1 => \N__24747\,
            in2 => \N__27377\,
            in3 => \N__26968\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_10_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_8_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__24859\,
            in1 => \N__24821\,
            in2 => \N__24833\,
            in3 => \N__24613\,
            lcout => \POWERLED.un1_dutycycle_53_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_12_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24746\,
            in2 => \_gnd_net_\,
            in3 => \N__26967\,
            lcout => \POWERLED.un1_dutycycle_53_9_a1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__24749\,
            in1 => \N__27369\,
            in2 => \N__24707\,
            in3 => \N__24614\,
            lcout => \POWERLED.un1_dutycycle_53_50_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25418\,
            in1 => \N__24508\,
            in2 => \N__24533\,
            in3 => \N__24532\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_1_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25404\,
            in1 => \N__25069\,
            in2 => \_gnd_net_\,
            in3 => \N__25055\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_2_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25419\,
            in1 => \N__25051\,
            in2 => \_gnd_net_\,
            in3 => \N__25037\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_3_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25405\,
            in1 => \N__25033\,
            in2 => \_gnd_net_\,
            in3 => \N__25019\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_4_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25420\,
            in1 => \N__25015\,
            in2 => \_gnd_net_\,
            in3 => \N__25001\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_5_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25406\,
            in1 => \N__24997\,
            in2 => \_gnd_net_\,
            in3 => \N__24983\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_6_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25421\,
            in1 => \N__24979\,
            in2 => \_gnd_net_\,
            in3 => \N__24965\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_7_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25407\,
            in1 => \N__24958\,
            in2 => \_gnd_net_\,
            in3 => \N__24944\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__32332\,
            ce => 'H',
            sr => \N__25801\
        );

    \VPP_VDDQ.count_8_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25433\,
            in1 => \N__24940\,
            in2 => \_gnd_net_\,
            in3 => \N__24923\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__32333\,
            ce => 'H',
            sr => \N__25800\
        );

    \VPP_VDDQ.count_9_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25417\,
            in1 => \N__25543\,
            in2 => \_gnd_net_\,
            in3 => \N__25526\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__32333\,
            ce => 'H',
            sr => \N__25800\
        );

    \VPP_VDDQ.count_10_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25430\,
            in1 => \N__25516\,
            in2 => \_gnd_net_\,
            in3 => \N__25502\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__32333\,
            ce => 'H',
            sr => \N__25800\
        );

    \VPP_VDDQ.count_11_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25415\,
            in1 => \N__25492\,
            in2 => \_gnd_net_\,
            in3 => \N__25478\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__32333\,
            ce => 'H',
            sr => \N__25800\
        );

    \VPP_VDDQ.count_12_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25431\,
            in1 => \N__25471\,
            in2 => \_gnd_net_\,
            in3 => \N__25457\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__32333\,
            ce => 'H',
            sr => \N__25800\
        );

    \VPP_VDDQ.count_13_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25416\,
            in1 => \N__25450\,
            in2 => \_gnd_net_\,
            in3 => \N__25436\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__32333\,
            ce => 'H',
            sr => \N__25800\
        );

    \VPP_VDDQ.count_14_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25432\,
            in1 => \N__25222\,
            in2 => \_gnd_net_\,
            in3 => \N__25205\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__32333\,
            ce => 'H',
            sr => \N__25800\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25180\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25096\,
            in2 => \_gnd_net_\,
            in3 => \N__25106\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32342\,
            ce => \N__25082\,
            sr => \N__25805\
        );

    \POWERLED.count_clk_RNIRJRN2_4_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25775\,
            in1 => \N__29060\,
            in2 => \_gnd_net_\,
            in3 => \N__28393\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_4_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32334\,
            ce => \N__29103\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNITMSN2_5_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25769\,
            in1 => \N__29061\,
            in2 => \_gnd_net_\,
            in3 => \N__28357\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_5_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32334\,
            ce => \N__29103\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIVPTN2_6_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25763\,
            in1 => \N__29062\,
            in2 => \_gnd_net_\,
            in3 => \N__28330\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_6_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28331\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32334\,
            ce => \N__29103\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIH9TE_10_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__26707\,
            in1 => \N__25634\,
            in2 => \_gnd_net_\,
            in3 => \N__25872\,
            lcout => \POWERLED.count_off_RNIH9TEZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8AQH_0_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__25586\,
            in1 => \N__28848\,
            in2 => \_gnd_net_\,
            in3 => \N__26708\,
            lcout => \POWERLED.func_state_RNI8AQHZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINH2G2_11_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__28168\,
            in1 => \N__29039\,
            in2 => \N__25886\,
            in3 => \N__28520\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__28071\,
            in1 => \_gnd_net_\,
            in2 => \N__28546\,
            in3 => \N__28714\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI118L2_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25892\,
            in2 => \N__25898\,
            in3 => \N__29038\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => \POWERLED.count_clkZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28522\,
            in1 => \_gnd_net_\,
            in2 => \N__25895\,
            in3 => \N__28716\,
            lcout => \POWERLED.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32423\,
            ce => \N__29118\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_0_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28717\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28516\,
            lcout => \POWERLED.count_clk_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_11_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28521\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28169\,
            lcout => \POWERLED.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32423\,
            ce => \N__29118\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28523\,
            lcout => \POWERLED.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32423\,
            ce => \N__29118\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__28070\,
            in1 => \N__28377\,
            in2 => \N__28652\,
            in3 => \N__28209\,
            lcout => \POWERLED.count_clk_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30157\,
            in2 => \_gnd_net_\,
            in3 => \N__25871\,
            lcout => \POWERLED.func_state_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__28382\,
            in1 => \N__28310\,
            in2 => \N__28076\,
            in3 => \N__28214\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPGQN2_3_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__28132\,
            in1 => \_gnd_net_\,
            in2 => \N__25808\,
            in3 => \N__28648\,
            lcout => \POWERLED.N_668\,
            ltout => \POWERLED.N_668_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNILPF34_3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__26010\,
            in1 => \N__26384\,
            in2 => \N__26147\,
            in3 => \N__27644\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIEAAR6_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011101100"
        )
    port map (
            in0 => \N__26454\,
            in1 => \N__26144\,
            in2 => \N__26135\,
            in3 => \N__30153\,
            lcout => \POWERLED.N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2VV9A_0_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__26386\,
            in1 => \N__26033\,
            in2 => \N__26014\,
            in3 => \N__26300\,
            lcout => \POWERLED.func_state_RNI2VV9A_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101010111"
        )
    port map (
            in0 => \N__26455\,
            in1 => \N__25978\,
            in2 => \N__25921\,
            in3 => \N__30152\,
            lcout => \POWERLED.un1_func_state25_6_0_0_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNINEAB6_1_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__25979\,
            in1 => \N__28088\,
            in2 => \N__30158\,
            in3 => \N__26385\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOI5P1_5_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111000000"
        )
    port map (
            in0 => \N__25970\,
            in1 => \N__29180\,
            in2 => \N__26180\,
            in3 => \N__31247\,
            lcout => \POWERLED.un1_dutycycle_172_m0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111110101"
        )
    port map (
            in0 => \N__31248\,
            in1 => \N__32954\,
            in2 => \N__29312\,
            in3 => \N__28843\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOGRS_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111000001"
        )
    port map (
            in0 => \N__26175\,
            in1 => \N__29308\,
            in2 => \N__25937\,
            in3 => \N__31587\,
            lcout => \POWERLED.un1_dutycycle_172_m1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001111"
        )
    port map (
            in0 => \N__26294\,
            in1 => \N__26709\,
            in2 => \N__25922\,
            in3 => \N__28844\,
            lcout => \POWERLED.count_clk_en_917_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__28842\,
            in1 => \N__26456\,
            in2 => \N__26390\,
            in3 => \N__30105\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI19L28_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26606\,
            in1 => \N__26309\,
            in2 => \N__26303\,
            in3 => \N__28597\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26293\,
            lcout => \func_state_RNI_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__26174\,
            in2 => \N__30145\,
            in3 => \N__26540\,
            lcout => \POWERLED.dutycycle_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__26192\,
            in1 => \N__30799\,
            in2 => \N__26459\,
            in3 => \N__30782\,
            lcout => \POWERLED.N_676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30783\,
            in1 => \N__26453\,
            in2 => \_gnd_net_\,
            in3 => \N__26191\,
            lcout => \func_state_RNI_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31276\,
            in1 => \N__31090\,
            in2 => \N__30920\,
            in3 => \N__26508\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_0\,
            ltout => \POWERLED.dutycycle_RNI_4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOGRS_0_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111111111"
        )
    port map (
            in0 => \N__29395\,
            in1 => \N__30784\,
            in2 => \N__26183\,
            in3 => \N__26179\,
            lcout => \POWERLED.un1_count_off_1_sqmuxa_8_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29456\,
            in1 => \N__31089\,
            in2 => \N__30919\,
            in3 => \N__26509\,
            lcout => OPEN,
            ltout => \POWERLED.N_546_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__29396\,
            in1 => \N__30839\,
            in2 => \N__26630\,
            in3 => \N__29292\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__29222\,
            in1 => \N__30728\,
            in2 => \N__30284\,
            in3 => \N__30079\,
            lcout => \POWERLED.N_482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIG2F54_1_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__32640\,
            in1 => \N__26396\,
            in2 => \N__26588\,
            in3 => \N__26600\,
            lcout => \POWERLED.g0_i_m2_rn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE0E38_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__26405\,
            in1 => \_gnd_net_\,
            in2 => \N__26471\,
            in3 => \N__26446\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => \POWERLED.dutycycleZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIIASA2_1_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111101"
        )
    port map (
            in0 => \N__32793\,
            in1 => \N__29604\,
            in2 => \N__26591\,
            in3 => \N__29485\,
            lcout => \POWERLED.dutycycle_eena_0_0\,
            ltout => \POWERLED.dutycycle_eena_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIUTUT3_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26579\,
            in1 => \N__30143\,
            in2 => \N__26564\,
            in3 => \N__32639\,
            lcout => \POWERLED.g0_i_m2_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIIASA2_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111101"
        )
    port map (
            in0 => \N__32792\,
            in1 => \N__26522\,
            in2 => \N__29618\,
            in3 => \N__29484\,
            lcout => \POWERLED.dutycycle_eena\,
            ltout => \POWERLED.dutycycle_eena_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIP8K44_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__26870\,
            in1 => \N__26851\,
            in2 => \N__26561\,
            in3 => \N__32638\,
            lcout => \POWERLED.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26470\,
            in2 => \N__26458\,
            in3 => \N__26404\,
            lcout => \POWERLED.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32462\,
            ce => 'H',
            sr => \N__31772\
        );

    \POWERLED.dutycycle_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__26869\,
            in1 => \N__26858\,
            in2 => \N__32668\,
            in3 => \N__26852\,
            lcout => \POWERLED.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32462\,
            ce => 'H',
            sr => \N__31772\
        );

    \POWERLED.dutycycle_RNI2MQD_7_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__30243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27099\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_36_and_i_0_a2_c_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI7JPT2_7_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26786\,
            in1 => \N__26843\,
            in2 => \N__26831\,
            in3 => \N__27451\,
            lcout => \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26828\,
            in2 => \_gnd_net_\,
            in3 => \N__29619\,
            lcout => \VCCIN_PWRGD.un10_outputZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_m1_0_a2_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001000000"
        )
    port map (
            in0 => \N__30580\,
            in1 => \N__30244\,
            in2 => \N__29912\,
            in3 => \N__26744\,
            lcout => \POWERLED.un1_clk_100khz_36_and_i_0_a2_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI99TE_7_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__27666\,
            in1 => \N__30578\,
            in2 => \N__27107\,
            in3 => \N__27891\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI48JN5_7_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__32811\,
            in1 => \N__26780\,
            in2 => \N__26774\,
            in3 => \N__29805\,
            lcout => \POWERLED.dutycycle_eena_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_43_and_i_0_o2_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__26743\,
            in1 => \N__30579\,
            in2 => \_gnd_net_\,
            in3 => \N__29900\,
            lcout => OPEN,
            ltout => \POWERLED.N_249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_4_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100101010"
        )
    port map (
            in0 => \N__30258\,
            in1 => \N__31435\,
            in2 => \N__26633\,
            in3 => \N__30123\,
            lcout => \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30265\,
            in3 => \N__30146\,
            lcout => \POWERLED.func_state_RNI2MQDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI12AS_6_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__29898\,
            in1 => \_gnd_net_\,
            in2 => \N__29223\,
            in3 => \N__30670\,
            lcout => \POWERLED.N_203\,
            ltout => \POWERLED.N_203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI12AS_0_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26888\,
            in3 => \N__27879\,
            lcout => \POWERLED.N_531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000001010"
        )
    port map (
            in0 => \N__30239\,
            in1 => \N__29744\,
            in2 => \N__31022\,
            in3 => \N__29899\,
            lcout => OPEN,
            ltout => \POWERLED.N_521_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5TUF2_3_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__27442\,
            in1 => \N__31003\,
            in2 => \N__26885\,
            in3 => \N__30147\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_43_and_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRUFD6_3_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__26879\,
            in1 => \N__32826\,
            in2 => \N__26882\,
            in3 => \N__32645\,
            lcout => \POWERLED.dutycycle_en_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_3_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001010"
        )
    port map (
            in0 => \N__27880\,
            in1 => \N__31002\,
            in2 => \N__27825\,
            in3 => \N__33129\,
            lcout => \POWERLED.N_523\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_9_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000001010000"
        )
    port map (
            in0 => \N__27374\,
            in1 => \N__29914\,
            in2 => \N__30264\,
            in3 => \N__29748\,
            lcout => OPEN,
            ltout => \POWERLED.N_503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5TUF2_9_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__30122\,
            in1 => \N__27373\,
            in2 => \N__26873\,
            in3 => \N__27456\,
            lcout => \POWERLED.dutycycle_eena_2_0_0_tz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI12AS_9_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__27372\,
            in1 => \N__29913\,
            in2 => \_gnd_net_\,
            in3 => \N__30720\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_30_and_i_0_a2_5_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_9_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101110"
        )
    port map (
            in0 => \N__27206\,
            in1 => \N__27810\,
            in2 => \N__27260\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_2_d_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRUFD6_9_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100000000"
        )
    port map (
            in0 => \N__27257\,
            in1 => \N__32827\,
            in2 => \N__27251\,
            in3 => \N__32646\,
            lcout => \POWERLED.dutycycle_RNIRUFD6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI02AS_1_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__30687\,
            in1 => \N__27205\,
            in2 => \_gnd_net_\,
            in3 => \N__27184\,
            lcout => \POWERLED.N_421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_3_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__31434\,
            in1 => \N__27103\,
            in2 => \_gnd_net_\,
            in3 => \N__31021\,
            lcout => \POWERLED.N_604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_12_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__26974\,
            in1 => \N__33130\,
            in2 => \N__27901\,
            in3 => \N__27819\,
            lcout => OPEN,
            ltout => \POWERLED.N_520_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRUFD6_12_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__26906\,
            in1 => \N__32831\,
            in2 => \N__26999\,
            in3 => \N__32669\,
            lcout => \POWERLED.dutycycle_RNIRUFD6Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_12_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__26976\,
            in1 => \N__30235\,
            in2 => \N__29759\,
            in3 => \N__29915\,
            lcout => OPEN,
            ltout => \POWERLED.N_518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5TUF2_12_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__30149\,
            in1 => \N__26975\,
            in2 => \N__26909\,
            in3 => \N__27458\,
            lcout => \POWERLED.un1_clk_100khz_42_and_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI99TE_4_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__27893\,
            in1 => \N__31433\,
            in2 => \N__30665\,
            in3 => \N__27673\,
            lcout => \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_14_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__27767\,
            in1 => \N__33128\,
            in2 => \N__27902\,
            in3 => \N__27832\,
            lcout => OPEN,
            ltout => \POWERLED.N_526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI36306_14_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__27698\,
            in1 => \N__32832\,
            in2 => \N__27920\,
            in3 => \N__32670\,
            lcout => \POWERLED.dutycycle_RNI36306Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24KO1_15_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__27897\,
            in1 => \N__33127\,
            in2 => \N__27476\,
            in3 => \N__27831\,
            lcout => \POWERLED.N_529\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE3861_14_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__30227\,
            in1 => \N__29757\,
            in2 => \N__27687\,
            in3 => \N__27769\,
            lcout => OPEN,
            ltout => \POWERLED.N_524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNID4I22_14_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27768\,
            in1 => \N__27459\,
            in2 => \N__27701\,
            in3 => \N__30150\,
            lcout => \POWERLED.un1_clk_100khz_47_and_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE3861_15_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__30228\,
            in1 => \N__29758\,
            in2 => \N__27688\,
            in3 => \N__27520\,
            lcout => OPEN,
            ltout => \POWERLED.N_527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNID4I22_1_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__27475\,
            in1 => \N__27460\,
            in2 => \N__27383\,
            in3 => \N__30151\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_48_and_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI36306_1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__32671\,
            in1 => \N__32833\,
            in2 => \N__27380\,
            in3 => \N__27968\,
            lcout => \POWERLED.dutycycle_en_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI300O2_8_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29080\,
            in1 => \N__27950\,
            in2 => \_gnd_net_\,
            in3 => \N__28228\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_8_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28229\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32261\,
            ce => \N__29106\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_15_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28463\,
            lcout => \POWERLED.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32261\,
            ce => \N__29106\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI531O2_9_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29081\,
            in1 => \N__27944\,
            in2 => \_gnd_net_\,
            in3 => \N__28189\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_9_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28190\,
            lcout => \POWERLED.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32261\,
            ce => \N__29106\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINDPN2_2_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27938\,
            in2 => \N__29104\,
            in3 => \N__28027\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_2_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32261\,
            ce => \N__29106\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_3_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32309\,
            ce => \N__29076\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPGQN2_3_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28147\,
            in1 => \N__29082\,
            in2 => \_gnd_net_\,
            in3 => \N__28002\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => \POWERLED.count_clkZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_3_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__28044\,
            in1 => \N__27987\,
            in2 => \N__28154\,
            in3 => \N__28245\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_6_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__28345\,
            in1 => \N__28314\,
            in2 => \N__28151\,
            in3 => \N__28110\,
            lcout => \POWERLED.count_clk_RNIZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPGQN2_0_3_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__28003\,
            in1 => \N__28148\,
            in2 => \N__29105\,
            in3 => \N__28246\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPGQN2_1_3_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__28346\,
            in1 => \N__27988\,
            in2 => \N__28136\,
            in3 => \N__28045\,
            lcout => \POWERLED.N_625\,
            ltout => \POWERLED.N_625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPGQN2_5_3_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__28111\,
            in1 => \_gnd_net_\,
            in2 => \N__28091\,
            in3 => \N__28319\,
            lcout => \POWERLED.count_clk_RNIPGQN2_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28721\,
            in2 => \N__28075\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28547\,
            in1 => \_gnd_net_\,
            in2 => \N__28049\,
            in3 => \N__28016\,
            lcout => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_1\,
            carryout => \POWERLED.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28551\,
            in1 => \_gnd_net_\,
            in2 => \N__28013\,
            in3 => \N__27992\,
            lcout => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_2\,
            carryout => \POWERLED.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28548\,
            in1 => \_gnd_net_\,
            in2 => \N__27989\,
            in3 => \N__28385\,
            lcout => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_3\,
            carryout => \POWERLED.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28552\,
            in1 => \_gnd_net_\,
            in2 => \N__28381\,
            in3 => \N__28349\,
            lcout => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_4\,
            carryout => \POWERLED.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28549\,
            in1 => \N__28344\,
            in2 => \_gnd_net_\,
            in3 => \N__28322\,
            lcout => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_5\,
            carryout => \POWERLED.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28553\,
            in1 => \_gnd_net_\,
            in2 => \N__28318\,
            in3 => \N__28250\,
            lcout => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_6\,
            carryout => \POWERLED.un1_count_clk_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28550\,
            in1 => \N__28247\,
            in2 => \_gnd_net_\,
            in3 => \N__28217\,
            lcout => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_7\,
            carryout => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28540\,
            in1 => \N__28213\,
            in2 => \_gnd_net_\,
            in3 => \N__28175\,
            lcout => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28543\,
            in1 => \N__28406\,
            in2 => \_gnd_net_\,
            in3 => \N__28172\,
            lcout => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_9\,
            carryout => \POWERLED.un1_count_clk_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28672\,
            in2 => \_gnd_net_\,
            in3 => \N__28160\,
            lcout => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_10\,
            carryout => \POWERLED.un1_count_clk_2_cry_11_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28544\,
            in1 => \_gnd_net_\,
            in2 => \N__28571\,
            in3 => \N__28157\,
            lcout => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_11_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28541\,
            in1 => \N__29144\,
            in2 => \_gnd_net_\,
            in3 => \N__28559\,
            lcout => \POWERLED.count_clk_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_12\,
            carryout => \POWERLED.un1_count_clk_2_cry_13_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_13_c_RNITQ5G2_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28545\,
            in1 => \N__28400\,
            in2 => \_gnd_net_\,
            in3 => \N__28556\,
            lcout => \POWERLED.count_clk_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_13_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28542\,
            in1 => \N__28448\,
            in2 => \_gnd_net_\,
            in3 => \N__28475\,
            lcout => \POWERLED.count_clk_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIVT6G2_15_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29075\,
            in1 => \N__28472\,
            in2 => \_gnd_net_\,
            in3 => \N__28459\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIECHG2_10_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__28436\,
            in1 => \N__28414\,
            in2 => \N__29119\,
            in3 => \N__28447\,
            lcout => \POWERLED.un2_count_clk_17_0_o2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28429\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32380\,
            ce => \N__29110\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIECHG2_0_10_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28991\,
            in1 => \N__28428\,
            in2 => \_gnd_net_\,
            in3 => \N__28415\,
            lcout => \POWERLED.un1_count_clk_2_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_14_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28695\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32380\,
            ce => \N__29110\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNILKND2_0_14_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28696\,
            in1 => \_gnd_net_\,
            in2 => \N__29120\,
            in3 => \N__28681\,
            lcout => \POWERLED.un1_count_clk_2_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI008L2_0_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28733\,
            in1 => \N__28990\,
            in2 => \_gnd_net_\,
            in3 => \N__28727\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => \POWERLED.count_clkZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNILKND2_14_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111000"
        )
    port map (
            in0 => \N__28697\,
            in1 => \N__29074\,
            in2 => \N__28685\,
            in3 => \N__28682\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_o2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNISLCE7_10_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28673\,
            in1 => \N__28931\,
            in2 => \N__28661\,
            in3 => \N__28658\,
            lcout => \POWERLED.count_clk_RNISLCE7Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5SKJ1_0_1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__30740\,
            in1 => \N__29608\,
            in2 => \N__28637\,
            in3 => \N__28892\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6GV92_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__28623\,
            in1 => \N__32644\,
            in2 => \N__28601\,
            in3 => \N__28598\,
            lcout => \POWERLED.count_clk_en\,
            ltout => \POWERLED.count_clk_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPK3G2_0_12_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29134\,
            in1 => \_gnd_net_\,
            in2 => \N__28574\,
            in3 => \N__28939\,
            lcout => \POWERLED.un1_count_clk_2_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_12_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29133\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32407\,
            ce => \N__29069\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_13_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29161\,
            lcout => \POWERLED.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32407\,
            ce => \N__29069\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIRN4G2_13_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29162\,
            in1 => \N__29150\,
            in2 => \_gnd_net_\,
            in3 => \N__29070\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => \POWERLED.count_clkZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPK3G2_12_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111000"
        )
    port map (
            in0 => \N__29135\,
            in1 => \N__29037\,
            in2 => \N__28943\,
            in3 => \N__28940\,
            lcout => \POWERLED.un2_count_clk_17_0_o2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_0_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28908\,
            lcout => \POWERLED.N_492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__28874\,
            in1 => \N__28885\,
            in2 => \N__32836\,
            in3 => \N__30434\,
            lcout => \POWERLED.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32465\,
            ce => 'H',
            sr => \N__31756\
        );

    \POWERLED.dutycycle_RNIKVDEF_5_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110000"
        )
    port map (
            in0 => \N__30433\,
            in1 => \N__32821\,
            in2 => \N__28886\,
            in3 => \N__28873\,
            lcout => \POWERLED.dutycycleZ1Z_5\,
            ltout => \POWERLED.dutycycleZ1Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_5_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29369\,
            in1 => \N__31105\,
            in2 => \N__28859\,
            in3 => \N__28845\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_5\,
            ltout => \POWERLED.dutycycle_RNI_3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__30785\,
            in1 => \_gnd_net_\,
            in2 => \N__28856\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011011111"
        )
    port map (
            in0 => \N__29173\,
            in1 => \N__31591\,
            in2 => \N__28853\,
            in3 => \N__28846\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_8Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__28739\,
            in1 => \N__30835\,
            in2 => \N__29762\,
            in3 => \N__29293\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_RNIOGRSZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNITCGG2_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111101110"
        )
    port map (
            in0 => \N__29725\,
            in1 => \N__29669\,
            in2 => \N__29633\,
            in3 => \N__29600\,
            lcout => \POWERLED.N_413_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101110011111100"
        )
    port map (
            in0 => \N__30812\,
            in1 => \N__29470\,
            in2 => \N__32492\,
            in3 => \N__32815\,
            lcout => \POWERLED.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32461\,
            ce => 'H',
            sr => \N__31755\
        );

    \POWERLED.dutycycle_RNIQCMNB_6_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110000"
        )
    port map (
            in0 => \N__32814\,
            in1 => \N__30811\,
            in2 => \N__29471\,
            in3 => \N__32488\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => \POWERLED.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_6_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__29364\,
            in1 => \_gnd_net_\,
            in2 => \N__29459\,
            in3 => \N__29455\,
            lcout => \POWERLED.N_672\,
            ltout => \POWERLED.N_672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_6_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29389\,
            in1 => \_gnd_net_\,
            in2 => \N__29411\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_168_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_6_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29388\,
            lcout => \POWERLED.N_412_i\,
            ltout => \POWERLED.N_412_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_3_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29365\,
            in2 => \N__29339\,
            in3 => \N__29336\,
            lcout => \POWERLED.dutycycle_RNI_6Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_5_1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__29291\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29209\,
            lcout => \POWERLED.func_state_RNI_5Z0Z_1\,
            ltout => \POWERLED.func_state_RNI_5Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_9_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30842\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_23_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIJM2T1_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100011"
        )
    port map (
            in0 => \N__30469\,
            in1 => \N__30824\,
            in2 => \N__30316\,
            in3 => \N__30442\,
            lcout => \POWERLED.N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI12AS_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__30598\,
            in1 => \N__29896\,
            in2 => \_gnd_net_\,
            in3 => \N__30124\,
            lcout => \POWERLED.func_state_RNI12ASZ0Z_1\,
            ltout => \POWERLED.func_state_RNI12ASZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI12AS_5_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__30803\,
            in1 => \_gnd_net_\,
            in2 => \N__30788\,
            in3 => \N__30769\,
            lcout => \POWERLED.dutycycle_eena_13_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI12AS_6_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__31088\,
            in1 => \N__30125\,
            in2 => \N__30664\,
            in3 => \N__29895\,
            lcout => \POWERLED.N_530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIIK1T1_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100011"
        )
    port map (
            in0 => \N__30470\,
            in1 => \N__30455\,
            in2 => \N__30315\,
            in3 => \N__30443\,
            lcout => \POWERLED.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI01AS_6_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31087\,
            in1 => \N__30289\,
            in2 => \N__30148\,
            in3 => \N__29897\,
            lcout => OPEN,
            ltout => \POWERLED.N_532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBD845_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29813\,
            in1 => \N__29789\,
            in2 => \N__29771\,
            in3 => \N__29768\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_51_and_i_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI0DF58_5_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__32849\,
            in1 => \N__32825\,
            in2 => \N__32678\,
            in3 => \N__32637\,
            lcout => \POWERLED.dutycycle_RNI0DF58Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__31498\,
            in1 => \N__31603\,
            in2 => \N__31637\,
            in3 => \N__31622\,
            lcout => \POWERLED.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32464\,
            ce => 'H',
            sr => \N__31773\
        );

    \POWERLED.dutycycle_RNIH92L6_3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__31633\,
            in1 => \N__31621\,
            in2 => \N__31604\,
            in3 => \N__31497\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => \POWERLED.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31103\,
            in2 => \N__31442\,
            in3 => \N__32944\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_5_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011110000"
        )
    port map (
            in0 => \N__31263\,
            in1 => \N__31426\,
            in2 => \N__31439\,
            in3 => \N__30917\,
            lcout => \POWERLED.un1_dutycycle_53_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_3_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__31104\,
            in1 => \N__30982\,
            in2 => \N__31436\,
            in3 => \N__30918\,
            lcout => OPEN,
            ltout => \POWERLED.un1_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_5_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__31264\,
            in1 => \N__30848\,
            in2 => \N__31190\,
            in3 => \N__31187\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_3_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__31102\,
            in1 => \N__30981\,
            in2 => \_gnd_net_\,
            in3 => \N__30916\,
            lcout => \POWERLED.d_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNISQ2V_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__33161\,
            in1 => \N__33123\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33020\,
            in1 => \N__33002\,
            in2 => \N__32987\,
            in3 => \N__32975\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_2_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32948\,
            in2 => \_gnd_net_\,
            in3 => \N__32864\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
