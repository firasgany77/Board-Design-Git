-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 7 2022 11:04:43

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : out std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \DSW_PWRGD.un1_curr_state10_0\ : std_logic;
signal v33dsw_ok : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\ : std_logic;
signal \G_27\ : std_logic;
signal \G_27_cascade_\ : std_logic;
signal \DSW_PWRGD.N_27_1\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_7_l_fx\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_4_l_fx\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_14_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_RNIZ0Z_1\ : std_logic;
signal \PCH_PWRGD.count_RNIZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_1\ : std_logic;
signal \DSW_PWRGD.countZ0Z_3\ : std_logic;
signal \DSW_PWRGD.countZ0Z_4\ : std_logic;
signal \DSW_PWRGD.countZ0Z_0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_1\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0_cascade_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_11\ : std_logic;
signal \DSW_PWRGD.countZ0Z_10\ : std_logic;
signal \DSW_PWRGD.countZ0Z_6\ : std_logic;
signal \DSW_PWRGD.countZ0Z_5\ : std_logic;
signal \DSW_PWRGD.countZ0Z_9\ : std_logic;
signal \DSW_PWRGD.countZ0Z_7\ : std_logic;
signal \DSW_PWRGD.countZ0Z_8\ : std_logic;
signal \DSW_PWRGD.countZ0Z_2\ : std_logic;
signal \PCH_PWRGD.N_2126_i_cascade_\ : std_logic;
signal \PCH_PWRGD.N_381_cascade_\ : std_logic;
signal \PCH_PWRGD.N_254_0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_12\ : std_logic;
signal \DSW_PWRGD.countZ0Z_13\ : std_logic;
signal \DSW_PWRGD.countZ0Z_14\ : std_logic;
signal \DSW_PWRGD.countZ0Z_15\ : std_logic;
signal \DSW_PWRGD.un4_count_11\ : std_logic;
signal \DSW_PWRGD.un4_count_10\ : std_logic;
signal \DSW_PWRGD.un4_count_8_cascade_\ : std_logic;
signal \DSW_PWRGD.un4_count_9\ : std_logic;
signal \DSW_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.N_381\ : std_logic;
signal \PCH_PWRGD.N_2126_i\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.N_255_0_cascade_\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \bfn_2_5_0_\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_cry_0_i\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \POWERLED.N_4527_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_0\ : std_logic;
signal \POWERLED.N_4528_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_1\ : std_logic;
signal \POWERLED.un85_clk_100khz_3\ : std_logic;
signal \POWERLED.N_4529_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_2\ : std_logic;
signal \POWERLED.un85_clk_100khz_4\ : std_logic;
signal \POWERLED.N_4530_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_3\ : std_logic;
signal \POWERLED.N_4531_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_4\ : std_logic;
signal \POWERLED.un85_clk_100khz_6\ : std_logic;
signal \POWERLED.N_4532_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_5\ : std_logic;
signal \POWERLED.N_4533_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_7\ : std_logic;
signal \POWERLED.N_4534_i\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \POWERLED.N_4535_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_8\ : std_logic;
signal \POWERLED.N_4536_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_9\ : std_logic;
signal \POWERLED.N_4537_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_10\ : std_logic;
signal \POWERLED.N_4538_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_11\ : std_logic;
signal \POWERLED.N_4539_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_12\ : std_logic;
signal \POWERLED.N_4540_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_13\ : std_logic;
signal \POWERLED.N_4541_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_14\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \POWERLED.un85_clk_100khz_1\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_9\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_11\ : std_logic;
signal v33a_enn : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_13\ : std_logic;
signal \POWERLED.un85_clk_100khz_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_7\ : std_logic;
signal \POWERLED.un85_clk_100khz_12\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_14\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.m4_0_0_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_6\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0\ : std_logic;
signal \PCH_PWRGD.curr_state_0_0\ : std_logic;
signal \PCH_PWRGD.count_rst_11\ : std_logic;
signal \PCH_PWRGD.count_rst_11_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_3_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.count_rst_10_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \PCH_PWRGD.count_rst_3_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_11_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_3\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_7\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_4_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_5\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_13_cascade_\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.N_1_i_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_7_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_8\ : std_logic;
signal \PCH_PWRGD.count_0_14\ : std_logic;
signal \PCH_PWRGD.count_0_13\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \N_187_cascade_\ : std_logic;
signal v33a_ok : std_logic;
signal v5a_ok : std_logic;
signal slp_susn : std_logic;
signal v1p8a_ok : std_logic;
signal \rsmrst_pwrgd_signal_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal v5s_enn : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2121\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_0\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_2\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_a2_5_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_46_0_cascade_\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \POWERLED.mult1_un47_sum_i\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_5_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_6\ : std_logic;
signal \PCH_PWRGD.count_rst_9\ : std_logic;
signal \PCH_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.count_rst_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.count_rst_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.count_rst\ : std_logic;
signal \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\ : std_logic;
signal \PCH_PWRGD.N_386\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_rst_5\ : std_logic;
signal \RSMRST_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_1_i\ : std_logic;
signal \RSMRST_PWRGD.un4_count_8\ : std_logic;
signal \RSMRST_PWRGD.un4_count_10\ : std_logic;
signal \RSMRST_PWRGD.un4_count_11\ : std_logic;
signal \POWERLED.g0_i_o3_0_cascade_\ : std_logic;
signal \POWERLED.pwm_outZ0\ : std_logic;
signal \POWERLED.g0_i_o3_0\ : std_logic;
signal pwrbtn_led : std_logic;
signal \POWERLED.curr_state_3_0_cascade_\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \POWERLED.count_RNIZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_8\ : std_logic;
signal \PCH_PWRGD.count_0_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_10\ : std_logic;
signal \RSMRST_PWRGD_curr_state_0\ : std_logic;
signal \N_187\ : std_logic;
signal \G_11_cascade_\ : std_logic;
signal \POWERLED.count_0_4\ : std_logic;
signal \POWERLED.count_0_2\ : std_logic;
signal \POWERLED.count_0_11\ : std_logic;
signal \POWERLED.count_0_3\ : std_logic;
signal \POWERLED.count_0_15\ : std_logic;
signal \POWERLED.count_0_7\ : std_logic;
signal \POWERLED.count_0_8\ : std_logic;
signal \POWERLED.count_0_10\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_0_cZ0\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_1_cZ0\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_2_cZ0\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_3_cZ0\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_4_cZ0\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_5_cZ0\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_7_cZ0\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_8_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_9_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_11\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2_c\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_c\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_c\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_c\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_c\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSCZ0\ : std_logic;
signal \PCH_PWRGD.count_0_2\ : std_logic;
signal \PCH_PWRGD.count_rst_12_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_3\ : std_logic;
signal \PCH_PWRGD.count_0_12\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.count_0_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_2\ : std_logic;
signal \RSMRST_PWRGD.N_256_i\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.N_27_2\ : std_logic;
signal \G_11\ : std_logic;
signal \POWERLED.un79_clk_100khzlto4_0_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlt15_0_cascade_\ : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_5\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_6_cascade_\ : std_logic;
signal \POWERLED.count_RNIZ0Z_15_cascade_\ : std_logic;
signal \POWERLED.N_8\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_cry_1_c_RNIBZ0Z209\ : std_logic;
signal \POWERLED.un1_count_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_cry_2_c_RNICZ0Z419\ : std_logic;
signal \POWERLED.un1_count_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\ : std_logic;
signal \POWERLED.un1_count_cry_3\ : std_logic;
signal \POWERLED.un1_count_cry_4\ : std_logic;
signal \POWERLED.un1_count_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59\ : std_logic;
signal \POWERLED.un1_count_cry_6\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69\ : std_logic;
signal \POWERLED.un1_count_cry_7\ : std_logic;
signal \POWERLED.un1_count_cry_8\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\ : std_logic;
signal \POWERLED.un1_count_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7\ : std_logic;
signal \POWERLED.un1_count_cry_10\ : std_logic;
signal \POWERLED.un1_count_cry_11\ : std_logic;
signal \POWERLED.un1_count_cry_12\ : std_logic;
signal \POWERLED.un1_count_cry_13\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.un1_count_cry_14\ : std_logic;
signal \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\ : std_logic;
signal \POWERLED.count_0_9\ : std_logic;
signal \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_eena_1_cascade_\ : std_logic;
signal \POWERLED.N_108_f0_1\ : std_logic;
signal \POWERLED.N_108_f0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_0\ : std_logic;
signal \POWERLED.dutycycle_eena_0_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_1\ : std_logic;
signal \POWERLED.dutycycle_eena_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_2\ : std_logic;
signal \POWERLED.func_state_0_sqmuxa_0_o2_xZ0Z1_cascade_\ : std_logic;
signal \POWERLED.g1_1_cascade_\ : std_logic;
signal \POWERLED.N_300_N_0_cascade_\ : std_logic;
signal \POWERLED.N_4548_0\ : std_logic;
signal \POWERLED.N_217_N_0\ : std_logic;
signal \POWERLED.N_353_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_14\ : std_logic;
signal \POWERLED.N_86_f0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_11\ : std_logic;
signal \POWERLED.dutycycle_en_11_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_15\ : std_logic;
signal \POWERLED.N_2215_i\ : std_logic;
signal \POWERLED.N_84_f0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_10_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ1Z_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.mult1_un47_sum\ : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_29\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_4_sf\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.dutycycle_en_12\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.dutycycle_RNI_11Z0Z_7_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_45_a0_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_45_a0_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_1\ : std_logic;
signal \HDA_STRAP.N_14_cascade_\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal hda_sdo_atp : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD_delayed_vccin_ok\ : std_logic;
signal \HDA_STRAP.curr_state_RNO_0Z0Z_0\ : std_logic;
signal \HDA_STRAP.N_5_0\ : std_logic;
signal \POWERLED.N_341_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_a3_1_0_2_cascade_\ : std_logic;
signal \POWERLED.N_64\ : std_logic;
signal \POWERLED.g0_0_a3_1_cascade_\ : std_logic;
signal \POWERLED.g0_3_1\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_2\ : std_logic;
signal \POWERLED.func_state_RNIMQ0FZ0Z_1\ : std_logic;
signal \POWERLED.N_309\ : std_logic;
signal \POWERLED.func_state_1_m0_1_cascade_\ : std_logic;
signal \POWERLED.count_RNI_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.func_state_RNIG5G37Z0Z_1\ : std_logic;
signal \POWERLED.func_state_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_1\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7\ : std_logic;
signal \POWERLED.count_0_13\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\ : std_logic;
signal \POWERLED.count_0_5\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\ : std_logic;
signal \POWERLED.count_0_14\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49\ : std_logic;
signal \POWERLED.count_0_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11_cascade_\ : std_logic;
signal \POWERLED.N_148_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_10\ : std_logic;
signal \POWERLED.dutycycle_en_10_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.un1_func_state25_4_i_a2_1\ : std_logic;
signal \POWERLED.N_301_cascade_\ : std_logic;
signal \POWERLED.N_341\ : std_logic;
signal \POWERLED.count_clk_en_1_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIBVNS_1Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_ns_1\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\ : std_logic;
signal \POWERLED.N_171\ : std_logic;
signal \POWERLED.N_283\ : std_logic;
signal \POWERLED.N_275_0\ : std_logic;
signal \POWERLED.dutycycle_set_0_0\ : std_logic;
signal \POWERLED.dutycycle_eena_13_0\ : std_logic;
signal \POWERLED.dutycycle_set_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_0_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_0\ : std_logic;
signal \POWERLED.d_i3_mux_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_13_4_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_13_4_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_13_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_11\ : std_logic;
signal \POWERLED.g0_0_1\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\ : std_logic;
signal \POWERLED.g0_i_1_cascade_\ : std_logic;
signal \POWERLED.g0_i_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9\ : std_logic;
signal \POWERLED.dutycycle_rst_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.g0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_14\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIEB706Z0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ1Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNIEB706Z0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_d_0\ : std_logic;
signal \POWERLED.N_143_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\ : std_logic;
signal \POWERLED.dutycycleZ1Z_8\ : std_logic;
signal \HDA_STRAP.un4_count_12\ : std_logic;
signal \HDA_STRAP.un4_count_9_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_13\ : std_logic;
signal \HDA_STRAP.un4_count_11\ : std_logic;
signal \HDA_STRAP.un4_count_10\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal \HDA_STRAP.un4_count\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_0\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_1_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m0_0_1_0\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_11_cascade_\ : std_logic;
signal \POWERLED.N_310\ : std_logic;
signal \POWERLED.N_314_cascade_\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_11\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIHDGK3_0Z0Z_1\ : std_logic;
signal \POWERLED.N_67\ : std_logic;
signal \POWERLED.func_state_1_m0_0\ : std_logic;
signal \POWERLED.func_state_RNIHDGK3_0Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_287_N\ : std_logic;
signal \POWERLED.func_state_RNI_1Z0Z_0\ : std_logic;
signal \POWERLED.func_state_RNI_1Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIBK1UZ0Z_0\ : std_logic;
signal \POWERLED.N_326_0\ : std_logic;
signal \POWERLED.func_stateZ1Z_0\ : std_logic;
signal \POWERLED.func_state_RNIB74H7Z0Z_1\ : std_logic;
signal \POWERLED.func_state_RNI6RANZ0Z_1\ : std_logic;
signal \POWERLED.func_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\ : std_logic;
signal \POWERLED.N_275_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_48_and_i_o2_2_0_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_48_and_i_o2_3_0\ : std_logic;
signal \POWERLED.N_197\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7\ : std_logic;
signal \POWERLED.count_0_12\ : std_logic;
signal \POWERLED.count_clk_0_2\ : std_logic;
signal \POWERLED.count_clk_0_13\ : std_logic;
signal \POWERLED.count_clk_0_14\ : std_logic;
signal \POWERLED.count_clk_0_3\ : std_logic;
signal \POWERLED.count_clk_0_4\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_10Z0Z_0\ : std_logic;
signal \POWERLED.N_337\ : std_logic;
signal \SUSWARN_N_fast\ : std_logic;
signal \POWERLED.N_390_cascade_\ : std_logic;
signal \SUSWARN_N_rep1\ : std_logic;
signal \POWERLED.dutycycle_eena_3_0_0_sx_cascade_\ : std_logic;
signal slp_s3n : std_logic;
signal rsmrstn : std_logic;
signal \POWERLED.N_222\ : std_logic;
signal \POWERLED.un1_dutycycle_172_sm3\ : std_logic;
signal \POWERLED.un1_clk_100khz_52_and_i_m2_1\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m4_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_52_and_i_0Z0Z_0\ : std_logic;
signal \POWERLED.N_225_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_14_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_14\ : std_logic;
signal \POWERLED.dutycycle_set_1\ : std_logic;
signal \POWERLED.dutycycle_0_5\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\ : std_logic;
signal \POWERLED.dutycycleZ1Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_13_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_4_1\ : std_logic;
signal \POWERLED.dutycycle_en_8\ : std_logic;
signal \POWERLED.dutycycle_eena_3_0_1\ : std_logic;
signal \POWERLED.dutycycle_eena_3_d_0\ : std_logic;
signal \POWERLED.dutycycle_en_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_1_0_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_1_0\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_a2_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\ : std_logic;
signal \POWERLED.dutycycle_RNI4VJH7Z0Z_4\ : std_logic;
signal \POWERLED.dutycycleZ1Z_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.dutycycle_RNI_11Z0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_a0_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_11\ : std_logic;
signal \POWERLED.N_209_iZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_a7_0\ : std_logic;
signal \POWERLED.N_144_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_7\ : std_logic;
signal \POWERLED.count_clk_RNIBVNSZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_51_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_4\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_15\ : std_logic;
signal \POWERLED.func_state_RNIBVNSZ0Z_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_7\ : std_logic;
signal \POWERLED.N_8_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_3\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.g0_i_a6_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_12\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.func_state_RNIC4OR2Z0Z_0\ : std_logic;
signal \POWERLED.N_390\ : std_logic;
signal \POWERLED.N_209\ : std_logic;
signal \POWERLED.N_145_N_cascade_\ : std_logic;
signal \G_154\ : std_logic;
signal \POWERLED.dutycycle_en_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \HDA_STRAP.curr_state_RNIH91AZ0Z_1\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_0\ : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_1\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.countZ0Z_3\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.countZ0Z_5\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7\ : std_logic;
signal \HDA_STRAP.countZ0Z_8\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_8\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_9\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_8\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_10\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_13\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.countZ0Z_15\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_16\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_16\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_17\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_a2_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_305_N_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_1\ : std_logic;
signal \POWERLED.N_150_i\ : std_logic;
signal \POWERLED.N_154\ : std_logic;
signal \POWERLED.N_389\ : std_logic;
signal \POWERLED.count_off_0_10\ : std_logic;
signal \POWERLED.count_off_1_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_offZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_4_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \POWERLED.count_RNIZ0Z_15\ : std_logic;
signal \POWERLED.curr_state_1_0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.count_0_1\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i\ : std_logic;
signal \POWERLED.count_0_0\ : std_logic;
signal slp_s4n : std_logic;
signal \RSMRST_PWRGD_RSMRSTn_2_fast\ : std_logic;
signal \POWERLED.count_clk_0_5\ : std_logic;
signal \POWERLED.count_clk_0_6\ : std_logic;
signal \POWERLED.count_clk_0_8\ : std_logic;
signal \POWERLED.count_clk_0_9\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_15\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_7\ : std_logic;
signal \POWERLED.N_392\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \POWERLED.func_state_RNIBVNS_0Z0Z_0\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m4_bm_rn_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIMUFP1Z0Z_2\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \G_9\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m4_bm_sn\ : std_logic;
signal \POWERLED.N_20_i\ : std_logic;
signal \POWERLED.dutycycle_N_3_mux_0\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_2_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIBVNS_0Z0Z_1\ : std_logic;
signal \POWERLED.N_2171_i\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m3_ns_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_0\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m3\ : std_logic;
signal \POWERLED.N_2200_i\ : std_logic;
signal \POWERLED.un1_dutycycle_96_0_a3_1\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \POWERLED.N_327\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_3_1_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_2\ : std_logic;
signal \POWERLED.N_342\ : std_logic;
signal \POWERLED.N_155\ : std_logic;
signal \POWERLED.N_336\ : std_logic;
signal \POWERLED.dutycycle_RNI_9Z0Z_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.un1_i3_mux\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un6_count_8_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \VPP_VDDQ.un6_count_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \POWERLED.count_off_0_5\ : std_logic;
signal \POWERLED.count_off_0_15\ : std_logic;
signal \POWERLED.count_off_0_8\ : std_logic;
signal \POWERLED.un34_clk_100khz_0_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_12\ : std_logic;
signal \POWERLED.un34_clk_100khz_1\ : std_logic;
signal \POWERLED.count_off_1_6\ : std_logic;
signal \POWERLED.count_off_1_6_cascade_\ : std_logic;
signal \POWERLED.count_off_1_2\ : std_logic;
signal \POWERLED.count_off_1_2_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.count_off_1_7\ : std_logic;
signal \POWERLED.count_off_1_7_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_3\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_off_1_11\ : std_logic;
signal \POWERLED.count_off_1_11_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_0\ : std_logic;
signal \POWERLED.func_state_RNI_2Z0Z_1\ : std_logic;
signal \POWERLED.N_289_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIBVNS_2Z0Z_0\ : std_logic;
signal \POWERLED.count_off_RNIG5N6N1Z0Z_11\ : std_logic;
signal \POWERLED.func_state_RNI_5Z0Z_1\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_2_tz_0_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_2\ : std_logic;
signal \POWERLED.func_state_RNI_2Z0Z_0\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_304_N\ : std_logic;
signal \POWERLED.un1_N_3_mux_0\ : std_logic;
signal \POWERLED.func_state\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_2_0\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_3_0\ : std_logic;
signal \POWERLED.N_352_cascade_\ : std_logic;
signal \POWERLED.N_394\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\ : std_logic;
signal \POWERLED.N_2182_i\ : std_logic;
signal \POWERLED.N_352\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_2_2_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_9\ : std_logic;
signal \POWERLED.count_clk_0_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_4_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.count_clk_0_0\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_2\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_0\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_1_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_3\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.count_2_1_4\ : std_logic;
signal \VPP_VDDQ.count_2_1_5\ : std_logic;
signal \VPP_VDDQ.count_2_1_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\ : std_logic;
signal \VPP_VDDQ.count_2_1_13_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal vpp_en : std_logic;
signal vccst_en : std_logic;
signal \VPP_VDDQ.N_360_cascade_\ : std_logic;
signal \VPP_VDDQ.N_264_i\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ.curr_state_RNITROD7Z0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_RNITROD7Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_27_0\ : std_logic;
signal \VPP_VDDQ.N_382\ : std_logic;
signal \VPP_VDDQ.N_186\ : std_logic;
signal \VPP_VDDQ.N_214\ : std_logic;
signal \VPP_VDDQ.un6_count\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ.N_360\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_0\ : std_logic;
signal \N_27_g\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_off_0_12\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1\ : std_logic;
signal \POWERLED.count_off_0_1\ : std_logic;
signal \POWERLED.count_off_0_13\ : std_logic;
signal \POWERLED.count_offZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_11\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_axb_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1_c_RNIN70FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4_c_RNIQD3FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un3_count_off_1_axb_6\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un3_count_off_1_axb_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6_c_RNISH5FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7_c_RNITJ6FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8\ : std_logic;
signal \POWERLED.un3_count_off_1_axb_9\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8_c_RNIUL7FZ0\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9_c_RNIVN8FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9\ : std_logic;
signal \POWERLED.un3_count_off_1_axb_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10_c_RNI7ULDZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11_c_RNI80NDZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12_c_RNI92ODZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14_c_RNIB6QDZ0\ : std_logic;
signal \POWERLED.count_off_0_14\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.count_offZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\ : std_logic;
signal \POWERLED.count_off_1_3\ : std_logic;
signal \POWERLED.count_off_1_3_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.un3_count_off_1_axb_3\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.count_offZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_0_0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\ : std_logic;
signal \POWERLED.N_116\ : std_logic;
signal \POWERLED.count_off_0_4\ : std_logic;
signal \POWERLED.count_off_enZ0\ : std_logic;
signal v33s_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal slp_s3n_signal : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal v5s_ok : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\ : std_logic;
signal dsw_pwrok : std_logic;
signal vccin_en : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0_cascade_\ : std_logic;
signal pch_pwrok : std_logic;
signal vccst_pwrgd : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_0\ : std_logic;
signal \VPP_VDDQ.N_53\ : std_logic;
signal \VPP_VDDQ.N_53_i\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_11\ : std_logic;
signal \POWERLED.count_clk_0_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.func_state_RNICAC53_0_0\ : std_logic;
signal \POWERLED.count_clk_0_1\ : std_logic;
signal \POWERLED.count_clk_en\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.N_163\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.N_176\ : std_logic;
signal \VPP_VDDQ.N_47_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\ : std_logic;
signal \VPP_VDDQ.count_2_1_2\ : std_logic;
signal \VPP_VDDQ.count_2_1_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.N_385\ : std_logic;
signal \VPP_VDDQ.N_385_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.m4_0_cascade_\ : std_logic;
signal suswarn_n : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \N_579_g\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_6\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_1\ : std_logic;
signal vddq_ok : std_logic;
signal \N_362\ : std_logic;
signal \VPP_VDDQ.count_2_1_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_12\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_4_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_11\ : std_logic;
signal \VPP_VDDQ.N_1_i_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_1_7\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_7_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_12_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_14\ : std_logic;
signal \VPP_VDDQ.count_2_1_14_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_0_6\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_1_8\ : std_logic;
signal \VPP_VDDQ.count_2_1_11_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_1_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.count_2_1_10_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_10\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\ : std_logic;
signal \VPP_VDDQ.N_1_i\ : std_logic;
signal \VPP_VDDQ.count_2_0_12\ : std_logic;
signal fpga_osc : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    SLP_S0n <= \SLP_S0n_wire\;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    SUSWARN_N <= \SUSWARN_N_wire\;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34245\,
            DIN => \N__34244\,
            DOUT => \N__34243\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34245\,
            PADOUT => \N__34244\,
            PADIN => \N__34243\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34236\,
            DIN => \N__34235\,
            DOUT => \N__34234\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34236\,
            PADOUT => \N__34235\,
            PADIN => \N__34234\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15452\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34227\,
            DIN => \N__34226\,
            DOUT => \N__34225\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34227\,
            PADOUT => \N__34226\,
            PADIN => \N__34225\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16306\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34218\,
            DIN => \N__34217\,
            DOUT => \N__34216\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34218\,
            PADOUT => \N__34217\,
            PADIN => \N__34216\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15761\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34209\,
            DIN => \N__34208\,
            DOUT => \N__34207\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34209\,
            PADOUT => \N__34208\,
            PADIN => \N__34207\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34200\,
            DIN => \N__34199\,
            DOUT => \N__34198\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34200\,
            PADOUT => \N__34199\,
            PADIN => \N__34198\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34191\,
            DIN => \N__34190\,
            DOUT => \N__34189\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34191\,
            PADOUT => \N__34190\,
            PADIN => \N__34189\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34182\,
            DIN => \N__34181\,
            DOUT => \N__34180\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34182\,
            PADOUT => \N__34181\,
            PADIN => \N__34180\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34173\,
            DIN => \N__34172\,
            DOUT => \N__34171\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34173\,
            PADOUT => \N__34172\,
            PADIN => \N__34171\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16333\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34164\,
            DIN => \N__34163\,
            DOUT => \N__34162\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34164\,
            PADOUT => \N__34163\,
            PADIN => \N__34162\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34155\,
            DIN => \N__34154\,
            DOUT => \N__34153\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34155\,
            PADOUT => \N__34154\,
            PADIN => \N__34153\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34146\,
            DIN => \N__34145\,
            DOUT => \N__34144\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34146\,
            PADOUT => \N__34145\,
            PADIN => \N__34144\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17582\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34137\,
            DIN => \N__34136\,
            DOUT => \N__34135\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34137\,
            PADOUT => \N__34136\,
            PADIN => \N__34135\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34128\,
            DIN => \N__34127\,
            DOUT => \N__34126\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34128\,
            PADOUT => \N__34127\,
            PADIN => \N__34126\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34119\,
            DIN => \N__34118\,
            DOUT => \N__34117\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34119\,
            PADOUT => \N__34118\,
            PADIN => \N__34117\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34110\,
            DIN => \N__34109\,
            DOUT => \N__34108\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34110\,
            PADOUT => \N__34109\,
            PADIN => \N__34108\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34101\,
            DIN => \N__34100\,
            DOUT => \N__34099\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34101\,
            PADOUT => \N__34100\,
            PADIN => \N__34099\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29269\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34092\,
            DIN => \N__34091\,
            DOUT => \N__34090\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34092\,
            PADOUT => \N__34091\,
            PADIN => \N__34090\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33dsw_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34083\,
            DIN => \N__34082\,
            DOUT => \N__34081\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34083\,
            PADOUT => \N__34082\,
            PADIN => \N__34081\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34074\,
            DIN => \N__34073\,
            DOUT => \N__34072\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34074\,
            PADOUT => \N__34073\,
            PADIN => \N__34072\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31958\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34065\,
            DIN => \N__34064\,
            DOUT => \N__34063\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34065\,
            PADOUT => \N__34064\,
            PADIN => \N__34063\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34056\,
            DIN => \N__34055\,
            DOUT => \N__34054\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34056\,
            PADOUT => \N__34055\,
            PADIN => \N__34054\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34047\,
            DIN => \N__34046\,
            DOUT => \N__34045\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34047\,
            PADOUT => \N__34046\,
            PADIN => \N__34045\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34038\,
            DIN => \N__34037\,
            DOUT => \N__34036\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34038\,
            PADOUT => \N__34037\,
            PADIN => \N__34036\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34029\,
            DIN => \N__34028\,
            DOUT => \N__34027\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34029\,
            PADOUT => \N__34028\,
            PADIN => \N__34027\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22406\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34020\,
            DIN => \N__34019\,
            DOUT => \N__34018\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34020\,
            PADOUT => \N__34019\,
            PADIN => \N__34018\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34011\,
            DIN => \N__34010\,
            DOUT => \N__34009\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34011\,
            PADOUT => \N__34010\,
            PADIN => \N__34009\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30275\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34002\,
            DIN => \N__34001\,
            DOUT => \N__34000\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34002\,
            PADOUT => \N__34001\,
            PADIN => \N__34000\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30335\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33993\,
            DIN => \N__33992\,
            DOUT => \N__33991\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33993\,
            PADOUT => \N__33992\,
            PADIN => \N__33991\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33984\,
            DIN => \N__33983\,
            DOUT => \N__33982\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33984\,
            PADOUT => \N__33983\,
            PADIN => \N__33982\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33975\,
            DIN => \N__33974\,
            DOUT => \N__33973\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33975\,
            PADOUT => \N__33974\,
            PADIN => \N__33973\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33966\,
            DIN => \N__33965\,
            DOUT => \N__33964\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33966\,
            PADOUT => \N__33965\,
            PADIN => \N__33964\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33957\,
            DIN => \N__33956\,
            DOUT => \N__33955\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33957\,
            PADOUT => \N__33956\,
            PADIN => \N__33955\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27460\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33948\,
            DIN => \N__33947\,
            DOUT => \N__33946\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33948\,
            PADOUT => \N__33947\,
            PADIN => \N__33946\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20366\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33939\,
            DIN => \N__33938\,
            DOUT => \N__33937\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33939\,
            PADOUT => \N__33938\,
            PADIN => \N__33937\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33930\,
            DIN => \N__33929\,
            DOUT => \N__33928\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33930\,
            PADOUT => \N__33929\,
            PADIN => \N__33928\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29288\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33921\,
            DIN => \N__33920\,
            DOUT => \N__33919\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33921\,
            PADOUT => \N__33920\,
            PADIN => \N__33919\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33912\,
            DIN => \N__33911\,
            DOUT => \N__33910\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33912\,
            PADOUT => \N__33911\,
            PADIN => \N__33910\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33903\,
            DIN => \N__33902\,
            DOUT => \N__33901\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33903\,
            PADOUT => \N__33902\,
            PADIN => \N__33901\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33894\,
            DIN => \N__33893\,
            DOUT => \N__33892\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33894\,
            PADOUT => \N__33893\,
            PADIN => \N__33892\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33885\,
            DIN => \N__33884\,
            DOUT => \N__33883\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33885\,
            PADOUT => \N__33884\,
            PADIN => \N__33883\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16223\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33876\,
            DIN => \N__33875\,
            DOUT => \N__33874\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33876\,
            PADOUT => \N__33875\,
            PADIN => \N__33874\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33867\,
            DIN => \N__33866\,
            DOUT => \N__33865\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33867\,
            PADOUT => \N__33866\,
            PADIN => \N__33865\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16337\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33858\,
            DIN => \N__33857\,
            DOUT => \N__33856\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33858\,
            PADOUT => \N__33857\,
            PADIN => \N__33856\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33849\,
            DIN => \N__33848\,
            DOUT => \N__33847\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33849\,
            PADOUT => \N__33848\,
            PADIN => \N__33847\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30385\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33840\,
            DIN => \N__33839\,
            DOUT => \N__33838\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33840\,
            PADOUT => \N__33839\,
            PADIN => \N__33838\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16307\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33831\,
            DIN => \N__33830\,
            DOUT => \N__33829\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33831\,
            PADOUT => \N__33830\,
            PADIN => \N__33829\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33822\,
            DIN => \N__33821\,
            DOUT => \N__33820\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33822\,
            PADOUT => \N__33821\,
            PADIN => \N__33820\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__33813\,
            DIN => \N__33812\,
            DOUT => \N__33811\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33813\,
            PADOUT => \N__33812\,
            PADIN => \N__33811\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33804\,
            DIN => \N__33803\,
            DOUT => \N__33802\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33804\,
            PADOUT => \N__33803\,
            PADIN => \N__33802\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33795\,
            DIN => \N__33794\,
            DOUT => \N__33793\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33795\,
            PADOUT => \N__33794\,
            PADIN => \N__33793\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30356\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33786\,
            DIN => \N__33785\,
            DOUT => \N__33784\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33786\,
            PADOUT => \N__33785\,
            PADIN => \N__33784\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33777\,
            DIN => \N__33776\,
            DOUT => \N__33775\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33777\,
            PADOUT => \N__33776\,
            PADIN => \N__33775\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33768\,
            DIN => \N__33767\,
            DOUT => \N__33766\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33768\,
            PADOUT => \N__33767\,
            PADIN => \N__33766\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33759\,
            DIN => \N__33758\,
            DOUT => \N__33757\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33759\,
            PADOUT => \N__33758\,
            PADIN => \N__33757\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33750\,
            DIN => \N__33749\,
            DOUT => \N__33748\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33750\,
            PADOUT => \N__33749\,
            PADIN => \N__33748\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33741\,
            DIN => \N__33740\,
            DOUT => \N__33739\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33741\,
            PADOUT => \N__33740\,
            PADIN => \N__33739\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33732\,
            DIN => \N__33731\,
            DOUT => \N__33730\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33732\,
            PADOUT => \N__33731\,
            PADIN => \N__33730\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30306\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33723\,
            DIN => \N__33722\,
            DOUT => \N__33721\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__33723\,
            PADOUT => \N__33722\,
            PADIN => \N__33721\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__7867\ : CascadeMux
    port map (
            O => \N__33704\,
            I => \N__33700\
        );

    \I__7866\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33695\
        );

    \I__7865\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33695\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__33695\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\
        );

    \I__7863\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33689\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__33689\,
            I => \VPP_VDDQ.count_2_1_10\
        );

    \I__7861\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33682\
        );

    \I__7860\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33679\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__33682\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__33679\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__33674\,
            I => \VPP_VDDQ.count_2_1_10_cascade_\
        );

    \I__7856\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__33668\,
            I => \VPP_VDDQ.un1_count_2_1_axb_10\
        );

    \I__7854\ : CascadeMux
    port map (
            O => \N__33665\,
            I => \N__33651\
        );

    \I__7853\ : CascadeMux
    port map (
            O => \N__33664\,
            I => \N__33648\
        );

    \I__7852\ : CascadeMux
    port map (
            O => \N__33663\,
            I => \N__33644\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__33662\,
            I => \N__33641\
        );

    \I__7850\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33638\
        );

    \I__7849\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33635\
        );

    \I__7848\ : CascadeMux
    port map (
            O => \N__33659\,
            I => \N__33627\
        );

    \I__7847\ : CascadeMux
    port map (
            O => \N__33658\,
            I => \N__33622\
        );

    \I__7846\ : CascadeMux
    port map (
            O => \N__33657\,
            I => \N__33612\
        );

    \I__7845\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33609\
        );

    \I__7844\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33598\
        );

    \I__7843\ : InMux
    port map (
            O => \N__33654\,
            I => \N__33598\
        );

    \I__7842\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33598\
        );

    \I__7841\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33598\
        );

    \I__7840\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33598\
        );

    \I__7839\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33593\
        );

    \I__7838\ : InMux
    port map (
            O => \N__33641\,
            I => \N__33593\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33588\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__33635\,
            I => \N__33588\
        );

    \I__7835\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33577\
        );

    \I__7834\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33577\
        );

    \I__7833\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33577\
        );

    \I__7832\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33577\
        );

    \I__7831\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33577\
        );

    \I__7830\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33568\
        );

    \I__7829\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33568\
        );

    \I__7828\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33568\
        );

    \I__7827\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33568\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__33621\,
            I => \N__33564\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__33620\,
            I => \N__33561\
        );

    \I__7824\ : CascadeMux
    port map (
            O => \N__33619\,
            I => \N__33551\
        );

    \I__7823\ : CascadeMux
    port map (
            O => \N__33618\,
            I => \N__33548\
        );

    \I__7822\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33538\
        );

    \I__7821\ : InMux
    port map (
            O => \N__33616\,
            I => \N__33538\
        );

    \I__7820\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33538\
        );

    \I__7819\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33535\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__33609\,
            I => \N__33522\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__33598\,
            I => \N__33522\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__33593\,
            I => \N__33522\
        );

    \I__7815\ : Span4Mux_v
    port map (
            O => \N__33588\,
            I => \N__33522\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__33577\,
            I => \N__33522\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__33568\,
            I => \N__33522\
        );

    \I__7812\ : InMux
    port map (
            O => \N__33567\,
            I => \N__33507\
        );

    \I__7811\ : InMux
    port map (
            O => \N__33564\,
            I => \N__33507\
        );

    \I__7810\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33507\
        );

    \I__7809\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33507\
        );

    \I__7808\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33507\
        );

    \I__7807\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33507\
        );

    \I__7806\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33507\
        );

    \I__7805\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33502\
        );

    \I__7804\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33502\
        );

    \I__7803\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33495\
        );

    \I__7802\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33495\
        );

    \I__7801\ : InMux
    port map (
            O => \N__33548\,
            I => \N__33495\
        );

    \I__7800\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33488\
        );

    \I__7799\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33488\
        );

    \I__7798\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33488\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__33538\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__33535\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7795\ : Odrv4
    port map (
            O => \N__33522\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__33507\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__33502\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__33495\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__33488\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__33473\,
            I => \N__33467\
        );

    \I__7789\ : CascadeMux
    port map (
            O => \N__33472\,
            I => \N__33461\
        );

    \I__7788\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33447\
        );

    \I__7787\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33436\
        );

    \I__7786\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33436\
        );

    \I__7785\ : InMux
    port map (
            O => \N__33466\,
            I => \N__33436\
        );

    \I__7784\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33436\
        );

    \I__7783\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33436\
        );

    \I__7782\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33419\
        );

    \I__7781\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33419\
        );

    \I__7780\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33419\
        );

    \I__7779\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33419\
        );

    \I__7778\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33406\
        );

    \I__7777\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33406\
        );

    \I__7776\ : InMux
    port map (
            O => \N__33455\,
            I => \N__33406\
        );

    \I__7775\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33406\
        );

    \I__7774\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33406\
        );

    \I__7773\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33406\
        );

    \I__7772\ : CascadeMux
    port map (
            O => \N__33451\,
            I => \N__33403\
        );

    \I__7771\ : CascadeMux
    port map (
            O => \N__33450\,
            I => \N__33394\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33386\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33386\
        );

    \I__7768\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33377\
        );

    \I__7767\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33377\
        );

    \I__7766\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33377\
        );

    \I__7765\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33377\
        );

    \I__7764\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33374\
        );

    \I__7763\ : InMux
    port map (
            O => \N__33430\,
            I => \N__33369\
        );

    \I__7762\ : InMux
    port map (
            O => \N__33429\,
            I => \N__33369\
        );

    \I__7761\ : InMux
    port map (
            O => \N__33428\,
            I => \N__33366\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__33419\,
            I => \N__33361\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__33406\,
            I => \N__33361\
        );

    \I__7758\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33346\
        );

    \I__7757\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33346\
        );

    \I__7756\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33346\
        );

    \I__7755\ : InMux
    port map (
            O => \N__33400\,
            I => \N__33346\
        );

    \I__7754\ : InMux
    port map (
            O => \N__33399\,
            I => \N__33346\
        );

    \I__7753\ : InMux
    port map (
            O => \N__33398\,
            I => \N__33346\
        );

    \I__7752\ : InMux
    port map (
            O => \N__33397\,
            I => \N__33346\
        );

    \I__7751\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33337\
        );

    \I__7750\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33337\
        );

    \I__7749\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33337\
        );

    \I__7748\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33337\
        );

    \I__7747\ : Span4Mux_v
    port map (
            O => \N__33386\,
            I => \N__33332\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__33377\,
            I => \N__33332\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__33374\,
            I => \N__33329\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__33369\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__33366\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7742\ : Odrv12
    port map (
            O => \N__33361\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__33346\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__33337\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__33332\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__33329\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7737\ : CascadeMux
    port map (
            O => \N__33314\,
            I => \N__33310\
        );

    \I__7736\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33307\
        );

    \I__7735\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33304\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__33307\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__33304\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__33299\,
            I => \N__33294\
        );

    \I__7731\ : CascadeMux
    port map (
            O => \N__33298\,
            I => \N__33287\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__33297\,
            I => \N__33274\
        );

    \I__7729\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33257\
        );

    \I__7728\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33257\
        );

    \I__7727\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33257\
        );

    \I__7726\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33257\
        );

    \I__7725\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33257\
        );

    \I__7724\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33254\
        );

    \I__7723\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33245\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33245\
        );

    \I__7721\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33245\
        );

    \I__7720\ : InMux
    port map (
            O => \N__33283\,
            I => \N__33245\
        );

    \I__7719\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33225\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33225\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33225\
        );

    \I__7716\ : InMux
    port map (
            O => \N__33279\,
            I => \N__33225\
        );

    \I__7715\ : InMux
    port map (
            O => \N__33278\,
            I => \N__33225\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33220\
        );

    \I__7713\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33220\
        );

    \I__7712\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33209\
        );

    \I__7711\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33209\
        );

    \I__7710\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33209\
        );

    \I__7709\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33209\
        );

    \I__7708\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33209\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33204\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__33257\,
            I => \N__33197\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33197\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33245\,
            I => \N__33197\
        );

    \I__7703\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33184\
        );

    \I__7702\ : InMux
    port map (
            O => \N__33243\,
            I => \N__33184\
        );

    \I__7701\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33184\
        );

    \I__7700\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33184\
        );

    \I__7699\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33184\
        );

    \I__7698\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33184\
        );

    \I__7697\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33177\
        );

    \I__7696\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33177\
        );

    \I__7695\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33177\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__33225\,
            I => \N__33170\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__33220\,
            I => \N__33170\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__33209\,
            I => \N__33170\
        );

    \I__7691\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33165\
        );

    \I__7690\ : InMux
    port map (
            O => \N__33207\,
            I => \N__33165\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__33204\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7688\ : Odrv4
    port map (
            O => \N__33197\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__33184\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__33177\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7685\ : Odrv4
    port map (
            O => \N__33170\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__33165\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7683\ : InMux
    port map (
            O => \N__33152\,
            I => \N__33149\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__33149\,
            I => \VPP_VDDQ.count_2_0_12\
        );

    \I__7681\ : ClkMux
    port map (
            O => \N__33146\,
            I => \N__33143\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N__33132\
        );

    \I__7679\ : ClkMux
    port map (
            O => \N__33142\,
            I => \N__33129\
        );

    \I__7678\ : ClkMux
    port map (
            O => \N__33141\,
            I => \N__33124\
        );

    \I__7677\ : ClkMux
    port map (
            O => \N__33140\,
            I => \N__33120\
        );

    \I__7676\ : ClkMux
    port map (
            O => \N__33139\,
            I => \N__33117\
        );

    \I__7675\ : ClkMux
    port map (
            O => \N__33138\,
            I => \N__33114\
        );

    \I__7674\ : ClkMux
    port map (
            O => \N__33137\,
            I => \N__33107\
        );

    \I__7673\ : ClkMux
    port map (
            O => \N__33136\,
            I => \N__33104\
        );

    \I__7672\ : ClkMux
    port map (
            O => \N__33135\,
            I => \N__33101\
        );

    \I__7671\ : Span4Mux_s2_h
    port map (
            O => \N__33132\,
            I => \N__33094\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__33129\,
            I => \N__33094\
        );

    \I__7669\ : ClkMux
    port map (
            O => \N__33128\,
            I => \N__33091\
        );

    \I__7668\ : ClkMux
    port map (
            O => \N__33127\,
            I => \N__33087\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__33124\,
            I => \N__33082\
        );

    \I__7666\ : ClkMux
    port map (
            O => \N__33123\,
            I => \N__33079\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__33120\,
            I => \N__33072\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33072\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__33114\,
            I => \N__33063\
        );

    \I__7662\ : ClkMux
    port map (
            O => \N__33113\,
            I => \N__33060\
        );

    \I__7661\ : ClkMux
    port map (
            O => \N__33112\,
            I => \N__33056\
        );

    \I__7660\ : ClkMux
    port map (
            O => \N__33111\,
            I => \N__33053\
        );

    \I__7659\ : ClkMux
    port map (
            O => \N__33110\,
            I => \N__33045\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__33107\,
            I => \N__33042\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__33104\,
            I => \N__33039\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__33101\,
            I => \N__33036\
        );

    \I__7655\ : ClkMux
    port map (
            O => \N__33100\,
            I => \N__33033\
        );

    \I__7654\ : ClkMux
    port map (
            O => \N__33099\,
            I => \N__33030\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__33094\,
            I => \N__33023\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__33091\,
            I => \N__33023\
        );

    \I__7651\ : ClkMux
    port map (
            O => \N__33090\,
            I => \N__33020\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__33087\,
            I => \N__33017\
        );

    \I__7649\ : ClkMux
    port map (
            O => \N__33086\,
            I => \N__33013\
        );

    \I__7648\ : ClkMux
    port map (
            O => \N__33085\,
            I => \N__33010\
        );

    \I__7647\ : Span4Mux_s2_h
    port map (
            O => \N__33082\,
            I => \N__33005\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__33079\,
            I => \N__33005\
        );

    \I__7645\ : ClkMux
    port map (
            O => \N__33078\,
            I => \N__33002\
        );

    \I__7644\ : ClkMux
    port map (
            O => \N__33077\,
            I => \N__32999\
        );

    \I__7643\ : Span4Mux_h
    port map (
            O => \N__33072\,
            I => \N__32996\
        );

    \I__7642\ : ClkMux
    port map (
            O => \N__33071\,
            I => \N__32993\
        );

    \I__7641\ : ClkMux
    port map (
            O => \N__33070\,
            I => \N__32990\
        );

    \I__7640\ : ClkMux
    port map (
            O => \N__33069\,
            I => \N__32986\
        );

    \I__7639\ : ClkMux
    port map (
            O => \N__33068\,
            I => \N__32982\
        );

    \I__7638\ : ClkMux
    port map (
            O => \N__33067\,
            I => \N__32978\
        );

    \I__7637\ : ClkMux
    port map (
            O => \N__33066\,
            I => \N__32975\
        );

    \I__7636\ : Span4Mux_v
    port map (
            O => \N__33063\,
            I => \N__32968\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__33060\,
            I => \N__32965\
        );

    \I__7634\ : ClkMux
    port map (
            O => \N__33059\,
            I => \N__32960\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__33056\,
            I => \N__32956\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__33053\,
            I => \N__32953\
        );

    \I__7631\ : ClkMux
    port map (
            O => \N__33052\,
            I => \N__32950\
        );

    \I__7630\ : ClkMux
    port map (
            O => \N__33051\,
            I => \N__32945\
        );

    \I__7629\ : ClkMux
    port map (
            O => \N__33050\,
            I => \N__32939\
        );

    \I__7628\ : ClkMux
    port map (
            O => \N__33049\,
            I => \N__32936\
        );

    \I__7627\ : ClkMux
    port map (
            O => \N__33048\,
            I => \N__32932\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__32929\
        );

    \I__7625\ : Span4Mux_v
    port map (
            O => \N__33042\,
            I => \N__32918\
        );

    \I__7624\ : Span4Mux_v
    port map (
            O => \N__33039\,
            I => \N__32918\
        );

    \I__7623\ : Span4Mux_s1_h
    port map (
            O => \N__33036\,
            I => \N__32918\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__33033\,
            I => \N__32918\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__33030\,
            I => \N__32915\
        );

    \I__7620\ : ClkMux
    port map (
            O => \N__33029\,
            I => \N__32912\
        );

    \I__7619\ : ClkMux
    port map (
            O => \N__33028\,
            I => \N__32908\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__33023\,
            I => \N__32901\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__33020\,
            I => \N__32901\
        );

    \I__7616\ : Span4Mux_s2_h
    port map (
            O => \N__33017\,
            I => \N__32896\
        );

    \I__7615\ : ClkMux
    port map (
            O => \N__33016\,
            I => \N__32893\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__33013\,
            I => \N__32888\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__33010\,
            I => \N__32888\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__33005\,
            I => \N__32884\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__33002\,
            I => \N__32879\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__32999\,
            I => \N__32879\
        );

    \I__7609\ : Span4Mux_v
    port map (
            O => \N__32996\,
            I => \N__32872\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__32993\,
            I => \N__32872\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__32990\,
            I => \N__32872\
        );

    \I__7606\ : ClkMux
    port map (
            O => \N__32989\,
            I => \N__32869\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__32986\,
            I => \N__32866\
        );

    \I__7604\ : ClkMux
    port map (
            O => \N__32985\,
            I => \N__32863\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32860\
        );

    \I__7602\ : ClkMux
    port map (
            O => \N__32981\,
            I => \N__32857\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32854\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32851\
        );

    \I__7599\ : ClkMux
    port map (
            O => \N__32974\,
            I => \N__32848\
        );

    \I__7598\ : ClkMux
    port map (
            O => \N__32973\,
            I => \N__32845\
        );

    \I__7597\ : ClkMux
    port map (
            O => \N__32972\,
            I => \N__32840\
        );

    \I__7596\ : ClkMux
    port map (
            O => \N__32971\,
            I => \N__32837\
        );

    \I__7595\ : Span4Mux_h
    port map (
            O => \N__32968\,
            I => \N__32832\
        );

    \I__7594\ : Span4Mux_v
    port map (
            O => \N__32965\,
            I => \N__32832\
        );

    \I__7593\ : ClkMux
    port map (
            O => \N__32964\,
            I => \N__32829\
        );

    \I__7592\ : ClkMux
    port map (
            O => \N__32963\,
            I => \N__32826\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32823\
        );

    \I__7590\ : ClkMux
    port map (
            O => \N__32959\,
            I => \N__32820\
        );

    \I__7589\ : Span4Mux_v
    port map (
            O => \N__32956\,
            I => \N__32814\
        );

    \I__7588\ : Span4Mux_s1_h
    port map (
            O => \N__32953\,
            I => \N__32814\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__32950\,
            I => \N__32811\
        );

    \I__7586\ : ClkMux
    port map (
            O => \N__32949\,
            I => \N__32808\
        );

    \I__7585\ : ClkMux
    port map (
            O => \N__32948\,
            I => \N__32805\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32802\
        );

    \I__7583\ : ClkMux
    port map (
            O => \N__32944\,
            I => \N__32799\
        );

    \I__7582\ : ClkMux
    port map (
            O => \N__32943\,
            I => \N__32795\
        );

    \I__7581\ : ClkMux
    port map (
            O => \N__32942\,
            I => \N__32791\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__32939\,
            I => \N__32788\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__32936\,
            I => \N__32785\
        );

    \I__7578\ : ClkMux
    port map (
            O => \N__32935\,
            I => \N__32782\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32777\
        );

    \I__7576\ : Span4Mux_h
    port map (
            O => \N__32929\,
            I => \N__32777\
        );

    \I__7575\ : ClkMux
    port map (
            O => \N__32928\,
            I => \N__32773\
        );

    \I__7574\ : ClkMux
    port map (
            O => \N__32927\,
            I => \N__32770\
        );

    \I__7573\ : Span4Mux_v
    port map (
            O => \N__32918\,
            I => \N__32764\
        );

    \I__7572\ : Span4Mux_h
    port map (
            O => \N__32915\,
            I => \N__32764\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__32912\,
            I => \N__32761\
        );

    \I__7570\ : ClkMux
    port map (
            O => \N__32911\,
            I => \N__32758\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__32908\,
            I => \N__32755\
        );

    \I__7568\ : ClkMux
    port map (
            O => \N__32907\,
            I => \N__32752\
        );

    \I__7567\ : ClkMux
    port map (
            O => \N__32906\,
            I => \N__32749\
        );

    \I__7566\ : Span4Mux_v
    port map (
            O => \N__32901\,
            I => \N__32744\
        );

    \I__7565\ : ClkMux
    port map (
            O => \N__32900\,
            I => \N__32741\
        );

    \I__7564\ : ClkMux
    port map (
            O => \N__32899\,
            I => \N__32738\
        );

    \I__7563\ : Span4Mux_h
    port map (
            O => \N__32896\,
            I => \N__32731\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__32893\,
            I => \N__32731\
        );

    \I__7561\ : Span4Mux_h
    port map (
            O => \N__32888\,
            I => \N__32731\
        );

    \I__7560\ : ClkMux
    port map (
            O => \N__32887\,
            I => \N__32728\
        );

    \I__7559\ : Span4Mux_v
    port map (
            O => \N__32884\,
            I => \N__32719\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__32879\,
            I => \N__32719\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__32872\,
            I => \N__32719\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__32869\,
            I => \N__32719\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__32866\,
            I => \N__32714\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__32863\,
            I => \N__32714\
        );

    \I__7553\ : Span4Mux_s2_h
    port map (
            O => \N__32860\,
            I => \N__32709\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32709\
        );

    \I__7551\ : Span4Mux_v
    port map (
            O => \N__32854\,
            I => \N__32700\
        );

    \I__7550\ : Span4Mux_v
    port map (
            O => \N__32851\,
            I => \N__32700\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__32848\,
            I => \N__32700\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__32845\,
            I => \N__32700\
        );

    \I__7547\ : ClkMux
    port map (
            O => \N__32844\,
            I => \N__32697\
        );

    \I__7546\ : ClkMux
    port map (
            O => \N__32843\,
            I => \N__32694\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32690\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32687\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__32832\,
            I => \N__32680\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__32829\,
            I => \N__32680\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__32826\,
            I => \N__32677\
        );

    \I__7540\ : Span4Mux_v
    port map (
            O => \N__32823\,
            I => \N__32672\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__32820\,
            I => \N__32672\
        );

    \I__7538\ : ClkMux
    port map (
            O => \N__32819\,
            I => \N__32669\
        );

    \I__7537\ : Span4Mux_h
    port map (
            O => \N__32814\,
            I => \N__32660\
        );

    \I__7536\ : Span4Mux_v
    port map (
            O => \N__32811\,
            I => \N__32660\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__32808\,
            I => \N__32660\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__32805\,
            I => \N__32660\
        );

    \I__7533\ : Span4Mux_s1_h
    port map (
            O => \N__32802\,
            I => \N__32655\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__32799\,
            I => \N__32655\
        );

    \I__7531\ : ClkMux
    port map (
            O => \N__32798\,
            I => \N__32652\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__32795\,
            I => \N__32649\
        );

    \I__7529\ : ClkMux
    port map (
            O => \N__32794\,
            I => \N__32646\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__32791\,
            I => \N__32643\
        );

    \I__7527\ : Span4Mux_v
    port map (
            O => \N__32788\,
            I => \N__32640\
        );

    \I__7526\ : Span4Mux_s1_h
    port map (
            O => \N__32785\,
            I => \N__32635\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__32782\,
            I => \N__32635\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__32777\,
            I => \N__32631\
        );

    \I__7523\ : ClkMux
    port map (
            O => \N__32776\,
            I => \N__32628\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__32773\,
            I => \N__32625\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__32770\,
            I => \N__32622\
        );

    \I__7520\ : ClkMux
    port map (
            O => \N__32769\,
            I => \N__32619\
        );

    \I__7519\ : Span4Mux_v
    port map (
            O => \N__32764\,
            I => \N__32612\
        );

    \I__7518\ : Span4Mux_v
    port map (
            O => \N__32761\,
            I => \N__32612\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__32758\,
            I => \N__32612\
        );

    \I__7516\ : Span4Mux_s1_h
    port map (
            O => \N__32755\,
            I => \N__32605\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__32752\,
            I => \N__32605\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__32749\,
            I => \N__32605\
        );

    \I__7513\ : ClkMux
    port map (
            O => \N__32748\,
            I => \N__32602\
        );

    \I__7512\ : ClkMux
    port map (
            O => \N__32747\,
            I => \N__32599\
        );

    \I__7511\ : Span4Mux_v
    port map (
            O => \N__32744\,
            I => \N__32592\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__32741\,
            I => \N__32592\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__32738\,
            I => \N__32592\
        );

    \I__7508\ : Span4Mux_v
    port map (
            O => \N__32731\,
            I => \N__32587\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__32728\,
            I => \N__32587\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__32719\,
            I => \N__32580\
        );

    \I__7505\ : Span4Mux_h
    port map (
            O => \N__32714\,
            I => \N__32580\
        );

    \I__7504\ : Span4Mux_h
    port map (
            O => \N__32709\,
            I => \N__32580\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__32700\,
            I => \N__32573\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__32697\,
            I => \N__32573\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__32694\,
            I => \N__32573\
        );

    \I__7500\ : ClkMux
    port map (
            O => \N__32693\,
            I => \N__32570\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__32690\,
            I => \N__32564\
        );

    \I__7498\ : Span4Mux_h
    port map (
            O => \N__32687\,
            I => \N__32564\
        );

    \I__7497\ : ClkMux
    port map (
            O => \N__32686\,
            I => \N__32561\
        );

    \I__7496\ : ClkMux
    port map (
            O => \N__32685\,
            I => \N__32558\
        );

    \I__7495\ : Span4Mux_v
    port map (
            O => \N__32680\,
            I => \N__32555\
        );

    \I__7494\ : Span4Mux_v
    port map (
            O => \N__32677\,
            I => \N__32548\
        );

    \I__7493\ : Span4Mux_s2_h
    port map (
            O => \N__32672\,
            I => \N__32548\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__32669\,
            I => \N__32548\
        );

    \I__7491\ : Span4Mux_v
    port map (
            O => \N__32660\,
            I => \N__32541\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__32655\,
            I => \N__32541\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__32652\,
            I => \N__32541\
        );

    \I__7488\ : Span4Mux_h
    port map (
            O => \N__32649\,
            I => \N__32534\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__32646\,
            I => \N__32534\
        );

    \I__7486\ : Span4Mux_h
    port map (
            O => \N__32643\,
            I => \N__32534\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__32640\,
            I => \N__32529\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__32635\,
            I => \N__32529\
        );

    \I__7483\ : ClkMux
    port map (
            O => \N__32634\,
            I => \N__32526\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__32631\,
            I => \N__32521\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__32628\,
            I => \N__32521\
        );

    \I__7480\ : Span4Mux_s2_h
    port map (
            O => \N__32625\,
            I => \N__32512\
        );

    \I__7479\ : Span4Mux_s2_h
    port map (
            O => \N__32622\,
            I => \N__32512\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__32619\,
            I => \N__32512\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__32612\,
            I => \N__32512\
        );

    \I__7476\ : Span4Mux_v
    port map (
            O => \N__32605\,
            I => \N__32507\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__32602\,
            I => \N__32507\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32504\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__32592\,
            I => \N__32493\
        );

    \I__7472\ : Span4Mux_v
    port map (
            O => \N__32587\,
            I => \N__32493\
        );

    \I__7471\ : IoSpan4Mux
    port map (
            O => \N__32580\,
            I => \N__32493\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__32573\,
            I => \N__32493\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32493\
        );

    \I__7468\ : ClkMux
    port map (
            O => \N__32569\,
            I => \N__32490\
        );

    \I__7467\ : Span4Mux_v
    port map (
            O => \N__32564\,
            I => \N__32482\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__32561\,
            I => \N__32482\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__32558\,
            I => \N__32482\
        );

    \I__7464\ : IoSpan4Mux
    port map (
            O => \N__32555\,
            I => \N__32479\
        );

    \I__7463\ : Span4Mux_h
    port map (
            O => \N__32548\,
            I => \N__32472\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__32541\,
            I => \N__32472\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__32534\,
            I => \N__32472\
        );

    \I__7460\ : Span4Mux_v
    port map (
            O => \N__32529\,
            I => \N__32467\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__32526\,
            I => \N__32467\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__32521\,
            I => \N__32460\
        );

    \I__7457\ : Span4Mux_h
    port map (
            O => \N__32512\,
            I => \N__32460\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__32507\,
            I => \N__32460\
        );

    \I__7455\ : IoSpan4Mux
    port map (
            O => \N__32504\,
            I => \N__32455\
        );

    \I__7454\ : IoSpan4Mux
    port map (
            O => \N__32493\,
            I => \N__32455\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__32490\,
            I => \N__32452\
        );

    \I__7452\ : ClkMux
    port map (
            O => \N__32489\,
            I => \N__32449\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__32482\,
            I => \N__32446\
        );

    \I__7450\ : Odrv4
    port map (
            O => \N__32479\,
            I => fpga_osc
        );

    \I__7449\ : Odrv4
    port map (
            O => \N__32472\,
            I => fpga_osc
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__32467\,
            I => fpga_osc
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__32460\,
            I => fpga_osc
        );

    \I__7446\ : Odrv4
    port map (
            O => \N__32455\,
            I => fpga_osc
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__32452\,
            I => fpga_osc
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__32449\,
            I => fpga_osc
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__32446\,
            I => fpga_osc
        );

    \I__7442\ : CEMux
    port map (
            O => \N__32429\,
            I => \N__32426\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__32426\,
            I => \N__32422\
        );

    \I__7440\ : CEMux
    port map (
            O => \N__32425\,
            I => \N__32419\
        );

    \I__7439\ : Span4Mux_v
    port map (
            O => \N__32422\,
            I => \N__32413\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__32419\,
            I => \N__32413\
        );

    \I__7437\ : CEMux
    port map (
            O => \N__32418\,
            I => \N__32410\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__32413\,
            I => \N__32404\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__32410\,
            I => \N__32404\
        );

    \I__7434\ : CEMux
    port map (
            O => \N__32409\,
            I => \N__32397\
        );

    \I__7433\ : Span4Mux_h
    port map (
            O => \N__32404\,
            I => \N__32394\
        );

    \I__7432\ : CEMux
    port map (
            O => \N__32403\,
            I => \N__32391\
        );

    \I__7431\ : InMux
    port map (
            O => \N__32402\,
            I => \N__32388\
        );

    \I__7430\ : InMux
    port map (
            O => \N__32401\,
            I => \N__32383\
        );

    \I__7429\ : InMux
    port map (
            O => \N__32400\,
            I => \N__32383\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__32397\,
            I => \N__32369\
        );

    \I__7427\ : Span4Mux_s0_h
    port map (
            O => \N__32394\,
            I => \N__32369\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__32391\,
            I => \N__32369\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__32388\,
            I => \N__32364\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__32383\,
            I => \N__32364\
        );

    \I__7423\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32351\
        );

    \I__7422\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32351\
        );

    \I__7421\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32346\
        );

    \I__7420\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32346\
        );

    \I__7419\ : InMux
    port map (
            O => \N__32378\,
            I => \N__32339\
        );

    \I__7418\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32339\
        );

    \I__7417\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32339\
        );

    \I__7416\ : Span4Mux_v
    port map (
            O => \N__32369\,
            I => \N__32334\
        );

    \I__7415\ : Span4Mux_h
    port map (
            O => \N__32364\,
            I => \N__32334\
        );

    \I__7414\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32328\
        );

    \I__7413\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32325\
        );

    \I__7412\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32312\
        );

    \I__7411\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32312\
        );

    \I__7410\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32312\
        );

    \I__7409\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32312\
        );

    \I__7408\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32312\
        );

    \I__7407\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32312\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32303\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__32346\,
            I => \N__32303\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__32339\,
            I => \N__32303\
        );

    \I__7403\ : Span4Mux_v
    port map (
            O => \N__32334\,
            I => \N__32303\
        );

    \I__7402\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32296\
        );

    \I__7401\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32296\
        );

    \I__7400\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32296\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__32328\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__32325\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__32312\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__7396\ : Odrv4
    port map (
            O => \N__32303\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__32296\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__32285\,
            I => \N__32282\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32282\,
            I => \N__32278\
        );

    \I__7392\ : InMux
    port map (
            O => \N__32281\,
            I => \N__32275\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__32278\,
            I => \N__32272\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__32275\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__32272\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__7388\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32264\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__7386\ : Odrv12
    port map (
            O => \N__32261\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__7385\ : CascadeMux
    port map (
            O => \N__32258\,
            I => \N__32255\
        );

    \I__7384\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32251\
        );

    \I__7383\ : InMux
    port map (
            O => \N__32254\,
            I => \N__32248\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__32251\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__32248\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32240\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__32240\,
            I => \N__32237\
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__32237\,
            I => \VPP_VDDQ.count_2_0_6\
        );

    \I__7377\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32231\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__32231\,
            I => \N__32228\
        );

    \I__7375\ : Span4Mux_h
    port map (
            O => \N__32228\,
            I => \N__32225\
        );

    \I__7374\ : Span4Mux_v
    port map (
            O => \N__32225\,
            I => \N__32222\
        );

    \I__7373\ : Odrv4
    port map (
            O => \N__32222\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__7372\ : CascadeMux
    port map (
            O => \N__32219\,
            I => \N__32215\
        );

    \I__7371\ : InMux
    port map (
            O => \N__32218\,
            I => \N__32210\
        );

    \I__7370\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32210\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__32210\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\
        );

    \I__7368\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32204\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__32204\,
            I => \N__32201\
        );

    \I__7366\ : Span12Mux_s11_v
    port map (
            O => \N__32201\,
            I => \N__32198\
        );

    \I__7365\ : Odrv12
    port map (
            O => \N__32198\,
            I => \VPP_VDDQ.count_2_1_8\
        );

    \I__7364\ : CascadeMux
    port map (
            O => \N__32195\,
            I => \VPP_VDDQ.count_2_1_11_cascade_\
        );

    \I__7363\ : InMux
    port map (
            O => \N__32192\,
            I => \N__32189\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__32189\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__32186\,
            I => \VPP_VDDQ.count_2Z0Z_11_cascade_\
        );

    \I__7360\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32180\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__32180\,
            I => \N__32177\
        );

    \I__7358\ : Odrv12
    port map (
            O => \N__32177\,
            I => \VPP_VDDQ.un9_clk_100khz_5\
        );

    \I__7357\ : CascadeMux
    port map (
            O => \N__32174\,
            I => \N__32170\
        );

    \I__7356\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32165\
        );

    \I__7355\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32165\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__32165\,
            I => \N__32162\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__32162\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\
        );

    \I__7352\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32156\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__32156\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__7350\ : CascadeMux
    port map (
            O => \N__32153\,
            I => \VPP_VDDQ.N_1_i_cascade_\
        );

    \I__7349\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32146\
        );

    \I__7348\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32143\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__32146\,
            I => \N__32138\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__32143\,
            I => \N__32138\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__32138\,
            I => \N__32132\
        );

    \I__7344\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32127\
        );

    \I__7343\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32127\
        );

    \I__7342\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32124\
        );

    \I__7341\ : Span4Mux_v
    port map (
            O => \N__32132\,
            I => \N__32121\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__32127\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__32124\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7338\ : Odrv4
    port map (
            O => \N__32121\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7337\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32111\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__32111\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__7335\ : CascadeMux
    port map (
            O => \N__32108\,
            I => \N__32105\
        );

    \I__7334\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32099\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32104\,
            I => \N__32099\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__32099\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\
        );

    \I__7331\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32093\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__32093\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__7329\ : CascadeMux
    port map (
            O => \N__32090\,
            I => \N__32087\
        );

    \I__7328\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32081\
        );

    \I__7327\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32081\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__32081\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__32078\,
            I => \VPP_VDDQ.count_2_1_7_cascade_\
        );

    \I__7324\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32072\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__32072\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__32069\,
            I => \VPP_VDDQ.count_2_1_12_cascade_\
        );

    \I__7321\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32060\
        );

    \I__7320\ : InMux
    port map (
            O => \N__32065\,
            I => \N__32060\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__32060\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__32057\,
            I => \N__32053\
        );

    \I__7317\ : CascadeMux
    port map (
            O => \N__32056\,
            I => \N__32050\
        );

    \I__7316\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32047\
        );

    \I__7315\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32044\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__32047\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__32044\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__7312\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32036\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__32036\,
            I => \VPP_VDDQ.count_2_0_14\
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__32033\,
            I => \VPP_VDDQ.count_2_1_14_cascade_\
        );

    \I__7309\ : InMux
    port map (
            O => \N__32030\,
            I => \N__32026\
        );

    \I__7308\ : InMux
    port map (
            O => \N__32029\,
            I => \N__32023\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__32026\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__32023\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__7305\ : InMux
    port map (
            O => \N__32018\,
            I => \N__32015\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__32015\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__7303\ : CascadeMux
    port map (
            O => \N__32012\,
            I => \VPP_VDDQ.m4_0_cascade_\
        );

    \I__7302\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32005\
        );

    \I__7301\ : InMux
    port map (
            O => \N__32008\,
            I => \N__31982\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__32005\,
            I => \N__31979\
        );

    \I__7299\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31976\
        );

    \I__7298\ : InMux
    port map (
            O => \N__32003\,
            I => \N__31973\
        );

    \I__7297\ : InMux
    port map (
            O => \N__32002\,
            I => \N__31970\
        );

    \I__7296\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31964\
        );

    \I__7295\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31961\
        );

    \I__7294\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31955\
        );

    \I__7293\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31952\
        );

    \I__7292\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31943\
        );

    \I__7291\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31943\
        );

    \I__7290\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31943\
        );

    \I__7289\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31943\
        );

    \I__7288\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31938\
        );

    \I__7287\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31938\
        );

    \I__7286\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31931\
        );

    \I__7285\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31931\
        );

    \I__7284\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31931\
        );

    \I__7283\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31928\
        );

    \I__7282\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31921\
        );

    \I__7281\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31921\
        );

    \I__7280\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31921\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31916\
        );

    \I__7278\ : Span4Mux_s1_h
    port map (
            O => \N__31979\,
            I => \N__31916\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31913\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__31973\,
            I => \N__31908\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__31970\,
            I => \N__31908\
        );

    \I__7274\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31901\
        );

    \I__7273\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31901\
        );

    \I__7272\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31901\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__31964\,
            I => \N__31896\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31896\
        );

    \I__7269\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31891\
        );

    \I__7268\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31891\
        );

    \I__7267\ : IoInMux
    port map (
            O => \N__31958\,
            I => \N__31886\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__31955\,
            I => \N__31882\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31879\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__31943\,
            I => \N__31872\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__31938\,
            I => \N__31872\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31872\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__31928\,
            I => \N__31865\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__31921\,
            I => \N__31865\
        );

    \I__7259\ : Span4Mux_h
    port map (
            O => \N__31916\,
            I => \N__31865\
        );

    \I__7258\ : Span4Mux_s1_v
    port map (
            O => \N__31913\,
            I => \N__31862\
        );

    \I__7257\ : Span4Mux_v
    port map (
            O => \N__31908\,
            I => \N__31857\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__31901\,
            I => \N__31857\
        );

    \I__7255\ : Span4Mux_v
    port map (
            O => \N__31896\,
            I => \N__31854\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__31891\,
            I => \N__31851\
        );

    \I__7253\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31846\
        );

    \I__7252\ : InMux
    port map (
            O => \N__31889\,
            I => \N__31846\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__31886\,
            I => \N__31843\
        );

    \I__7250\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31840\
        );

    \I__7249\ : Span4Mux_v
    port map (
            O => \N__31882\,
            I => \N__31835\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__31879\,
            I => \N__31835\
        );

    \I__7247\ : Span12Mux_v
    port map (
            O => \N__31872\,
            I => \N__31832\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__31865\,
            I => \N__31827\
        );

    \I__7245\ : Span4Mux_h
    port map (
            O => \N__31862\,
            I => \N__31827\
        );

    \I__7244\ : Span4Mux_h
    port map (
            O => \N__31857\,
            I => \N__31818\
        );

    \I__7243\ : Span4Mux_h
    port map (
            O => \N__31854\,
            I => \N__31818\
        );

    \I__7242\ : Span4Mux_h
    port map (
            O => \N__31851\,
            I => \N__31818\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__31846\,
            I => \N__31818\
        );

    \I__7240\ : Odrv12
    port map (
            O => \N__31843\,
            I => suswarn_n
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__31840\,
            I => suswarn_n
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__31835\,
            I => suswarn_n
        );

    \I__7237\ : Odrv12
    port map (
            O => \N__31832\,
            I => suswarn_n
        );

    \I__7236\ : Odrv4
    port map (
            O => \N__31827\,
            I => suswarn_n
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__31818\,
            I => suswarn_n
        );

    \I__7234\ : CascadeMux
    port map (
            O => \N__31805\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__31802\,
            I => \N__31796\
        );

    \I__7232\ : InMux
    port map (
            O => \N__31801\,
            I => \N__31790\
        );

    \I__7231\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31787\
        );

    \I__7230\ : InMux
    port map (
            O => \N__31799\,
            I => \N__31784\
        );

    \I__7229\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31779\
        );

    \I__7228\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31779\
        );

    \I__7227\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31776\
        );

    \I__7226\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31773\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__31790\,
            I => \N__31760\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__31787\,
            I => \N__31757\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__31784\,
            I => \N__31754\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31751\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__31776\,
            I => \N__31748\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__31773\,
            I => \N__31745\
        );

    \I__7219\ : CEMux
    port map (
            O => \N__31772\,
            I => \N__31712\
        );

    \I__7218\ : CEMux
    port map (
            O => \N__31771\,
            I => \N__31712\
        );

    \I__7217\ : CEMux
    port map (
            O => \N__31770\,
            I => \N__31712\
        );

    \I__7216\ : CEMux
    port map (
            O => \N__31769\,
            I => \N__31712\
        );

    \I__7215\ : CEMux
    port map (
            O => \N__31768\,
            I => \N__31712\
        );

    \I__7214\ : CEMux
    port map (
            O => \N__31767\,
            I => \N__31712\
        );

    \I__7213\ : CEMux
    port map (
            O => \N__31766\,
            I => \N__31712\
        );

    \I__7212\ : CEMux
    port map (
            O => \N__31765\,
            I => \N__31712\
        );

    \I__7211\ : CEMux
    port map (
            O => \N__31764\,
            I => \N__31712\
        );

    \I__7210\ : CEMux
    port map (
            O => \N__31763\,
            I => \N__31712\
        );

    \I__7209\ : Glb2LocalMux
    port map (
            O => \N__31760\,
            I => \N__31712\
        );

    \I__7208\ : Glb2LocalMux
    port map (
            O => \N__31757\,
            I => \N__31712\
        );

    \I__7207\ : Glb2LocalMux
    port map (
            O => \N__31754\,
            I => \N__31712\
        );

    \I__7206\ : Glb2LocalMux
    port map (
            O => \N__31751\,
            I => \N__31712\
        );

    \I__7205\ : Glb2LocalMux
    port map (
            O => \N__31748\,
            I => \N__31712\
        );

    \I__7204\ : Glb2LocalMux
    port map (
            O => \N__31745\,
            I => \N__31712\
        );

    \I__7203\ : GlobalMux
    port map (
            O => \N__31712\,
            I => \N__31709\
        );

    \I__7202\ : gio2CtrlBuf
    port map (
            O => \N__31709\,
            I => \N_579_g\
        );

    \I__7201\ : CascadeMux
    port map (
            O => \N__31706\,
            I => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_\
        );

    \I__7200\ : CascadeMux
    port map (
            O => \N__31703\,
            I => \N__31700\
        );

    \I__7199\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31697\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__31697\,
            I => \N__31693\
        );

    \I__7197\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31690\
        );

    \I__7196\ : Odrv4
    port map (
            O => \N__31693\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__31690\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__7194\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31682\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__31682\,
            I => \VPP_VDDQ.count_2_1_6\
        );

    \I__7192\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31667\
        );

    \I__7191\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31667\
        );

    \I__7190\ : InMux
    port map (
            O => \N__31677\,
            I => \N__31667\
        );

    \I__7189\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31667\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__31667\,
            I => \N__31664\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__31664\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__31661\,
            I => \N__31655\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__31660\,
            I => \N__31650\
        );

    \I__7184\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31643\
        );

    \I__7183\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31643\
        );

    \I__7182\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31643\
        );

    \I__7181\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31636\
        );

    \I__7180\ : InMux
    port map (
            O => \N__31653\,
            I => \N__31636\
        );

    \I__7179\ : InMux
    port map (
            O => \N__31650\,
            I => \N__31636\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__31643\,
            I => \N__31633\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__31636\,
            I => \N__31630\
        );

    \I__7176\ : Span4Mux_v
    port map (
            O => \N__31633\,
            I => \N__31626\
        );

    \I__7175\ : Span4Mux_s1_h
    port map (
            O => \N__31630\,
            I => \N__31623\
        );

    \I__7174\ : InMux
    port map (
            O => \N__31629\,
            I => \N__31620\
        );

    \I__7173\ : Span4Mux_v
    port map (
            O => \N__31626\,
            I => \N__31617\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__31623\,
            I => \N__31612\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__31620\,
            I => \N__31612\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__31617\,
            I => vddq_ok
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__31612\,
            I => vddq_ok
        );

    \I__7168\ : InMux
    port map (
            O => \N__31607\,
            I => \N__31604\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__31604\,
            I => \N__31600\
        );

    \I__7166\ : CascadeMux
    port map (
            O => \N__31603\,
            I => \N__31596\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__31600\,
            I => \N__31592\
        );

    \I__7164\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31587\
        );

    \I__7163\ : InMux
    port map (
            O => \N__31596\,
            I => \N__31587\
        );

    \I__7162\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31584\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__31592\,
            I => \N_362\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__31587\,
            I => \N_362\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__31584\,
            I => \N_362\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__31577\,
            I => \VPP_VDDQ.count_2_1_0_cascade_\
        );

    \I__7157\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31570\
        );

    \I__7156\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31567\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__31570\,
            I => \N__31562\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__31567\,
            I => \N__31562\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__31562\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__7152\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31556\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__31556\,
            I => \VPP_VDDQ.un9_clk_100khz_12\
        );

    \I__7150\ : CascadeMux
    port map (
            O => \N__31553\,
            I => \VPP_VDDQ.un9_clk_100khz_4_cascade_\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31547\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__31547\,
            I => \VPP_VDDQ.un9_clk_100khz_11\
        );

    \I__7147\ : CascadeMux
    port map (
            O => \N__31544\,
            I => \VPP_VDDQ.N_47_cascade_\
        );

    \I__7146\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31537\
        );

    \I__7145\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31534\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__31537\,
            I => \N__31529\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__31534\,
            I => \N__31529\
        );

    \I__7142\ : Span4Mux_s2_h
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__31526\,
            I => \N__31523\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__31523\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_1\
        );

    \I__7139\ : CascadeMux
    port map (
            O => \N__31520\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\
        );

    \I__7138\ : CascadeMux
    port map (
            O => \N__31517\,
            I => \N__31514\
        );

    \I__7137\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31511\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31507\
        );

    \I__7135\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31504\
        );

    \I__7134\ : Span4Mux_h
    port map (
            O => \N__31507\,
            I => \N__31499\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__31504\,
            I => \N__31499\
        );

    \I__7132\ : Span4Mux_s3_h
    port map (
            O => \N__31499\,
            I => \N__31496\
        );

    \I__7131\ : Span4Mux_v
    port map (
            O => \N__31496\,
            I => \N__31493\
        );

    \I__7130\ : Odrv4
    port map (
            O => \N__31493\,
            I => \VPP_VDDQ.count_2_1_1\
        );

    \I__7129\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31487\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__31487\,
            I => \VPP_VDDQ.curr_state_2_0_1\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__31484\,
            I => \N__31480\
        );

    \I__7126\ : CascadeMux
    port map (
            O => \N__31483\,
            I => \N__31477\
        );

    \I__7125\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31474\
        );

    \I__7124\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31471\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__31474\,
            I => \N__31468\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__31471\,
            I => \N__31465\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__31468\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__31465\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\
        );

    \I__7119\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31454\
        );

    \I__7118\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31454\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__31454\,
            I => \VPP_VDDQ.count_2_1_2\
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__31451\,
            I => \VPP_VDDQ.count_2_1_3_cascade_\
        );

    \I__7115\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31444\
        );

    \I__7114\ : InMux
    port map (
            O => \N__31447\,
            I => \N__31441\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__31444\,
            I => \N__31438\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__31441\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__7111\ : Odrv4
    port map (
            O => \N__31438\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__7110\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31430\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__31430\,
            I => \VPP_VDDQ.N_385\
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__31427\,
            I => \VPP_VDDQ.N_385_cascade_\
        );

    \I__7107\ : InMux
    port map (
            O => \N__31424\,
            I => \N__31420\
        );

    \I__7106\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31417\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__31420\,
            I => \N__31414\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__31417\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__7103\ : Odrv12
    port map (
            O => \N__31414\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__31409\,
            I => \N__31406\
        );

    \I__7101\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31400\
        );

    \I__7100\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31400\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__31400\,
            I => \N__31397\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__31397\,
            I => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\
        );

    \I__7097\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31391\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__31391\,
            I => \POWERLED.count_clk_0_11\
        );

    \I__7095\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31385\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__31385\,
            I => \POWERLED.count_clk_0_12\
        );

    \I__7093\ : CascadeMux
    port map (
            O => \N__31382\,
            I => \N__31379\
        );

    \I__7092\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31373\
        );

    \I__7091\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31373\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31370\
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__31370\,
            I => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\
        );

    \I__7088\ : InMux
    port map (
            O => \N__31367\,
            I => \N__31363\
        );

    \I__7087\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31360\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__31363\,
            I => \N__31355\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31360\,
            I => \N__31355\
        );

    \I__7084\ : Odrv12
    port map (
            O => \N__31355\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__7083\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31349\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31342\
        );

    \I__7081\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31339\
        );

    \I__7080\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31332\
        );

    \I__7079\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31332\
        );

    \I__7078\ : InMux
    port map (
            O => \N__31345\,
            I => \N__31332\
        );

    \I__7077\ : Span4Mux_h
    port map (
            O => \N__31342\,
            I => \N__31329\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__31339\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__31332\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__31329\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31304\
        );

    \I__7072\ : InMux
    port map (
            O => \N__31321\,
            I => \N__31304\
        );

    \I__7071\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31299\
        );

    \I__7070\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31299\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31290\
        );

    \I__7068\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31290\
        );

    \I__7067\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31290\
        );

    \I__7066\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31290\
        );

    \I__7065\ : CascadeMux
    port map (
            O => \N__31314\,
            I => \N__31287\
        );

    \I__7064\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31272\
        );

    \I__7063\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31272\
        );

    \I__7062\ : InMux
    port map (
            O => \N__31311\,
            I => \N__31272\
        );

    \I__7061\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31272\
        );

    \I__7060\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31272\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31265\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__31299\,
            I => \N__31265\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__31290\,
            I => \N__31265\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31254\
        );

    \I__7055\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31254\
        );

    \I__7054\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31254\
        );

    \I__7053\ : InMux
    port map (
            O => \N__31284\,
            I => \N__31254\
        );

    \I__7052\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31254\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__31272\,
            I => \N__31244\
        );

    \I__7050\ : Span4Mux_v
    port map (
            O => \N__31265\,
            I => \N__31244\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31244\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31237\
        );

    \I__7047\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31237\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31251\,
            I => \N__31237\
        );

    \I__7045\ : Span4Mux_s3_h
    port map (
            O => \N__31244\,
            I => \N__31234\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__31237\,
            I => \POWERLED.func_state_RNICAC53_0_0\
        );

    \I__7043\ : Odrv4
    port map (
            O => \N__31234\,
            I => \POWERLED.func_state_RNICAC53_0_0\
        );

    \I__7042\ : InMux
    port map (
            O => \N__31229\,
            I => \N__31226\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__31226\,
            I => \POWERLED.count_clk_0_1\
        );

    \I__7040\ : CEMux
    port map (
            O => \N__31223\,
            I => \N__31220\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__31220\,
            I => \N__31214\
        );

    \I__7038\ : CEMux
    port map (
            O => \N__31219\,
            I => \N__31211\
        );

    \I__7037\ : CEMux
    port map (
            O => \N__31218\,
            I => \N__31208\
        );

    \I__7036\ : CEMux
    port map (
            O => \N__31217\,
            I => \N__31198\
        );

    \I__7035\ : Span4Mux_v
    port map (
            O => \N__31214\,
            I => \N__31193\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__31211\,
            I => \N__31193\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31188\
        );

    \I__7032\ : CEMux
    port map (
            O => \N__31207\,
            I => \N__31183\
        );

    \I__7031\ : InMux
    port map (
            O => \N__31206\,
            I => \N__31183\
        );

    \I__7030\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31174\
        );

    \I__7029\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31174\
        );

    \I__7028\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31174\
        );

    \I__7027\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31174\
        );

    \I__7026\ : CEMux
    port map (
            O => \N__31201\,
            I => \N__31171\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__31198\,
            I => \N__31166\
        );

    \I__7024\ : Span4Mux_s2_h
    port map (
            O => \N__31193\,
            I => \N__31166\
        );

    \I__7023\ : InMux
    port map (
            O => \N__31192\,
            I => \N__31163\
        );

    \I__7022\ : CascadeMux
    port map (
            O => \N__31191\,
            I => \N__31157\
        );

    \I__7021\ : Span4Mux_v
    port map (
            O => \N__31188\,
            I => \N__31152\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31152\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__31174\,
            I => \N__31149\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__31171\,
            I => \N__31136\
        );

    \I__7017\ : Span4Mux_h
    port map (
            O => \N__31166\,
            I => \N__31136\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__31163\,
            I => \N__31136\
        );

    \I__7015\ : InMux
    port map (
            O => \N__31162\,
            I => \N__31131\
        );

    \I__7014\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31131\
        );

    \I__7013\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31126\
        );

    \I__7012\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31126\
        );

    \I__7011\ : Span4Mux_h
    port map (
            O => \N__31152\,
            I => \N__31123\
        );

    \I__7010\ : Span4Mux_h
    port map (
            O => \N__31149\,
            I => \N__31120\
        );

    \I__7009\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31107\
        );

    \I__7008\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31107\
        );

    \I__7007\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31107\
        );

    \I__7006\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31107\
        );

    \I__7005\ : InMux
    port map (
            O => \N__31144\,
            I => \N__31107\
        );

    \I__7004\ : InMux
    port map (
            O => \N__31143\,
            I => \N__31107\
        );

    \I__7003\ : Sp12to4
    port map (
            O => \N__31136\,
            I => \N__31100\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__31131\,
            I => \N__31100\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__31126\,
            I => \N__31100\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__31123\,
            I => \POWERLED.count_clk_en\
        );

    \I__6999\ : Odrv4
    port map (
            O => \N__31120\,
            I => \POWERLED.count_clk_en\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__31107\,
            I => \POWERLED.count_clk_en\
        );

    \I__6997\ : Odrv12
    port map (
            O => \N__31100\,
            I => \POWERLED.count_clk_en\
        );

    \I__6996\ : InMux
    port map (
            O => \N__31091\,
            I => \N__31088\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__31088\,
            I => \POWERLED.count_clk_RNIZ0Z_0\
        );

    \I__6994\ : CascadeMux
    port map (
            O => \N__31085\,
            I => \N__31082\
        );

    \I__6993\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__31079\,
            I => \N__31073\
        );

    \I__6991\ : InMux
    port map (
            O => \N__31078\,
            I => \N__31070\
        );

    \I__6990\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31067\
        );

    \I__6989\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31064\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__31073\,
            I => \N__31061\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__31070\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__31067\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__31064\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__31061\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6983\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31048\
        );

    \I__6982\ : InMux
    port map (
            O => \N__31051\,
            I => \N__31045\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__31048\,
            I => \POWERLED.N_163\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__31045\,
            I => \POWERLED.N_163\
        );

    \I__6979\ : InMux
    port map (
            O => \N__31040\,
            I => \N__31036\
        );

    \I__6978\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31033\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__31036\,
            I => \N__31029\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__31033\,
            I => \N__31026\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31023\
        );

    \I__6974\ : Span4Mux_s3_h
    port map (
            O => \N__31029\,
            I => \N__31020\
        );

    \I__6973\ : Span4Mux_s2_h
    port map (
            O => \N__31026\,
            I => \N__31017\
        );

    \I__6972\ : InMux
    port map (
            O => \N__31023\,
            I => \N__31014\
        );

    \I__6971\ : Odrv4
    port map (
            O => \N__31020\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__6970\ : Odrv4
    port map (
            O => \N__31017\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__31014\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__6968\ : CascadeMux
    port map (
            O => \N__31007\,
            I => \POWERLED.count_clkZ0Z_1_cascade_\
        );

    \I__6967\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30999\
        );

    \I__6966\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30996\
        );

    \I__6965\ : CascadeMux
    port map (
            O => \N__31002\,
            I => \N__30993\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30990\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30987\
        );

    \I__6962\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30984\
        );

    \I__6961\ : Span4Mux_v
    port map (
            O => \N__30990\,
            I => \N__30981\
        );

    \I__6960\ : Span4Mux_s2_h
    port map (
            O => \N__30987\,
            I => \N__30978\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30975\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__30981\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__6957\ : Odrv4
    port map (
            O => \N__30978\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__6956\ : Odrv4
    port map (
            O => \N__30975\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__6955\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30962\
        );

    \I__6954\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30962\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__30962\,
            I => \POWERLED.N_176\
        );

    \I__6952\ : CascadeMux
    port map (
            O => \N__30959\,
            I => \POWERLED.count_offZ0Z_0_cascade_\
        );

    \I__6951\ : InMux
    port map (
            O => \N__30956\,
            I => \N__30953\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__30953\,
            I => \POWERLED.count_off_0_0\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__30950\,
            I => \N__30947\
        );

    \I__6948\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30943\
        );

    \I__6947\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30940\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__30943\,
            I => \N__30935\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__30940\,
            I => \N__30935\
        );

    \I__6944\ : Odrv4
    port map (
            O => \N__30935\,
            I => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\
        );

    \I__6943\ : CascadeMux
    port map (
            O => \N__30932\,
            I => \N__30926\
        );

    \I__6942\ : InMux
    port map (
            O => \N__30931\,
            I => \N__30903\
        );

    \I__6941\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30903\
        );

    \I__6940\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30903\
        );

    \I__6939\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30894\
        );

    \I__6938\ : InMux
    port map (
            O => \N__30925\,
            I => \N__30894\
        );

    \I__6937\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30894\
        );

    \I__6936\ : InMux
    port map (
            O => \N__30923\,
            I => \N__30894\
        );

    \I__6935\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30889\
        );

    \I__6934\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30889\
        );

    \I__6933\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30877\
        );

    \I__6932\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30877\
        );

    \I__6931\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30877\
        );

    \I__6930\ : InMux
    port map (
            O => \N__30917\,
            I => \N__30877\
        );

    \I__6929\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30877\
        );

    \I__6928\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30864\
        );

    \I__6927\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30864\
        );

    \I__6926\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30864\
        );

    \I__6925\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30864\
        );

    \I__6924\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30864\
        );

    \I__6923\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30864\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__30903\,
            I => \N__30848\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__30894\,
            I => \N__30848\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__30889\,
            I => \N__30845\
        );

    \I__6919\ : InMux
    port map (
            O => \N__30888\,
            I => \N__30842\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__30877\,
            I => \N__30839\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__30864\,
            I => \N__30836\
        );

    \I__6916\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30823\
        );

    \I__6915\ : InMux
    port map (
            O => \N__30862\,
            I => \N__30823\
        );

    \I__6914\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30823\
        );

    \I__6913\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30823\
        );

    \I__6912\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30823\
        );

    \I__6911\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30823\
        );

    \I__6910\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30812\
        );

    \I__6909\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30812\
        );

    \I__6908\ : InMux
    port map (
            O => \N__30855\,
            I => \N__30812\
        );

    \I__6907\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30812\
        );

    \I__6906\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30812\
        );

    \I__6905\ : Span4Mux_h
    port map (
            O => \N__30848\,
            I => \N__30809\
        );

    \I__6904\ : Odrv12
    port map (
            O => \N__30845\,
            I => \POWERLED.N_116\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__30842\,
            I => \POWERLED.N_116\
        );

    \I__6902\ : Odrv4
    port map (
            O => \N__30839\,
            I => \POWERLED.N_116\
        );

    \I__6901\ : Odrv4
    port map (
            O => \N__30836\,
            I => \POWERLED.N_116\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__30823\,
            I => \POWERLED.N_116\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__30812\,
            I => \POWERLED.N_116\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__30809\,
            I => \POWERLED.N_116\
        );

    \I__6897\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__30791\,
            I => \POWERLED.count_off_0_4\
        );

    \I__6895\ : CEMux
    port map (
            O => \N__30788\,
            I => \N__30779\
        );

    \I__6894\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30768\
        );

    \I__6893\ : CEMux
    port map (
            O => \N__30786\,
            I => \N__30768\
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__30785\,
            I => \N__30762\
        );

    \I__6891\ : CascadeMux
    port map (
            O => \N__30784\,
            I => \N__30758\
        );

    \I__6890\ : CEMux
    port map (
            O => \N__30783\,
            I => \N__30748\
        );

    \I__6889\ : CEMux
    port map (
            O => \N__30782\,
            I => \N__30745\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30742\
        );

    \I__6887\ : CascadeMux
    port map (
            O => \N__30778\,
            I => \N__30739\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__30777\,
            I => \N__30736\
        );

    \I__6885\ : InMux
    port map (
            O => \N__30776\,
            I => \N__30727\
        );

    \I__6884\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30727\
        );

    \I__6883\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30727\
        );

    \I__6882\ : InMux
    port map (
            O => \N__30773\,
            I => \N__30724\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__30768\,
            I => \N__30721\
        );

    \I__6880\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30716\
        );

    \I__6879\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30716\
        );

    \I__6878\ : CEMux
    port map (
            O => \N__30765\,
            I => \N__30711\
        );

    \I__6877\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30704\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30704\
        );

    \I__6875\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30704\
        );

    \I__6874\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30695\
        );

    \I__6873\ : InMux
    port map (
            O => \N__30756\,
            I => \N__30695\
        );

    \I__6872\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30695\
        );

    \I__6871\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30695\
        );

    \I__6870\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30688\
        );

    \I__6869\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30688\
        );

    \I__6868\ : CEMux
    port map (
            O => \N__30751\,
            I => \N__30688\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__30748\,
            I => \N__30683\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__30745\,
            I => \N__30683\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__30742\,
            I => \N__30680\
        );

    \I__6864\ : InMux
    port map (
            O => \N__30739\,
            I => \N__30671\
        );

    \I__6863\ : InMux
    port map (
            O => \N__30736\,
            I => \N__30671\
        );

    \I__6862\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30671\
        );

    \I__6861\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30671\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__30727\,
            I => \N__30668\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__30724\,
            I => \N__30665\
        );

    \I__6858\ : Span4Mux_v
    port map (
            O => \N__30721\,
            I => \N__30662\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__30716\,
            I => \N__30659\
        );

    \I__6856\ : InMux
    port map (
            O => \N__30715\,
            I => \N__30654\
        );

    \I__6855\ : InMux
    port map (
            O => \N__30714\,
            I => \N__30654\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__30711\,
            I => \N__30649\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__30704\,
            I => \N__30649\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30646\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__30688\,
            I => \N__30643\
        );

    \I__6850\ : Span4Mux_s3_v
    port map (
            O => \N__30683\,
            I => \N__30632\
        );

    \I__6849\ : Span4Mux_s0_h
    port map (
            O => \N__30680\,
            I => \N__30632\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__30671\,
            I => \N__30632\
        );

    \I__6847\ : Span4Mux_s3_v
    port map (
            O => \N__30668\,
            I => \N__30632\
        );

    \I__6846\ : Span4Mux_v
    port map (
            O => \N__30665\,
            I => \N__30632\
        );

    \I__6845\ : Span4Mux_s1_h
    port map (
            O => \N__30662\,
            I => \N__30623\
        );

    \I__6844\ : Span4Mux_v
    port map (
            O => \N__30659\,
            I => \N__30623\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__30654\,
            I => \N__30623\
        );

    \I__6842\ : Span4Mux_s3_v
    port map (
            O => \N__30649\,
            I => \N__30623\
        );

    \I__6841\ : Span4Mux_s3_h
    port map (
            O => \N__30646\,
            I => \N__30620\
        );

    \I__6840\ : Odrv12
    port map (
            O => \N__30643\,
            I => \POWERLED.count_off_enZ0\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__30632\,
            I => \POWERLED.count_off_enZ0\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__30623\,
            I => \POWERLED.count_off_enZ0\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__30620\,
            I => \POWERLED.count_off_enZ0\
        );

    \I__6836\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30608\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__30608\,
            I => \N__30605\
        );

    \I__6834\ : Span12Mux_v
    port map (
            O => \N__30605\,
            I => \N__30602\
        );

    \I__6833\ : Odrv12
    port map (
            O => \N__30602\,
            I => v33s_ok
        );

    \I__6832\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30596\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__30596\,
            I => \N__30593\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__30593\,
            I => \N__30590\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__30590\,
            I => vccst_cpu_ok
        );

    \I__6828\ : CascadeMux
    port map (
            O => \N__30587\,
            I => \N__30580\
        );

    \I__6827\ : CascadeMux
    port map (
            O => \N__30586\,
            I => \N__30577\
        );

    \I__6826\ : InMux
    port map (
            O => \N__30585\,
            I => \N__30571\
        );

    \I__6825\ : InMux
    port map (
            O => \N__30584\,
            I => \N__30571\
        );

    \I__6824\ : InMux
    port map (
            O => \N__30583\,
            I => \N__30568\
        );

    \I__6823\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30565\
        );

    \I__6822\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30562\
        );

    \I__6821\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30559\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30556\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__30568\,
            I => \N__30551\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30543\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__30562\,
            I => \N__30536\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30536\
        );

    \I__6815\ : Span4Mux_s3_h
    port map (
            O => \N__30556\,
            I => \N__30536\
        );

    \I__6814\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30531\
        );

    \I__6813\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30531\
        );

    \I__6812\ : Span4Mux_v
    port map (
            O => \N__30551\,
            I => \N__30528\
        );

    \I__6811\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30525\
        );

    \I__6810\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30516\
        );

    \I__6809\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30516\
        );

    \I__6808\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30510\
        );

    \I__6807\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30510\
        );

    \I__6806\ : Span4Mux_v
    port map (
            O => \N__30543\,
            I => \N__30506\
        );

    \I__6805\ : Span4Mux_h
    port map (
            O => \N__30536\,
            I => \N__30501\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__30531\,
            I => \N__30501\
        );

    \I__6803\ : Span4Mux_v
    port map (
            O => \N__30528\,
            I => \N__30498\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__30525\,
            I => \N__30495\
        );

    \I__6801\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30488\
        );

    \I__6800\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30488\
        );

    \I__6799\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30488\
        );

    \I__6798\ : CascadeMux
    port map (
            O => \N__30521\,
            I => \N__30485\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30479\
        );

    \I__6796\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30476\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__30510\,
            I => \N__30473\
        );

    \I__6794\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30470\
        );

    \I__6793\ : Span4Mux_h
    port map (
            O => \N__30506\,
            I => \N__30465\
        );

    \I__6792\ : Span4Mux_v
    port map (
            O => \N__30501\,
            I => \N__30465\
        );

    \I__6791\ : Span4Mux_h
    port map (
            O => \N__30498\,
            I => \N__30458\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__30495\,
            I => \N__30458\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__30488\,
            I => \N__30458\
        );

    \I__6788\ : InMux
    port map (
            O => \N__30485\,
            I => \N__30453\
        );

    \I__6787\ : InMux
    port map (
            O => \N__30484\,
            I => \N__30453\
        );

    \I__6786\ : InMux
    port map (
            O => \N__30483\,
            I => \N__30448\
        );

    \I__6785\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30448\
        );

    \I__6784\ : Span12Mux_s7_h
    port map (
            O => \N__30479\,
            I => \N__30441\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__30476\,
            I => \N__30441\
        );

    \I__6782\ : Span12Mux_s4_h
    port map (
            O => \N__30473\,
            I => \N__30441\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__30470\,
            I => slp_s3n_signal
        );

    \I__6780\ : Odrv4
    port map (
            O => \N__30465\,
            I => slp_s3n_signal
        );

    \I__6779\ : Odrv4
    port map (
            O => \N__30458\,
            I => slp_s3n_signal
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__30453\,
            I => slp_s3n_signal
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__30448\,
            I => slp_s3n_signal
        );

    \I__6776\ : Odrv12
    port map (
            O => \N__30441\,
            I => slp_s3n_signal
        );

    \I__6775\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30425\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__30425\,
            I => \N__30422\
        );

    \I__6773\ : Span4Mux_s3_h
    port map (
            O => \N__30422\,
            I => \N__30419\
        );

    \I__6772\ : Span4Mux_h
    port map (
            O => \N__30419\,
            I => \N__30412\
        );

    \I__6771\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30403\
        );

    \I__6770\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30403\
        );

    \I__6769\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30403\
        );

    \I__6768\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30403\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__30412\,
            I => rsmrst_pwrgd_signal
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__30403\,
            I => rsmrst_pwrgd_signal
        );

    \I__6765\ : InMux
    port map (
            O => \N__30398\,
            I => \N__30395\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__30395\,
            I => v5s_ok
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__30392\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\
        );

    \I__6762\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30386\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30386\,
            I => \N__30382\
        );

    \I__6760\ : IoInMux
    port map (
            O => \N__30385\,
            I => \N__30379\
        );

    \I__6759\ : Span4Mux_v
    port map (
            O => \N__30382\,
            I => \N__30376\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__30379\,
            I => \N__30373\
        );

    \I__6757\ : Sp12to4
    port map (
            O => \N__30376\,
            I => \N__30370\
        );

    \I__6756\ : Span4Mux_s0_h
    port map (
            O => \N__30373\,
            I => \N__30367\
        );

    \I__6755\ : Span12Mux_s4_h
    port map (
            O => \N__30370\,
            I => \N__30364\
        );

    \I__6754\ : Span4Mux_v
    port map (
            O => \N__30367\,
            I => \N__30361\
        );

    \I__6753\ : Odrv12
    port map (
            O => \N__30364\,
            I => dsw_pwrok
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__30361\,
            I => dsw_pwrok
        );

    \I__6751\ : IoInMux
    port map (
            O => \N__30356\,
            I => \N__30353\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__6749\ : Span4Mux_s1_v
    port map (
            O => \N__30350\,
            I => \N__30347\
        );

    \I__6748\ : Span4Mux_v
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__6747\ : Span4Mux_v
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__6746\ : Odrv4
    port map (
            O => \N__30341\,
            I => vccin_en
        );

    \I__6745\ : CascadeMux
    port map (
            O => \N__30338\,
            I => \VPP_VDDQ.delayed_vddq_okZ0_cascade_\
        );

    \I__6744\ : IoInMux
    port map (
            O => \N__30335\,
            I => \N__30332\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__30332\,
            I => \N__30329\
        );

    \I__6742\ : Span4Mux_s2_h
    port map (
            O => \N__30329\,
            I => \N__30325\
        );

    \I__6741\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30322\
        );

    \I__6740\ : Span4Mux_v
    port map (
            O => \N__30325\,
            I => \N__30319\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__30322\,
            I => \N__30316\
        );

    \I__6738\ : Span4Mux_v
    port map (
            O => \N__30319\,
            I => \N__30311\
        );

    \I__6737\ : Span4Mux_s2_h
    port map (
            O => \N__30316\,
            I => \N__30311\
        );

    \I__6736\ : Span4Mux_h
    port map (
            O => \N__30311\,
            I => \N__30307\
        );

    \I__6735\ : CascadeMux
    port map (
            O => \N__30310\,
            I => \N__30303\
        );

    \I__6734\ : Span4Mux_h
    port map (
            O => \N__30307\,
            I => \N__30299\
        );

    \I__6733\ : IoInMux
    port map (
            O => \N__30306\,
            I => \N__30296\
        );

    \I__6732\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30293\
        );

    \I__6731\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30290\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__30299\,
            I => \N__30287\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__30296\,
            I => \N__30280\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30280\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__30290\,
            I => \N__30280\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__30287\,
            I => pch_pwrok
        );

    \I__6725\ : Odrv12
    port map (
            O => \N__30280\,
            I => pch_pwrok
        );

    \I__6724\ : IoInMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__6722\ : IoSpan4Mux
    port map (
            O => \N__30269\,
            I => \N__30266\
        );

    \I__6721\ : Span4Mux_s2_v
    port map (
            O => \N__30266\,
            I => \N__30263\
        );

    \I__6720\ : Span4Mux_v
    port map (
            O => \N__30263\,
            I => \N__30260\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__30257\,
            I => vccst_pwrgd
        );

    \I__6717\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30251\,
            I => \VPP_VDDQ.delayed_vddq_ok_en\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__30248\,
            I => \VPP_VDDQ.delayed_vddq_ok_en_cascade_\
        );

    \I__6714\ : CascadeMux
    port map (
            O => \N__30245\,
            I => \N__30242\
        );

    \I__6713\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30236\
        );

    \I__6712\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30236\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__30236\,
            I => \N__30233\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__30233\,
            I => \VPP_VDDQ.delayed_vddq_ok_0\
        );

    \I__6709\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30218\
        );

    \I__6708\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30218\
        );

    \I__6707\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30218\
        );

    \I__6706\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30218\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__30218\,
            I => \VPP_VDDQ.N_53\
        );

    \I__6704\ : SRMux
    port map (
            O => \N__30215\,
            I => \N__30212\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__30212\,
            I => \N__30209\
        );

    \I__6702\ : Sp12to4
    port map (
            O => \N__30209\,
            I => \N__30206\
        );

    \I__6701\ : Odrv12
    port map (
            O => \N__30206\,
            I => \VPP_VDDQ.N_53_i\
        );

    \I__6700\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30200\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__30200\,
            I => \N__30196\
        );

    \I__6698\ : InMux
    port map (
            O => \N__30199\,
            I => \N__30193\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__30196\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__30193\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__6695\ : InMux
    port map (
            O => \N__30188\,
            I => \POWERLED.un3_count_off_1_cry_14\
        );

    \I__6694\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30179\
        );

    \I__6693\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30179\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__30179\,
            I => \N__30176\
        );

    \I__6691\ : Odrv4
    port map (
            O => \N__30176\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNIB6QDZ0\
        );

    \I__6690\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30170\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__6688\ : Span4Mux_v
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__6687\ : Odrv4
    port map (
            O => \N__30164\,
            I => \POWERLED.count_off_0_14\
        );

    \I__6686\ : CascadeMux
    port map (
            O => \N__30161\,
            I => \N__30157\
        );

    \I__6685\ : InMux
    port map (
            O => \N__30160\,
            I => \N__30154\
        );

    \I__6684\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30151\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30148\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__30151\,
            I => \POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__30148\,
            I => \POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0\
        );

    \I__6680\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30136\
        );

    \I__6678\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30133\
        );

    \I__6677\ : Odrv12
    port map (
            O => \N__30136\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__30133\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__6675\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30125\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__30125\,
            I => \N__30122\
        );

    \I__6673\ : Odrv12
    port map (
            O => \N__30122\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__30119\,
            I => \POWERLED.count_offZ0Z_4_cascade_\
        );

    \I__6671\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30113\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__30113\,
            I => \N__30110\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__30110\,
            I => \POWERLED.un34_clk_100khz_2\
        );

    \I__6668\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30101\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30101\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__30098\,
            I => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\
        );

    \I__6664\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30092\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__30092\,
            I => \POWERLED.count_off_1_3\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__30089\,
            I => \POWERLED.count_off_1_3_cascade_\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30080\
        );

    \I__6660\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30080\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__30080\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__6658\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30074\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__30074\,
            I => \N__30071\
        );

    \I__6656\ : Odrv12
    port map (
            O => \N__30071\,
            I => \POWERLED.un3_count_off_1_axb_3\
        );

    \I__6655\ : CascadeMux
    port map (
            O => \N__30068\,
            I => \N__30062\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__30067\,
            I => \N__30059\
        );

    \I__6653\ : InMux
    port map (
            O => \N__30066\,
            I => \N__30054\
        );

    \I__6652\ : InMux
    port map (
            O => \N__30065\,
            I => \N__30054\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30051\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30048\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__30054\,
            I => \N__30043\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__30051\,
            I => \N__30043\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__30048\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__6646\ : Odrv4
    port map (
            O => \N__30043\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__6645\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__30035\,
            I => \POWERLED.un3_count_off_1_axb_7\
        );

    \I__6643\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30026\
        );

    \I__6642\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30026\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__30026\,
            I => \POWERLED.un3_count_off_1_cry_6_c_RNISH5FZ0\
        );

    \I__6640\ : InMux
    port map (
            O => \N__30023\,
            I => \POWERLED.un3_count_off_1_cry_6\
        );

    \I__6639\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30017\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__30017\,
            I => \N__30013\
        );

    \I__6637\ : InMux
    port map (
            O => \N__30016\,
            I => \N__30010\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__30013\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__30010\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__6634\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29999\
        );

    \I__6633\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29999\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__29999\,
            I => \POWERLED.un3_count_off_1_cry_7_c_RNITJ6FZ0\
        );

    \I__6631\ : InMux
    port map (
            O => \N__29996\,
            I => \POWERLED.un3_count_off_1_cry_7\
        );

    \I__6630\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29990\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29987\
        );

    \I__6628\ : Span4Mux_s2_h
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__6627\ : Odrv4
    port map (
            O => \N__29984\,
            I => \POWERLED.un3_count_off_1_axb_9\
        );

    \I__6626\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29975\
        );

    \I__6625\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29975\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__6623\ : Span4Mux_v
    port map (
            O => \N__29972\,
            I => \N__29969\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__29969\,
            I => \POWERLED.un3_count_off_1_cry_8_c_RNIUL7FZ0\
        );

    \I__6621\ : InMux
    port map (
            O => \N__29966\,
            I => \bfn_12_5_0_\
        );

    \I__6620\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29960\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__29960\,
            I => \N__29957\
        );

    \I__6618\ : Span4Mux_v
    port map (
            O => \N__29957\,
            I => \N__29954\
        );

    \I__6617\ : Sp12to4
    port map (
            O => \N__29954\,
            I => \N__29951\
        );

    \I__6616\ : Odrv12
    port map (
            O => \N__29951\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__6614\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29939\
        );

    \I__6613\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29939\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__6611\ : Span4Mux_v
    port map (
            O => \N__29936\,
            I => \N__29933\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__29933\,
            I => \POWERLED.un3_count_off_1_cry_9_c_RNIVN8FZ0\
        );

    \I__6609\ : InMux
    port map (
            O => \N__29930\,
            I => \POWERLED.un3_count_off_1_cry_9\
        );

    \I__6608\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29924\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__29924\,
            I => \POWERLED.un3_count_off_1_axb_11\
        );

    \I__6606\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29915\
        );

    \I__6605\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29915\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__29915\,
            I => \POWERLED.un3_count_off_1_cry_10_c_RNI7ULDZ0\
        );

    \I__6603\ : InMux
    port map (
            O => \N__29912\,
            I => \POWERLED.un3_count_off_1_cry_10\
        );

    \I__6602\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29906\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__29906\,
            I => \N__29902\
        );

    \I__6600\ : InMux
    port map (
            O => \N__29905\,
            I => \N__29899\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__29902\,
            I => \N__29896\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__29899\,
            I => \N__29893\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__29896\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__6596\ : Odrv4
    port map (
            O => \N__29893\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__29888\,
            I => \N__29885\
        );

    \I__6594\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29879\
        );

    \I__6593\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29879\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__29879\,
            I => \N__29876\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__29876\,
            I => \POWERLED.un3_count_off_1_cry_11_c_RNI80NDZ0\
        );

    \I__6590\ : InMux
    port map (
            O => \N__29873\,
            I => \POWERLED.un3_count_off_1_cry_11\
        );

    \I__6589\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__29867\,
            I => \N__29864\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__29864\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__6586\ : CascadeMux
    port map (
            O => \N__29861\,
            I => \N__29858\
        );

    \I__6585\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29852\
        );

    \I__6584\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29852\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29849\
        );

    \I__6582\ : Odrv12
    port map (
            O => \N__29849\,
            I => \POWERLED.un3_count_off_1_cry_12_c_RNI92ODZ0\
        );

    \I__6581\ : InMux
    port map (
            O => \N__29846\,
            I => \POWERLED.un3_count_off_1_cry_12\
        );

    \I__6580\ : InMux
    port map (
            O => \N__29843\,
            I => \POWERLED.un3_count_off_1_cry_13\
        );

    \I__6579\ : InMux
    port map (
            O => \N__29840\,
            I => \N__29837\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__29837\,
            I => \POWERLED.count_off_0_13\
        );

    \I__6577\ : CascadeMux
    port map (
            O => \N__29834\,
            I => \POWERLED.count_offZ0Z_13_cascade_\
        );

    \I__6576\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29828\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__6574\ : Span4Mux_h
    port map (
            O => \N__29825\,
            I => \N__29822\
        );

    \I__6573\ : Odrv4
    port map (
            O => \N__29822\,
            I => \POWERLED.un34_clk_100khz_11\
        );

    \I__6572\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29814\
        );

    \I__6571\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29811\
        );

    \I__6570\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29808\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__29814\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__29811\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__29808\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__6566\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__29798\,
            I => \POWERLED.un3_count_off_1_axb_2\
        );

    \I__6564\ : InMux
    port map (
            O => \N__29795\,
            I => \N__29789\
        );

    \I__6563\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29789\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__29789\,
            I => \POWERLED.un3_count_off_1_cry_1_c_RNIN70FZ0\
        );

    \I__6561\ : InMux
    port map (
            O => \N__29786\,
            I => \POWERLED.un3_count_off_1_cry_1\
        );

    \I__6560\ : InMux
    port map (
            O => \N__29783\,
            I => \POWERLED.un3_count_off_1_cry_2\
        );

    \I__6559\ : InMux
    port map (
            O => \N__29780\,
            I => \POWERLED.un3_count_off_1_cry_3\
        );

    \I__6558\ : CascadeMux
    port map (
            O => \N__29777\,
            I => \N__29773\
        );

    \I__6557\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29770\
        );

    \I__6556\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29767\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__29770\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__29767\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__6553\ : CascadeMux
    port map (
            O => \N__29762\,
            I => \N__29758\
        );

    \I__6552\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29753\
        );

    \I__6551\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29753\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__29753\,
            I => \POWERLED.un3_count_off_1_cry_4_c_RNIQD3FZ0\
        );

    \I__6549\ : InMux
    port map (
            O => \N__29750\,
            I => \POWERLED.un3_count_off_1_cry_4\
        );

    \I__6548\ : InMux
    port map (
            O => \N__29747\,
            I => \N__29744\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__29744\,
            I => \POWERLED.un3_count_off_1_axb_6\
        );

    \I__6546\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29737\
        );

    \I__6545\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29734\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__29737\,
            I => \POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__29734\,
            I => \POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0\
        );

    \I__6542\ : InMux
    port map (
            O => \N__29729\,
            I => \POWERLED.un3_count_off_1_cry_5\
        );

    \I__6541\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29722\
        );

    \I__6540\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29719\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__29722\,
            I => \VPP_VDDQ.N_186\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__29719\,
            I => \VPP_VDDQ.N_186\
        );

    \I__6537\ : CascadeMux
    port map (
            O => \N__29714\,
            I => \N__29711\
        );

    \I__6536\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29708\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__29708\,
            I => \VPP_VDDQ.N_214\
        );

    \I__6534\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29701\
        );

    \I__6533\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29695\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__29698\,
            I => \N__29692\
        );

    \I__6530\ : Span4Mux_v
    port map (
            O => \N__29695\,
            I => \N__29689\
        );

    \I__6529\ : Span4Mux_s3_h
    port map (
            O => \N__29692\,
            I => \N__29686\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__29689\,
            I => \VPP_VDDQ.un6_count\
        );

    \I__6527\ : Odrv4
    port map (
            O => \N__29686\,
            I => \VPP_VDDQ.un6_count\
        );

    \I__6526\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29676\
        );

    \I__6525\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29668\
        );

    \I__6524\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29668\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__29676\,
            I => \N__29665\
        );

    \I__6522\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29658\
        );

    \I__6521\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29658\
        );

    \I__6520\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29658\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__29668\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6518\ : Odrv4
    port map (
            O => \N__29665\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__29658\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6516\ : CascadeMux
    port map (
            O => \N__29651\,
            I => \N__29647\
        );

    \I__6515\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29641\
        );

    \I__6514\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29641\
        );

    \I__6513\ : InMux
    port map (
            O => \N__29646\,
            I => \N__29637\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29634\
        );

    \I__6511\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29631\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__29637\,
            I => \VPP_VDDQ.N_360\
        );

    \I__6509\ : Odrv4
    port map (
            O => \N__29634\,
            I => \VPP_VDDQ.N_360\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__29631\,
            I => \VPP_VDDQ.N_360\
        );

    \I__6507\ : CascadeMux
    port map (
            O => \N__29624\,
            I => \N__29621\
        );

    \I__6506\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29611\
        );

    \I__6505\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29611\
        );

    \I__6504\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29608\
        );

    \I__6503\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29601\
        );

    \I__6502\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29601\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29601\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__29611\,
            I => \N__29598\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__29608\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__29601\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__6497\ : Odrv4
    port map (
            O => \N__29598\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__6496\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29530\
        );

    \I__6495\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29530\
        );

    \I__6494\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29530\
        );

    \I__6493\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29530\
        );

    \I__6492\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29521\
        );

    \I__6491\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29521\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29521\
        );

    \I__6489\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29521\
        );

    \I__6488\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29512\
        );

    \I__6487\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29512\
        );

    \I__6486\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29512\
        );

    \I__6485\ : InMux
    port map (
            O => \N__29580\,
            I => \N__29512\
        );

    \I__6484\ : InMux
    port map (
            O => \N__29579\,
            I => \N__29505\
        );

    \I__6483\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29505\
        );

    \I__6482\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29505\
        );

    \I__6481\ : InMux
    port map (
            O => \N__29576\,
            I => \N__29500\
        );

    \I__6480\ : InMux
    port map (
            O => \N__29575\,
            I => \N__29500\
        );

    \I__6479\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29491\
        );

    \I__6478\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29491\
        );

    \I__6477\ : InMux
    port map (
            O => \N__29572\,
            I => \N__29491\
        );

    \I__6476\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29491\
        );

    \I__6475\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29484\
        );

    \I__6474\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29484\
        );

    \I__6473\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29484\
        );

    \I__6472\ : InMux
    port map (
            O => \N__29567\,
            I => \N__29475\
        );

    \I__6471\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29475\
        );

    \I__6470\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29475\
        );

    \I__6469\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29475\
        );

    \I__6468\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29468\
        );

    \I__6467\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29468\
        );

    \I__6466\ : InMux
    port map (
            O => \N__29561\,
            I => \N__29468\
        );

    \I__6465\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29459\
        );

    \I__6464\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29459\
        );

    \I__6463\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29459\
        );

    \I__6462\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29459\
        );

    \I__6461\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29450\
        );

    \I__6460\ : InMux
    port map (
            O => \N__29555\,
            I => \N__29450\
        );

    \I__6459\ : InMux
    port map (
            O => \N__29554\,
            I => \N__29450\
        );

    \I__6458\ : InMux
    port map (
            O => \N__29553\,
            I => \N__29450\
        );

    \I__6457\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29441\
        );

    \I__6456\ : InMux
    port map (
            O => \N__29551\,
            I => \N__29441\
        );

    \I__6455\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29441\
        );

    \I__6454\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29441\
        );

    \I__6453\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29436\
        );

    \I__6452\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29436\
        );

    \I__6451\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29427\
        );

    \I__6450\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29427\
        );

    \I__6449\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29427\
        );

    \I__6448\ : InMux
    port map (
            O => \N__29543\,
            I => \N__29427\
        );

    \I__6447\ : InMux
    port map (
            O => \N__29542\,
            I => \N__29422\
        );

    \I__6446\ : InMux
    port map (
            O => \N__29541\,
            I => \N__29422\
        );

    \I__6445\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29417\
        );

    \I__6444\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29417\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__29530\,
            I => \N__29412\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__29521\,
            I => \N__29409\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__29512\,
            I => \N__29405\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__29505\,
            I => \N__29402\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__29500\,
            I => \N__29398\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__29491\,
            I => \N__29392\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29389\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__29475\,
            I => \N__29386\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__29468\,
            I => \N__29383\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29380\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__29450\,
            I => \N__29377\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29441\,
            I => \N__29374\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__29436\,
            I => \N__29371\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29368\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__29422\,
            I => \N__29365\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__29417\,
            I => \N__29362\
        );

    \I__6427\ : CEMux
    port map (
            O => \N__29416\,
            I => \N__29315\
        );

    \I__6426\ : CEMux
    port map (
            O => \N__29415\,
            I => \N__29315\
        );

    \I__6425\ : Glb2LocalMux
    port map (
            O => \N__29412\,
            I => \N__29315\
        );

    \I__6424\ : Glb2LocalMux
    port map (
            O => \N__29409\,
            I => \N__29315\
        );

    \I__6423\ : CEMux
    port map (
            O => \N__29408\,
            I => \N__29315\
        );

    \I__6422\ : Glb2LocalMux
    port map (
            O => \N__29405\,
            I => \N__29315\
        );

    \I__6421\ : Glb2LocalMux
    port map (
            O => \N__29402\,
            I => \N__29315\
        );

    \I__6420\ : CEMux
    port map (
            O => \N__29401\,
            I => \N__29315\
        );

    \I__6419\ : Glb2LocalMux
    port map (
            O => \N__29398\,
            I => \N__29315\
        );

    \I__6418\ : CEMux
    port map (
            O => \N__29397\,
            I => \N__29315\
        );

    \I__6417\ : CEMux
    port map (
            O => \N__29396\,
            I => \N__29315\
        );

    \I__6416\ : CEMux
    port map (
            O => \N__29395\,
            I => \N__29315\
        );

    \I__6415\ : Glb2LocalMux
    port map (
            O => \N__29392\,
            I => \N__29315\
        );

    \I__6414\ : Glb2LocalMux
    port map (
            O => \N__29389\,
            I => \N__29315\
        );

    \I__6413\ : Glb2LocalMux
    port map (
            O => \N__29386\,
            I => \N__29315\
        );

    \I__6412\ : Glb2LocalMux
    port map (
            O => \N__29383\,
            I => \N__29315\
        );

    \I__6411\ : Glb2LocalMux
    port map (
            O => \N__29380\,
            I => \N__29315\
        );

    \I__6410\ : Glb2LocalMux
    port map (
            O => \N__29377\,
            I => \N__29315\
        );

    \I__6409\ : Glb2LocalMux
    port map (
            O => \N__29374\,
            I => \N__29315\
        );

    \I__6408\ : Glb2LocalMux
    port map (
            O => \N__29371\,
            I => \N__29315\
        );

    \I__6407\ : Glb2LocalMux
    port map (
            O => \N__29368\,
            I => \N__29315\
        );

    \I__6406\ : Glb2LocalMux
    port map (
            O => \N__29365\,
            I => \N__29315\
        );

    \I__6405\ : Glb2LocalMux
    port map (
            O => \N__29362\,
            I => \N__29315\
        );

    \I__6404\ : GlobalMux
    port map (
            O => \N__29315\,
            I => \N__29312\
        );

    \I__6403\ : gio2CtrlBuf
    port map (
            O => \N__29312\,
            I => \N_27_g\
        );

    \I__6402\ : CascadeMux
    port map (
            O => \N__29309\,
            I => \POWERLED.count_off_RNIZ0Z_1_cascade_\
        );

    \I__6401\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29303\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__29303\,
            I => \POWERLED.count_off_0_12\
        );

    \I__6399\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29297\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__29297\,
            I => \POWERLED.count_off_RNIZ0Z_1\
        );

    \I__6397\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29291\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__29291\,
            I => \POWERLED.count_off_0_1\
        );

    \I__6395\ : IoInMux
    port map (
            O => \N__29288\,
            I => \N__29285\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29282\
        );

    \I__6393\ : IoSpan4Mux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__29279\,
            I => vpp_en
        );

    \I__6391\ : InMux
    port map (
            O => \N__29276\,
            I => \N__29273\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__29273\,
            I => \N__29270\
        );

    \I__6389\ : Span4Mux_v
    port map (
            O => \N__29270\,
            I => \N__29264\
        );

    \I__6388\ : IoInMux
    port map (
            O => \N__29269\,
            I => \N__29261\
        );

    \I__6387\ : InMux
    port map (
            O => \N__29268\,
            I => \N__29256\
        );

    \I__6386\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29256\
        );

    \I__6385\ : IoSpan4Mux
    port map (
            O => \N__29264\,
            I => \N__29251\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__29261\,
            I => \N__29251\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29246\
        );

    \I__6382\ : IoSpan4Mux
    port map (
            O => \N__29251\,
            I => \N__29243\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__29250\,
            I => \N__29239\
        );

    \I__6380\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29235\
        );

    \I__6379\ : Span4Mux_s3_v
    port map (
            O => \N__29246\,
            I => \N__29232\
        );

    \I__6378\ : Span4Mux_s0_h
    port map (
            O => \N__29243\,
            I => \N__29228\
        );

    \I__6377\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29225\
        );

    \I__6376\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29222\
        );

    \I__6375\ : CascadeMux
    port map (
            O => \N__29238\,
            I => \N__29219\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29216\
        );

    \I__6373\ : Span4Mux_v
    port map (
            O => \N__29232\,
            I => \N__29213\
        );

    \I__6372\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29210\
        );

    \I__6371\ : Span4Mux_h
    port map (
            O => \N__29228\,
            I => \N__29207\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__29225\,
            I => \N__29202\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__29222\,
            I => \N__29202\
        );

    \I__6368\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29197\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__29216\,
            I => \N__29190\
        );

    \I__6366\ : Span4Mux_v
    port map (
            O => \N__29213\,
            I => \N__29190\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29190\
        );

    \I__6364\ : Span4Mux_h
    port map (
            O => \N__29207\,
            I => \N__29185\
        );

    \I__6363\ : Span4Mux_h
    port map (
            O => \N__29202\,
            I => \N__29185\
        );

    \I__6362\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29182\
        );

    \I__6361\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29179\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29176\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__29190\,
            I => vccst_en
        );

    \I__6358\ : Odrv4
    port map (
            O => \N__29185\,
            I => vccst_en
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__29182\,
            I => vccst_en
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__29179\,
            I => vccst_en
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__29176\,
            I => vccst_en
        );

    \I__6354\ : CascadeMux
    port map (
            O => \N__29165\,
            I => \VPP_VDDQ.N_360_cascade_\
        );

    \I__6353\ : CascadeMux
    port map (
            O => \N__29162\,
            I => \N__29158\
        );

    \I__6352\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29155\
        );

    \I__6351\ : InMux
    port map (
            O => \N__29158\,
            I => \N__29152\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__29155\,
            I => \N__29147\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__29152\,
            I => \N__29147\
        );

    \I__6348\ : Span4Mux_h
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__6347\ : Odrv4
    port map (
            O => \N__29144\,
            I => \VPP_VDDQ.N_264_i\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__29141\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\
        );

    \I__6345\ : InMux
    port map (
            O => \N__29138\,
            I => \N__29132\
        );

    \I__6344\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29132\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__29132\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__6342\ : SRMux
    port map (
            O => \N__29129\,
            I => \N__29125\
        );

    \I__6341\ : SRMux
    port map (
            O => \N__29128\,
            I => \N__29122\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__29125\,
            I => \N__29118\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__29122\,
            I => \N__29115\
        );

    \I__6338\ : SRMux
    port map (
            O => \N__29121\,
            I => \N__29112\
        );

    \I__6337\ : Span4Mux_h
    port map (
            O => \N__29118\,
            I => \N__29109\
        );

    \I__6336\ : Span4Mux_v
    port map (
            O => \N__29115\,
            I => \N__29106\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__29112\,
            I => \N__29103\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__29109\,
            I => \VPP_VDDQ.curr_state_RNITROD7Z0Z_0\
        );

    \I__6333\ : Odrv4
    port map (
            O => \N__29106\,
            I => \VPP_VDDQ.curr_state_RNITROD7Z0Z_0\
        );

    \I__6332\ : Odrv12
    port map (
            O => \N__29103\,
            I => \VPP_VDDQ.curr_state_RNITROD7Z0Z_0\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__29096\,
            I => \VPP_VDDQ.curr_state_RNITROD7Z0Z_0_cascade_\
        );

    \I__6330\ : CEMux
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__29090\,
            I => \N__29087\
        );

    \I__6328\ : Odrv4
    port map (
            O => \N__29087\,
            I => \VPP_VDDQ.N_27_0\
        );

    \I__6327\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29081\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__29081\,
            I => \VPP_VDDQ.N_382\
        );

    \I__6325\ : InMux
    port map (
            O => \N__29078\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__6324\ : InMux
    port map (
            O => \N__29075\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__6323\ : InMux
    port map (
            O => \N__29072\,
            I => \N__29066\
        );

    \I__6322\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29066\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__29066\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__29063\,
            I => \VPP_VDDQ.count_2_1_13_cascade_\
        );

    \I__6319\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29057\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__29057\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__29054\,
            I => \N__29050\
        );

    \I__6316\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29045\
        );

    \I__6315\ : InMux
    port map (
            O => \N__29050\,
            I => \N__29045\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__29045\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__29042\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__29039\,
            I => \N__29035\
        );

    \I__6311\ : InMux
    port map (
            O => \N__29038\,
            I => \N__29030\
        );

    \I__6310\ : InMux
    port map (
            O => \N__29035\,
            I => \N__29030\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__29030\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__6308\ : InMux
    port map (
            O => \N__29027\,
            I => \N__29021\
        );

    \I__6307\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29021\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__29021\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\
        );

    \I__6305\ : InMux
    port map (
            O => \N__29018\,
            I => \N__29015\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__29015\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29012\,
            I => \N__29009\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__29009\,
            I => \VPP_VDDQ.un1_count_2_1_axb_5\
        );

    \I__6301\ : InMux
    port map (
            O => \N__29006\,
            I => \N__29003\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__29003\,
            I => \N__28999\
        );

    \I__6299\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28996\
        );

    \I__6298\ : Odrv4
    port map (
            O => \N__28999\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__28996\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\
        );

    \I__6296\ : InMux
    port map (
            O => \N__28991\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__6295\ : InMux
    port map (
            O => \N__28988\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__6294\ : InMux
    port map (
            O => \N__28985\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__6293\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28978\
        );

    \I__6292\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28975\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__28978\,
            I => \N__28972\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__28975\,
            I => \N__28969\
        );

    \I__6289\ : Span4Mux_s2_h
    port map (
            O => \N__28972\,
            I => \N__28966\
        );

    \I__6288\ : Span4Mux_s2_h
    port map (
            O => \N__28969\,
            I => \N__28963\
        );

    \I__6287\ : Span4Mux_v
    port map (
            O => \N__28966\,
            I => \N__28960\
        );

    \I__6286\ : Span4Mux_v
    port map (
            O => \N__28963\,
            I => \N__28957\
        );

    \I__6285\ : Odrv4
    port map (
            O => \N__28960\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__6284\ : Odrv4
    port map (
            O => \N__28957\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__6283\ : InMux
    port map (
            O => \N__28952\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__6282\ : CascadeMux
    port map (
            O => \N__28949\,
            I => \N__28945\
        );

    \I__6281\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28940\
        );

    \I__6280\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28940\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__28940\,
            I => \N__28937\
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__28937\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\
        );

    \I__6277\ : InMux
    port map (
            O => \N__28934\,
            I => \bfn_11_12_0_\
        );

    \I__6276\ : InMux
    port map (
            O => \N__28931\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__6275\ : InMux
    port map (
            O => \N__28928\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__6274\ : InMux
    port map (
            O => \N__28925\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__6273\ : InMux
    port map (
            O => \N__28922\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__28919\,
            I => \N__28915\
        );

    \I__6271\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28910\
        );

    \I__6270\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28910\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__28910\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__6268\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28901\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28901\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__28901\,
            I => \VPP_VDDQ.count_2_1_4\
        );

    \I__6265\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28895\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__28895\,
            I => \VPP_VDDQ.count_2_1_5\
        );

    \I__6263\ : CascadeMux
    port map (
            O => \N__28892\,
            I => \VPP_VDDQ.count_2_1_5_cascade_\
        );

    \I__6262\ : CascadeMux
    port map (
            O => \N__28889\,
            I => \N__28886\
        );

    \I__6261\ : InMux
    port map (
            O => \N__28886\,
            I => \N__28880\
        );

    \I__6260\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28880\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__28880\,
            I => \N__28877\
        );

    \I__6258\ : Odrv12
    port map (
            O => \N__28877\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__28874\,
            I => \N__28871\
        );

    \I__6256\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28865\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28865\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__28865\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__6253\ : CascadeMux
    port map (
            O => \N__28862\,
            I => \N__28859\
        );

    \I__6252\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28856\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__6250\ : Span4Mux_v
    port map (
            O => \N__28853\,
            I => \N__28850\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__28850\,
            I => \N__28847\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__28847\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__6247\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__28841\,
            I => \VPP_VDDQ.un1_count_2_1_axb_2\
        );

    \I__6245\ : InMux
    port map (
            O => \N__28838\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__6244\ : InMux
    port map (
            O => \N__28835\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__6243\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28829\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__28829\,
            I => \VPP_VDDQ.un1_count_2_1_axb_4\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__28826\,
            I => \N__28823\
        );

    \I__6240\ : InMux
    port map (
            O => \N__28823\,
            I => \N__28817\
        );

    \I__6239\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28817\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__28817\,
            I => \N__28814\
        );

    \I__6237\ : Odrv4
    port map (
            O => \N__28814\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\
        );

    \I__6236\ : InMux
    port map (
            O => \N__28811\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__28808\,
            I => \VPP_VDDQ.count_2_1_9_cascade_\
        );

    \I__6234\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28802\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__28802\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__6232\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28796\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__28796\,
            I => \N__28792\
        );

    \I__6230\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28789\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__28792\,
            I => \N__28784\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28784\
        );

    \I__6227\ : Span4Mux_h
    port map (
            O => \N__28784\,
            I => \N__28781\
        );

    \I__6226\ : Span4Mux_s0_h
    port map (
            O => \N__28781\,
            I => \N__28778\
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__28778\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__6224\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28772\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__28772\,
            I => \N__28769\
        );

    \I__6222\ : Span4Mux_v
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__6221\ : Span4Mux_v
    port map (
            O => \N__28766\,
            I => \N__28763\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__28763\,
            I => \VPP_VDDQ.un9_clk_100khz_2\
        );

    \I__6219\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28757\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__28757\,
            I => \VPP_VDDQ.un9_clk_100khz_0\
        );

    \I__6217\ : CascadeMux
    port map (
            O => \N__28754\,
            I => \VPP_VDDQ.un9_clk_100khz_1_cascade_\
        );

    \I__6216\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__28748\,
            I => \VPP_VDDQ.un9_clk_100khz_3\
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__28745\,
            I => \N__28742\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28742\,
            I => \N__28739\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__28739\,
            I => \POWERLED.count_clk_0_10\
        );

    \I__6211\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28730\
        );

    \I__6210\ : InMux
    port map (
            O => \N__28735\,
            I => \N__28730\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__28730\,
            I => \N__28727\
        );

    \I__6208\ : Odrv4
    port map (
            O => \N__28727\,
            I => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\
        );

    \I__6207\ : CascadeMux
    port map (
            O => \N__28724\,
            I => \N__28721\
        );

    \I__6206\ : InMux
    port map (
            O => \N__28721\,
            I => \N__28718\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__28718\,
            I => \N__28715\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__28715\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__6203\ : CascadeMux
    port map (
            O => \N__28712\,
            I => \POWERLED.count_clkZ0Z_10_cascade_\
        );

    \I__6202\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28705\
        );

    \I__6201\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28702\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28699\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__28702\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__28699\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__6197\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28690\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__28693\,
            I => \N__28687\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__28690\,
            I => \N__28684\
        );

    \I__6194\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28681\
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__28684\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__28681\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__28676\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_4_cascade_\
        );

    \I__6190\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28669\
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__28672\,
            I => \N__28666\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__28669\,
            I => \N__28663\
        );

    \I__6187\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28660\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__28663\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__28660\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__6184\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28652\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__28652\,
            I => \POWERLED.count_clk_0_0\
        );

    \I__6182\ : CascadeMux
    port map (
            O => \N__28649\,
            I => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__28646\,
            I => \POWERLED.count_clkZ0Z_0_cascade_\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__28643\,
            I => \POWERLED.N_352_cascade_\
        );

    \I__6179\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28637\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__28637\,
            I => \N__28634\
        );

    \I__6177\ : Span4Mux_h
    port map (
            O => \N__28634\,
            I => \N__28629\
        );

    \I__6176\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28626\
        );

    \I__6175\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28623\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__28629\,
            I => \POWERLED.N_394\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__28626\,
            I => \POWERLED.N_394\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__28623\,
            I => \POWERLED.N_394\
        );

    \I__6171\ : InMux
    port map (
            O => \N__28616\,
            I => \N__28610\
        );

    \I__6170\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28610\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__28610\,
            I => \N__28606\
        );

    \I__6168\ : CascadeMux
    port map (
            O => \N__28609\,
            I => \N__28603\
        );

    \I__6167\ : Span4Mux_s3_h
    port map (
            O => \N__28606\,
            I => \N__28600\
        );

    \I__6166\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28597\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__28600\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__28597\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28586\
        );

    \I__6162\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28586\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__28586\,
            I => \N__28582\
        );

    \I__6160\ : CascadeMux
    port map (
            O => \N__28585\,
            I => \N__28579\
        );

    \I__6159\ : Span4Mux_s3_h
    port map (
            O => \N__28582\,
            I => \N__28576\
        );

    \I__6158\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28573\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__28576\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__28573\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__6155\ : CascadeMux
    port map (
            O => \N__28568\,
            I => \N__28565\
        );

    \I__6154\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28562\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__28562\,
            I => \N__28557\
        );

    \I__6152\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28554\
        );

    \I__6151\ : CascadeMux
    port map (
            O => \N__28560\,
            I => \N__28551\
        );

    \I__6150\ : Span4Mux_s2_h
    port map (
            O => \N__28557\,
            I => \N__28548\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__28554\,
            I => \N__28545\
        );

    \I__6148\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28542\
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__28548\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__28545\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__28542\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__6144\ : InMux
    port map (
            O => \N__28535\,
            I => \N__28529\
        );

    \I__6143\ : InMux
    port map (
            O => \N__28534\,
            I => \N__28529\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__28529\,
            I => \N__28525\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__28528\,
            I => \N__28522\
        );

    \I__6140\ : Span4Mux_v
    port map (
            O => \N__28525\,
            I => \N__28519\
        );

    \I__6139\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28516\
        );

    \I__6138\ : Odrv4
    port map (
            O => \N__28519\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__28516\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__6136\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28507\
        );

    \I__6135\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28504\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__28507\,
            I => \N__28500\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__28504\,
            I => \N__28497\
        );

    \I__6132\ : CascadeMux
    port map (
            O => \N__28503\,
            I => \N__28494\
        );

    \I__6131\ : Span4Mux_h
    port map (
            O => \N__28500\,
            I => \N__28491\
        );

    \I__6130\ : Span4Mux_s3_h
    port map (
            O => \N__28497\,
            I => \N__28488\
        );

    \I__6129\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28485\
        );

    \I__6128\ : Odrv4
    port map (
            O => \N__28491\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__28488\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__28485\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__6125\ : CascadeMux
    port map (
            O => \N__28478\,
            I => \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__28475\,
            I => \N__28467\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__28474\,
            I => \N__28463\
        );

    \I__6122\ : InMux
    port map (
            O => \N__28473\,
            I => \N__28457\
        );

    \I__6121\ : InMux
    port map (
            O => \N__28472\,
            I => \N__28453\
        );

    \I__6120\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28450\
        );

    \I__6119\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28439\
        );

    \I__6118\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28439\
        );

    \I__6117\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28439\
        );

    \I__6116\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28436\
        );

    \I__6115\ : CascadeMux
    port map (
            O => \N__28462\,
            I => \N__28433\
        );

    \I__6114\ : CascadeMux
    port map (
            O => \N__28461\,
            I => \N__28430\
        );

    \I__6113\ : InMux
    port map (
            O => \N__28460\,
            I => \N__28425\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__28457\,
            I => \N__28421\
        );

    \I__6111\ : InMux
    port map (
            O => \N__28456\,
            I => \N__28418\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__28453\,
            I => \N__28415\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__28450\,
            I => \N__28412\
        );

    \I__6108\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28409\
        );

    \I__6107\ : InMux
    port map (
            O => \N__28448\,
            I => \N__28404\
        );

    \I__6106\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28404\
        );

    \I__6105\ : InMux
    port map (
            O => \N__28446\,
            I => \N__28401\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__28439\,
            I => \N__28398\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__28436\,
            I => \N__28395\
        );

    \I__6102\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28388\
        );

    \I__6101\ : InMux
    port map (
            O => \N__28430\,
            I => \N__28388\
        );

    \I__6100\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28388\
        );

    \I__6099\ : InMux
    port map (
            O => \N__28428\,
            I => \N__28385\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__28425\,
            I => \N__28382\
        );

    \I__6097\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28379\
        );

    \I__6096\ : Span4Mux_h
    port map (
            O => \N__28421\,
            I => \N__28368\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__28418\,
            I => \N__28368\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__28415\,
            I => \N__28368\
        );

    \I__6093\ : Span4Mux_v
    port map (
            O => \N__28412\,
            I => \N__28368\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__28409\,
            I => \N__28368\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__28404\,
            I => \N__28365\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__28401\,
            I => \N__28360\
        );

    \I__6089\ : Span4Mux_s2_v
    port map (
            O => \N__28398\,
            I => \N__28360\
        );

    \I__6088\ : Span4Mux_v
    port map (
            O => \N__28395\,
            I => \N__28349\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__28388\,
            I => \N__28349\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28349\
        );

    \I__6085\ : Span4Mux_v
    port map (
            O => \N__28382\,
            I => \N__28349\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__28379\,
            I => \N__28349\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__28368\,
            I => \N__28346\
        );

    \I__6082\ : Span4Mux_h
    port map (
            O => \N__28365\,
            I => \N__28341\
        );

    \I__6081\ : Span4Mux_h
    port map (
            O => \N__28360\,
            I => \N__28341\
        );

    \I__6080\ : Span4Mux_v
    port map (
            O => \N__28349\,
            I => \N__28337\
        );

    \I__6079\ : Span4Mux_h
    port map (
            O => \N__28346\,
            I => \N__28332\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__28341\,
            I => \N__28332\
        );

    \I__6077\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28329\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__28337\,
            I => \POWERLED.N_2182_i\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__28332\,
            I => \POWERLED.N_2182_i\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__28329\,
            I => \POWERLED.N_2182_i\
        );

    \I__6073\ : InMux
    port map (
            O => \N__28322\,
            I => \N__28319\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__28319\,
            I => \POWERLED.N_352\
        );

    \I__6071\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28306\
        );

    \I__6070\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28306\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28314\,
            I => \N__28306\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__28313\,
            I => \N__28303\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__28306\,
            I => \N__28300\
        );

    \I__6066\ : InMux
    port map (
            O => \N__28303\,
            I => \N__28297\
        );

    \I__6065\ : Span4Mux_s2_h
    port map (
            O => \N__28300\,
            I => \N__28294\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28291\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__28294\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__6062\ : Odrv4
    port map (
            O => \N__28291\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__6061\ : CascadeMux
    port map (
            O => \N__28286\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_2_2_cascade_\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28274\
        );

    \I__6059\ : InMux
    port map (
            O => \N__28282\,
            I => \N__28274\
        );

    \I__6058\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28274\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__28274\,
            I => \POWERLED.count_clk_RNIZ0Z_9\
        );

    \I__6056\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28265\
        );

    \I__6055\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28265\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__28265\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__6053\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__28259\,
            I => \N__28256\
        );

    \I__6051\ : Span4Mux_v
    port map (
            O => \N__28256\,
            I => \N__28253\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__28253\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_0\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__28250\,
            I => \N__28246\
        );

    \I__6048\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28243\
        );

    \I__6047\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28238\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__28243\,
            I => \N__28235\
        );

    \I__6045\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28232\
        );

    \I__6044\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28229\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__28238\,
            I => \N__28226\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__28235\,
            I => \N__28221\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__28232\,
            I => \N__28221\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__28229\,
            I => \N__28218\
        );

    \I__6039\ : Odrv4
    port map (
            O => \N__28226\,
            I => \POWERLED.func_state_RNI_2Z0Z_1\
        );

    \I__6038\ : Odrv4
    port map (
            O => \N__28221\,
            I => \POWERLED.func_state_RNI_2Z0Z_1\
        );

    \I__6037\ : Odrv12
    port map (
            O => \N__28218\,
            I => \POWERLED.func_state_RNI_2Z0Z_1\
        );

    \I__6036\ : CascadeMux
    port map (
            O => \N__28211\,
            I => \POWERLED.N_289_cascade_\
        );

    \I__6035\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28204\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28201\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28197\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__28201\,
            I => \N__28194\
        );

    \I__6031\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28191\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__28197\,
            I => \N__28188\
        );

    \I__6029\ : Span4Mux_v
    port map (
            O => \N__28194\,
            I => \N__28185\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__28191\,
            I => \POWERLED.func_state_RNIBVNS_2Z0Z_0\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__28188\,
            I => \POWERLED.func_state_RNIBVNS_2Z0Z_0\
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__28185\,
            I => \POWERLED.func_state_RNIBVNS_2Z0Z_0\
        );

    \I__6025\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28174\
        );

    \I__6024\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28171\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__28174\,
            I => \N__28167\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__28171\,
            I => \N__28164\
        );

    \I__6021\ : InMux
    port map (
            O => \N__28170\,
            I => \N__28161\
        );

    \I__6020\ : Span4Mux_v
    port map (
            O => \N__28167\,
            I => \N__28153\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__28164\,
            I => \N__28148\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__28161\,
            I => \N__28148\
        );

    \I__6017\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28145\
        );

    \I__6016\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28140\
        );

    \I__6015\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28140\
        );

    \I__6014\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28135\
        );

    \I__6013\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28135\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__28153\,
            I => \POWERLED.count_off_RNIG5N6N1Z0Z_11\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__28148\,
            I => \POWERLED.count_off_RNIG5N6N1Z0Z_11\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__28145\,
            I => \POWERLED.count_off_RNIG5N6N1Z0Z_11\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__28140\,
            I => \POWERLED.count_off_RNIG5N6N1Z0Z_11\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__28135\,
            I => \POWERLED.count_off_RNIG5N6N1Z0Z_11\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__28124\,
            I => \N__28121\
        );

    \I__6006\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28117\
        );

    \I__6005\ : InMux
    port map (
            O => \N__28120\,
            I => \N__28114\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__28117\,
            I => \N__28111\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__28114\,
            I => \N__28108\
        );

    \I__6002\ : Span4Mux_h
    port map (
            O => \N__28111\,
            I => \N__28105\
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__28108\,
            I => \POWERLED.func_state_RNI_5Z0Z_1\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__28105\,
            I => \POWERLED.func_state_RNI_5Z0Z_1\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__28100\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_2_tz_0_cascade_\
        );

    \I__5998\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__5996\ : Odrv12
    port map (
            O => \N__28091\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_2\
        );

    \I__5995\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28084\
        );

    \I__5994\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28081\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__28084\,
            I => \N__28076\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__28081\,
            I => \N__28076\
        );

    \I__5991\ : Odrv4
    port map (
            O => \N__28076\,
            I => \POWERLED.func_state_RNI_2Z0Z_0\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__28073\,
            I => \N__28069\
        );

    \I__5989\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28060\
        );

    \I__5988\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28060\
        );

    \I__5987\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28057\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__28067\,
            I => \N__28049\
        );

    \I__5985\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28045\
        );

    \I__5984\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28042\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__28060\,
            I => \N__28038\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28035\
        );

    \I__5981\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28032\
        );

    \I__5980\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28024\
        );

    \I__5979\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28021\
        );

    \I__5978\ : InMux
    port map (
            O => \N__28053\,
            I => \N__28018\
        );

    \I__5977\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28015\
        );

    \I__5976\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28010\
        );

    \I__5975\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28010\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__28045\,
            I => \N__28005\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__28042\,
            I => \N__28005\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__28041\,
            I => \N__28002\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__28038\,
            I => \N__27996\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__28035\,
            I => \N__27996\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__28032\,
            I => \N__27993\
        );

    \I__5968\ : InMux
    port map (
            O => \N__28031\,
            I => \N__27990\
        );

    \I__5967\ : InMux
    port map (
            O => \N__28030\,
            I => \N__27983\
        );

    \I__5966\ : InMux
    port map (
            O => \N__28029\,
            I => \N__27983\
        );

    \I__5965\ : InMux
    port map (
            O => \N__28028\,
            I => \N__27983\
        );

    \I__5964\ : InMux
    port map (
            O => \N__28027\,
            I => \N__27980\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__28024\,
            I => \N__27976\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__28021\,
            I => \N__27973\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__28018\,
            I => \N__27970\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__28015\,
            I => \N__27965\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__28010\,
            I => \N__27965\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__28005\,
            I => \N__27962\
        );

    \I__5957\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27957\
        );

    \I__5956\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27957\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__27996\,
            I => \N__27952\
        );

    \I__5954\ : Span4Mux_v
    port map (
            O => \N__27993\,
            I => \N__27952\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__27990\,
            I => \N__27949\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__27983\,
            I => \N__27946\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__27980\,
            I => \N__27943\
        );

    \I__5950\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27940\
        );

    \I__5949\ : Span4Mux_v
    port map (
            O => \N__27976\,
            I => \N__27931\
        );

    \I__5948\ : Span4Mux_s3_v
    port map (
            O => \N__27973\,
            I => \N__27931\
        );

    \I__5947\ : Span4Mux_s3_v
    port map (
            O => \N__27970\,
            I => \N__27931\
        );

    \I__5946\ : Span4Mux_v
    port map (
            O => \N__27965\,
            I => \N__27931\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__27962\,
            I => \N__27926\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__27957\,
            I => \N__27926\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__27952\,
            I => \N__27919\
        );

    \I__5942\ : Span4Mux_h
    port map (
            O => \N__27949\,
            I => \N__27919\
        );

    \I__5941\ : Span4Mux_s3_v
    port map (
            O => \N__27946\,
            I => \N__27919\
        );

    \I__5940\ : Span12Mux_s3_v
    port map (
            O => \N__27943\,
            I => \N__27914\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27914\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__27931\,
            I => \N__27909\
        );

    \I__5937\ : Span4Mux_v
    port map (
            O => \N__27926\,
            I => \N__27909\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__27919\,
            I => gpio_fpga_soc_4
        );

    \I__5935\ : Odrv12
    port map (
            O => \N__27914\,
            I => gpio_fpga_soc_4
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__27909\,
            I => gpio_fpga_soc_4
        );

    \I__5933\ : InMux
    port map (
            O => \N__27902\,
            I => \N__27899\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__5931\ : Span4Mux_h
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__5930\ : Odrv4
    port map (
            O => \N__27893\,
            I => \POWERLED.un1_func_state25_6_0_o_N_304_N\
        );

    \I__5929\ : InMux
    port map (
            O => \N__27890\,
            I => \N__27886\
        );

    \I__5928\ : CascadeMux
    port map (
            O => \N__27889\,
            I => \N__27877\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27873\
        );

    \I__5926\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27870\
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__27884\,
            I => \N__27867\
        );

    \I__5924\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27860\
        );

    \I__5923\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27860\
        );

    \I__5922\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27860\
        );

    \I__5921\ : CascadeMux
    port map (
            O => \N__27880\,
            I => \N__27856\
        );

    \I__5920\ : InMux
    port map (
            O => \N__27877\,
            I => \N__27853\
        );

    \I__5919\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27850\
        );

    \I__5918\ : Sp12to4
    port map (
            O => \N__27873\,
            I => \N__27845\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__27870\,
            I => \N__27845\
        );

    \I__5916\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27842\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__27860\,
            I => \N__27839\
        );

    \I__5914\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27836\
        );

    \I__5913\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27832\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__27853\,
            I => \N__27827\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__27850\,
            I => \N__27827\
        );

    \I__5910\ : Span12Mux_s11_v
    port map (
            O => \N__27845\,
            I => \N__27824\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__27842\,
            I => \N__27819\
        );

    \I__5908\ : Span4Mux_s3_h
    port map (
            O => \N__27839\,
            I => \N__27819\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__27836\,
            I => \N__27816\
        );

    \I__5906\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27813\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__27832\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__27827\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5903\ : Odrv12
    port map (
            O => \N__27824\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__27819\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5901\ : Odrv12
    port map (
            O => \N__27816\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__27813\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5899\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27791\
        );

    \I__5898\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27788\
        );

    \I__5897\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27783\
        );

    \I__5896\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27783\
        );

    \I__5895\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27780\
        );

    \I__5894\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27772\
        );

    \I__5893\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27769\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__27791\,
            I => \N__27764\
        );

    \I__5891\ : InMux
    port map (
            O => \N__27788\,
            I => \N__27761\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__27783\,
            I => \N__27756\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__27780\,
            I => \N__27756\
        );

    \I__5888\ : InMux
    port map (
            O => \N__27779\,
            I => \N__27749\
        );

    \I__5887\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27749\
        );

    \I__5886\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27749\
        );

    \I__5885\ : InMux
    port map (
            O => \N__27776\,
            I => \N__27744\
        );

    \I__5884\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27744\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__27772\,
            I => \N__27741\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__27769\,
            I => \N__27729\
        );

    \I__5881\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27726\
        );

    \I__5880\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27723\
        );

    \I__5879\ : Span4Mux_v
    port map (
            O => \N__27764\,
            I => \N__27720\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__27761\,
            I => \N__27717\
        );

    \I__5877\ : Span4Mux_v
    port map (
            O => \N__27756\,
            I => \N__27714\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__27749\,
            I => \N__27709\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__27744\,
            I => \N__27709\
        );

    \I__5874\ : Span4Mux_v
    port map (
            O => \N__27741\,
            I => \N__27706\
        );

    \I__5873\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27703\
        );

    \I__5872\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27694\
        );

    \I__5871\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27694\
        );

    \I__5870\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27694\
        );

    \I__5869\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27694\
        );

    \I__5868\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27685\
        );

    \I__5867\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27685\
        );

    \I__5866\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27685\
        );

    \I__5865\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27685\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__27729\,
            I => \N__27678\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27678\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__27723\,
            I => \N__27678\
        );

    \I__5861\ : Odrv4
    port map (
            O => \N__27720\,
            I => \POWERLED.func_state\
        );

    \I__5860\ : Odrv12
    port map (
            O => \N__27717\,
            I => \POWERLED.func_state\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__27714\,
            I => \POWERLED.func_state\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__27709\,
            I => \POWERLED.func_state\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__27706\,
            I => \POWERLED.func_state\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__27703\,
            I => \POWERLED.func_state\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__27694\,
            I => \POWERLED.func_state\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__27685\,
            I => \POWERLED.func_state\
        );

    \I__5853\ : Odrv4
    port map (
            O => \N__27678\,
            I => \POWERLED.func_state\
        );

    \I__5852\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27656\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__27656\,
            I => \N__27653\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__27653\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_2_0\
        );

    \I__5849\ : CascadeMux
    port map (
            O => \N__27650\,
            I => \N__27647\
        );

    \I__5848\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27644\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__27644\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_3_0\
        );

    \I__5846\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27638\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__27638\,
            I => \POWERLED.count_off_1_2\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__27635\,
            I => \POWERLED.count_off_1_2_cascade_\
        );

    \I__5843\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27626\
        );

    \I__5842\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27626\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__27626\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__5840\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27620\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__27620\,
            I => \POWERLED.count_off_1_7\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__27617\,
            I => \POWERLED.count_off_1_7_cascade_\
        );

    \I__5837\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__27611\,
            I => \POWERLED.un34_clk_100khz_3\
        );

    \I__5835\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27602\
        );

    \I__5834\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27602\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__27602\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__5832\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27596\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__27596\,
            I => \N__27593\
        );

    \I__5830\ : Span4Mux_v
    port map (
            O => \N__27593\,
            I => \N__27590\
        );

    \I__5829\ : Odrv4
    port map (
            O => \N__27590\,
            I => \POWERLED.count_off_1_11\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__27587\,
            I => \POWERLED.count_off_1_11_cascade_\
        );

    \I__5827\ : CascadeMux
    port map (
            O => \N__27584\,
            I => \N__27581\
        );

    \I__5826\ : InMux
    port map (
            O => \N__27581\,
            I => \N__27578\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__27578\,
            I => \N__27575\
        );

    \I__5824\ : Span4Mux_v
    port map (
            O => \N__27575\,
            I => \N__27571\
        );

    \I__5823\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27568\
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__27571\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__27568\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__5820\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27560\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__27560\,
            I => \POWERLED.count_off_0_15\
        );

    \I__5818\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27554\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__27554\,
            I => \POWERLED.count_off_0_8\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__27551\,
            I => \POWERLED.un34_clk_100khz_0_cascade_\
        );

    \I__5815\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__5813\ : Odrv12
    port map (
            O => \N__27542\,
            I => \POWERLED.un34_clk_100khz_12\
        );

    \I__5812\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__27536\,
            I => \POWERLED.un34_clk_100khz_1\
        );

    \I__5810\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27530\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__27530\,
            I => \POWERLED.count_off_1_6\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__27527\,
            I => \POWERLED.count_off_1_6_cascade_\
        );

    \I__5807\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27520\
        );

    \I__5806\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27517\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__27517\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__5803\ : Odrv4
    port map (
            O => \N__27514\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__5802\ : InMux
    port map (
            O => \N__27509\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__5801\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27502\
        );

    \I__5800\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27499\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__27502\,
            I => \N__27496\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__27499\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__27496\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__5796\ : InMux
    port map (
            O => \N__27491\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27484\
        );

    \I__5794\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27481\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__27484\,
            I => \N__27478\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__27481\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__27478\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__5790\ : InMux
    port map (
            O => \N__27473\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__5789\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27465\
        );

    \I__5788\ : InMux
    port map (
            O => \N__27469\,
            I => \N__27462\
        );

    \I__5787\ : InMux
    port map (
            O => \N__27468\,
            I => \N__27457\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__27465\,
            I => \N__27454\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__27462\,
            I => \N__27450\
        );

    \I__5784\ : InMux
    port map (
            O => \N__27461\,
            I => \N__27446\
        );

    \I__5783\ : IoInMux
    port map (
            O => \N__27460\,
            I => \N__27442\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__27457\,
            I => \N__27439\
        );

    \I__5781\ : Span4Mux_s1_h
    port map (
            O => \N__27454\,
            I => \N__27436\
        );

    \I__5780\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27433\
        );

    \I__5779\ : Span4Mux_v
    port map (
            O => \N__27450\,
            I => \N__27430\
        );

    \I__5778\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27427\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27424\
        );

    \I__5776\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27421\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27418\
        );

    \I__5774\ : Span4Mux_v
    port map (
            O => \N__27439\,
            I => \N__27415\
        );

    \I__5773\ : Span4Mux_h
    port map (
            O => \N__27436\,
            I => \N__27410\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__27433\,
            I => \N__27410\
        );

    \I__5771\ : Span4Mux_h
    port map (
            O => \N__27430\,
            I => \N__27405\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__27427\,
            I => \N__27405\
        );

    \I__5769\ : Span4Mux_v
    port map (
            O => \N__27424\,
            I => \N__27400\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__27421\,
            I => \N__27400\
        );

    \I__5767\ : Span4Mux_s3_h
    port map (
            O => \N__27418\,
            I => \N__27397\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__27415\,
            I => \N__27392\
        );

    \I__5765\ : Span4Mux_v
    port map (
            O => \N__27410\,
            I => \N__27392\
        );

    \I__5764\ : Span4Mux_v
    port map (
            O => \N__27405\,
            I => \N__27387\
        );

    \I__5763\ : Span4Mux_h
    port map (
            O => \N__27400\,
            I => \N__27387\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__27397\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__27392\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__27387\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5759\ : InMux
    port map (
            O => \N__27380\,
            I => \bfn_9_15_0_\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__27377\,
            I => \N__27374\
        );

    \I__5757\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27370\
        );

    \I__5756\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27367\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__27370\,
            I => \N__27364\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__27367\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__5753\ : Odrv12
    port map (
            O => \N__27364\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__5751\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__27353\,
            I => \POWERLED.count_off_0_5\
        );

    \I__5749\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27346\
        );

    \I__5748\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27343\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__27346\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__27343\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__5745\ : InMux
    port map (
            O => \N__27338\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__5744\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27331\
        );

    \I__5743\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27328\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__27331\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__27328\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__5740\ : InMux
    port map (
            O => \N__27323\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__5739\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27316\
        );

    \I__5738\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27313\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__27316\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__27313\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__5735\ : InMux
    port map (
            O => \N__27308\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__5734\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27301\
        );

    \I__5733\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27298\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__27301\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__27298\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__5730\ : InMux
    port map (
            O => \N__27293\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__27290\,
            I => \N__27286\
        );

    \I__5728\ : InMux
    port map (
            O => \N__27289\,
            I => \N__27283\
        );

    \I__5727\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27280\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__27283\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__27280\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__5724\ : InMux
    port map (
            O => \N__27275\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__5723\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27268\
        );

    \I__5722\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27265\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__27268\,
            I => \N__27262\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__27265\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__27262\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__5718\ : InMux
    port map (
            O => \N__27257\,
            I => \bfn_9_14_0_\
        );

    \I__5717\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27250\
        );

    \I__5716\ : InMux
    port map (
            O => \N__27253\,
            I => \N__27247\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__27250\,
            I => \N__27244\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__27247\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__5713\ : Odrv4
    port map (
            O => \N__27244\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__5712\ : InMux
    port map (
            O => \N__27239\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__5710\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27229\
        );

    \I__5709\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27226\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27223\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__27226\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__5706\ : Odrv4
    port map (
            O => \N__27223\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__5705\ : InMux
    port map (
            O => \N__27218\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__5704\ : CascadeMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__5703\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27208\
        );

    \I__5702\ : InMux
    port map (
            O => \N__27211\,
            I => \N__27205\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__27208\,
            I => \N__27202\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__27205\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__5699\ : Odrv4
    port map (
            O => \N__27202\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__5698\ : InMux
    port map (
            O => \N__27197\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__27194\,
            I => \N__27191\
        );

    \I__5696\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27188\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__27188\,
            I => \N__27185\
        );

    \I__5694\ : Odrv12
    port map (
            O => \N__27185\,
            I => \POWERLED.dutycycle_RNIZ0Z_1\
        );

    \I__5693\ : InMux
    port map (
            O => \N__27182\,
            I => \N__27179\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__27179\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__5691\ : CascadeMux
    port map (
            O => \N__27176\,
            I => \VPP_VDDQ.un6_count_8_cascade_\
        );

    \I__5690\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27170\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__27170\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__5688\ : InMux
    port map (
            O => \N__27167\,
            I => \N__27164\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__27164\,
            I => \VPP_VDDQ.un6_count_9\
        );

    \I__5686\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27157\
        );

    \I__5685\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27154\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__27157\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__27154\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__5682\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27145\
        );

    \I__5681\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27142\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__27145\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__27142\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__5678\ : InMux
    port map (
            O => \N__27137\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__5677\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27130\
        );

    \I__5676\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27127\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__27130\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__27127\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__5673\ : InMux
    port map (
            O => \N__27122\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__5672\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__27116\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_0\
        );

    \I__5670\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__27110\,
            I => \POWERLED.un1_dutycycle_172_m3\
        );

    \I__5668\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27099\
        );

    \I__5667\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27094\
        );

    \I__5666\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27089\
        );

    \I__5665\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27086\
        );

    \I__5664\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27081\
        );

    \I__5663\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27081\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27099\,
            I => \N__27078\
        );

    \I__5661\ : CascadeMux
    port map (
            O => \N__27098\,
            I => \N__27074\
        );

    \I__5660\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27071\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__27094\,
            I => \N__27068\
        );

    \I__5658\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27065\
        );

    \I__5657\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27062\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__27089\,
            I => \N__27055\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__27086\,
            I => \N__27055\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__27081\,
            I => \N__27055\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__27078\,
            I => \N__27049\
        );

    \I__5652\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27046\
        );

    \I__5651\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27043\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__27071\,
            I => \N__27039\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__27068\,
            I => \N__27030\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__27065\,
            I => \N__27030\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__27062\,
            I => \N__27030\
        );

    \I__5646\ : Span4Mux_v
    port map (
            O => \N__27055\,
            I => \N__27030\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__27054\,
            I => \N__27026\
        );

    \I__5644\ : CascadeMux
    port map (
            O => \N__27053\,
            I => \N__27014\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__27052\,
            I => \N__27010\
        );

    \I__5642\ : Span4Mux_v
    port map (
            O => \N__27049\,
            I => \N__27005\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__27046\,
            I => \N__27005\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__27043\,
            I => \N__27002\
        );

    \I__5639\ : InMux
    port map (
            O => \N__27042\,
            I => \N__26999\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__27039\,
            I => \N__26994\
        );

    \I__5637\ : Span4Mux_v
    port map (
            O => \N__27030\,
            I => \N__26994\
        );

    \I__5636\ : InMux
    port map (
            O => \N__27029\,
            I => \N__26985\
        );

    \I__5635\ : InMux
    port map (
            O => \N__27026\,
            I => \N__26985\
        );

    \I__5634\ : InMux
    port map (
            O => \N__27025\,
            I => \N__26985\
        );

    \I__5633\ : InMux
    port map (
            O => \N__27024\,
            I => \N__26985\
        );

    \I__5632\ : InMux
    port map (
            O => \N__27023\,
            I => \N__26976\
        );

    \I__5631\ : InMux
    port map (
            O => \N__27022\,
            I => \N__26976\
        );

    \I__5630\ : InMux
    port map (
            O => \N__27021\,
            I => \N__26976\
        );

    \I__5629\ : InMux
    port map (
            O => \N__27020\,
            I => \N__26976\
        );

    \I__5628\ : InMux
    port map (
            O => \N__27019\,
            I => \N__26963\
        );

    \I__5627\ : InMux
    port map (
            O => \N__27018\,
            I => \N__26963\
        );

    \I__5626\ : InMux
    port map (
            O => \N__27017\,
            I => \N__26963\
        );

    \I__5625\ : InMux
    port map (
            O => \N__27014\,
            I => \N__26963\
        );

    \I__5624\ : InMux
    port map (
            O => \N__27013\,
            I => \N__26963\
        );

    \I__5623\ : InMux
    port map (
            O => \N__27010\,
            I => \N__26963\
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__27005\,
            I => \POWERLED.N_2200_i\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__27002\,
            I => \POWERLED.N_2200_i\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__26999\,
            I => \POWERLED.N_2200_i\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__26994\,
            I => \POWERLED.N_2200_i\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__26985\,
            I => \POWERLED.N_2200_i\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__26976\,
            I => \POWERLED.N_2200_i\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__26963\,
            I => \POWERLED.N_2200_i\
        );

    \I__5615\ : InMux
    port map (
            O => \N__26948\,
            I => \N__26945\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__26945\,
            I => \POWERLED.un1_dutycycle_96_0_a3_1\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__26942\,
            I => \N__26934\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \N__26929\
        );

    \I__5611\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26924\
        );

    \I__5610\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26924\
        );

    \I__5609\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26918\
        );

    \I__5608\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26913\
        );

    \I__5607\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26913\
        );

    \I__5606\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26910\
        );

    \I__5605\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26907\
        );

    \I__5604\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26904\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__26924\,
            I => \N__26901\
        );

    \I__5602\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26894\
        );

    \I__5601\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26894\
        );

    \I__5600\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26894\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__26918\,
            I => \N__26891\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__26913\,
            I => \N__26888\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__26910\,
            I => \N__26885\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26879\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26879\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__26901\,
            I => \N__26870\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__26894\,
            I => \N__26870\
        );

    \I__5592\ : Span4Mux_v
    port map (
            O => \N__26891\,
            I => \N__26870\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__26888\,
            I => \N__26870\
        );

    \I__5590\ : Span4Mux_h
    port map (
            O => \N__26885\,
            I => \N__26867\
        );

    \I__5589\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26864\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__26879\,
            I => \N__26859\
        );

    \I__5587\ : Span4Mux_v
    port map (
            O => \N__26870\,
            I => \N__26859\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__26867\,
            I => \POWERLED.dutycycle\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__26864\,
            I => \POWERLED.dutycycle\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__26859\,
            I => \POWERLED.dutycycle\
        );

    \I__5583\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26848\
        );

    \I__5582\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26845\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__26848\,
            I => \POWERLED.N_327\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__26845\,
            I => \POWERLED.N_327\
        );

    \I__5579\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26837\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__26837\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_0\
        );

    \I__5577\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26828\
        );

    \I__5576\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26823\
        );

    \I__5575\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26823\
        );

    \I__5574\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26820\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__26828\,
            I => \N__26817\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__26823\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_5\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__26820\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_5\
        );

    \I__5570\ : Odrv4
    port map (
            O => \N__26817\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_5\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__26810\,
            I => \POWERLED.un1_dutycycle_53_axb_3_1_0_cascade_\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__26807\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_1_cascade_\
        );

    \I__5567\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26801\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26798\
        );

    \I__5565\ : Odrv12
    port map (
            O => \N__26798\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_2\
        );

    \I__5564\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26792\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__26792\,
            I => \N__26789\
        );

    \I__5562\ : Span4Mux_v
    port map (
            O => \N__26789\,
            I => \N__26785\
        );

    \I__5561\ : InMux
    port map (
            O => \N__26788\,
            I => \N__26782\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__26785\,
            I => \POWERLED.N_342\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__26782\,
            I => \POWERLED.N_342\
        );

    \I__5558\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__5556\ : Span4Mux_v
    port map (
            O => \N__26771\,
            I => \N__26766\
        );

    \I__5555\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26763\
        );

    \I__5554\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26760\
        );

    \I__5553\ : Span4Mux_h
    port map (
            O => \N__26766\,
            I => \N__26755\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__26763\,
            I => \N__26755\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__26760\,
            I => \POWERLED.N_155\
        );

    \I__5550\ : Odrv4
    port map (
            O => \N__26755\,
            I => \POWERLED.N_155\
        );

    \I__5549\ : CascadeMux
    port map (
            O => \N__26750\,
            I => \N__26746\
        );

    \I__5548\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26743\
        );

    \I__5547\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26740\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__26743\,
            I => \N__26736\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__26740\,
            I => \N__26733\
        );

    \I__5544\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26730\
        );

    \I__5543\ : Span4Mux_s3_h
    port map (
            O => \N__26736\,
            I => \N__26727\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__26733\,
            I => \N__26724\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__26730\,
            I => \N__26721\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__26727\,
            I => \N__26718\
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__26724\,
            I => \POWERLED.N_336\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__26721\,
            I => \POWERLED.N_336\
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__26718\,
            I => \POWERLED.N_336\
        );

    \I__5536\ : InMux
    port map (
            O => \N__26711\,
            I => \N__26708\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__26708\,
            I => \N__26704\
        );

    \I__5534\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26701\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__26704\,
            I => \POWERLED.dutycycle_RNI_9Z0Z_0\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__26701\,
            I => \POWERLED.dutycycle_RNI_9Z0Z_0\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__26696\,
            I => \N__26689\
        );

    \I__5530\ : InMux
    port map (
            O => \N__26695\,
            I => \N__26686\
        );

    \I__5529\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26683\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__26693\,
            I => \N__26678\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__26692\,
            I => \N__26672\
        );

    \I__5526\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26669\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__26686\,
            I => \N__26666\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__26683\,
            I => \N__26663\
        );

    \I__5523\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26660\
        );

    \I__5522\ : InMux
    port map (
            O => \N__26681\,
            I => \N__26655\
        );

    \I__5521\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26655\
        );

    \I__5520\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26652\
        );

    \I__5519\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26647\
        );

    \I__5518\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26647\
        );

    \I__5517\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26644\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__26669\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5515\ : Odrv12
    port map (
            O => \N__26666\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5514\ : Odrv12
    port map (
            O => \N__26663\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__26660\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__26655\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__26652\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__26647\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__26644\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__26627\,
            I => \N__26623\
        );

    \I__5507\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26619\
        );

    \I__5506\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26614\
        );

    \I__5505\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26614\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__26619\,
            I => \N__26608\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__26614\,
            I => \N__26608\
        );

    \I__5502\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26603\
        );

    \I__5501\ : Span4Mux_v
    port map (
            O => \N__26608\,
            I => \N__26596\
        );

    \I__5500\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26591\
        );

    \I__5499\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26591\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__26603\,
            I => \N__26588\
        );

    \I__5497\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26579\
        );

    \I__5496\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26579\
        );

    \I__5495\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26579\
        );

    \I__5494\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26579\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__26596\,
            I => \N__26569\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26569\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__26588\,
            I => \N__26559\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__26579\,
            I => \N__26559\
        );

    \I__5489\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26556\
        );

    \I__5488\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26551\
        );

    \I__5487\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26548\
        );

    \I__5486\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26543\
        );

    \I__5485\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26543\
        );

    \I__5484\ : Span4Mux_h
    port map (
            O => \N__26569\,
            I => \N__26540\
        );

    \I__5483\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26529\
        );

    \I__5482\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26529\
        );

    \I__5481\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26529\
        );

    \I__5480\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26529\
        );

    \I__5479\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26529\
        );

    \I__5478\ : Sp12to4
    port map (
            O => \N__26559\,
            I => \N__26524\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__26556\,
            I => \N__26524\
        );

    \I__5476\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26519\
        );

    \I__5475\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26519\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__26551\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__26548\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__26543\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__26540\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__26529\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__5469\ : Odrv12
    port map (
            O => \N__26524\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__26519\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__5467\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26498\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__26495\,
            I => \POWERLED.un1_i3_mux\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__26492\,
            I => \N__26484\
        );

    \I__5462\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26479\
        );

    \I__5461\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26476\
        );

    \I__5460\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26472\
        );

    \I__5459\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26463\
        );

    \I__5458\ : InMux
    port map (
            O => \N__26487\,
            I => \N__26463\
        );

    \I__5457\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26463\
        );

    \I__5456\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26463\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__26482\,
            I => \N__26459\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__26479\,
            I => \N__26452\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__26476\,
            I => \N__26449\
        );

    \I__5452\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26446\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__26472\,
            I => \N__26441\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__26463\,
            I => \N__26441\
        );

    \I__5449\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26438\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26435\
        );

    \I__5447\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26426\
        );

    \I__5446\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26426\
        );

    \I__5445\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26426\
        );

    \I__5444\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26426\
        );

    \I__5443\ : Span4Mux_v
    port map (
            O => \N__26452\,
            I => \N__26417\
        );

    \I__5442\ : Span4Mux_h
    port map (
            O => \N__26449\,
            I => \N__26417\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__26446\,
            I => \N__26417\
        );

    \I__5440\ : Span4Mux_v
    port map (
            O => \N__26441\,
            I => \N__26417\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26412\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__26435\,
            I => \N__26412\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__26426\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__26417\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__5435\ : Odrv4
    port map (
            O => \N__26412\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__5433\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26398\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__26401\,
            I => \N__26384\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__26398\,
            I => \N__26377\
        );

    \I__5430\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26372\
        );

    \I__5429\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26372\
        );

    \I__5428\ : InMux
    port map (
            O => \N__26395\,
            I => \N__26367\
        );

    \I__5427\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26367\
        );

    \I__5426\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26364\
        );

    \I__5425\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26359\
        );

    \I__5424\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26359\
        );

    \I__5423\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26354\
        );

    \I__5422\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26347\
        );

    \I__5421\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26347\
        );

    \I__5420\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26347\
        );

    \I__5419\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26344\
        );

    \I__5418\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26335\
        );

    \I__5417\ : InMux
    port map (
            O => \N__26382\,
            I => \N__26335\
        );

    \I__5416\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26335\
        );

    \I__5415\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26335\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__26377\,
            I => \N__26332\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26325\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__26367\,
            I => \N__26325\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__26364\,
            I => \N__26325\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26322\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__26358\,
            I => \N__26319\
        );

    \I__5408\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26316\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__26354\,
            I => \N__26311\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__26347\,
            I => \N__26311\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__26344\,
            I => \N__26300\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__26335\,
            I => \N__26300\
        );

    \I__5403\ : Span4Mux_s1_v
    port map (
            O => \N__26332\,
            I => \N__26300\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__26325\,
            I => \N__26300\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__26322\,
            I => \N__26300\
        );

    \I__5400\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26297\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__26316\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__26311\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5397\ : Odrv4
    port map (
            O => \N__26300\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__26297\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__26288\,
            I => \N__26283\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__26287\,
            I => \N__26279\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__26286\,
            I => \N__26275\
        );

    \I__5392\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26270\
        );

    \I__5391\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26267\
        );

    \I__5390\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26260\
        );

    \I__5389\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26260\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26253\
        );

    \I__5387\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26253\
        );

    \I__5386\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26253\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26248\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__26267\,
            I => \N__26248\
        );

    \I__5383\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26245\
        );

    \I__5382\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26242\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__26260\,
            I => \N__26237\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__26253\,
            I => \N__26234\
        );

    \I__5379\ : Span4Mux_h
    port map (
            O => \N__26248\,
            I => \N__26229\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__26245\,
            I => \N__26229\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__26242\,
            I => \N__26226\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__26241\,
            I => \N__26223\
        );

    \I__5375\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26220\
        );

    \I__5374\ : Span4Mux_h
    port map (
            O => \N__26237\,
            I => \N__26215\
        );

    \I__5373\ : Span4Mux_h
    port map (
            O => \N__26234\,
            I => \N__26215\
        );

    \I__5372\ : Span4Mux_h
    port map (
            O => \N__26229\,
            I => \N__26210\
        );

    \I__5371\ : Span4Mux_v
    port map (
            O => \N__26226\,
            I => \N__26210\
        );

    \I__5370\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26207\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__26220\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__26215\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__26210\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26207\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__26198\,
            I => \N__26195\
        );

    \I__5364\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26185\
        );

    \I__5363\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26185\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__26193\,
            I => \N__26181\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__26192\,
            I => \N__26178\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__26191\,
            I => \N__26175\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__26190\,
            I => \N__26172\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__26185\,
            I => \N__26167\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__26184\,
            I => \N__26162\
        );

    \I__5356\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26157\
        );

    \I__5355\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26157\
        );

    \I__5354\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26154\
        );

    \I__5353\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26150\
        );

    \I__5352\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26145\
        );

    \I__5351\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26145\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__26167\,
            I => \N__26142\
        );

    \I__5349\ : InMux
    port map (
            O => \N__26166\,
            I => \N__26139\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26136\
        );

    \I__5347\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26133\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26128\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__26154\,
            I => \N__26128\
        );

    \I__5344\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26125\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__26150\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__26145\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5341\ : Odrv4
    port map (
            O => \N__26142\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__26139\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__26136\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__26133\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__26128\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__26125\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5335\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__26105\,
            I => \N__26102\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__26102\,
            I => \N__26099\
        );

    \I__5332\ : Span4Mux_v
    port map (
            O => \N__26099\,
            I => \N__26094\
        );

    \I__5331\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26091\
        );

    \I__5330\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26088\
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__26094\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__26091\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__26088\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__5326\ : CascadeMux
    port map (
            O => \N__26081\,
            I => \N__26078\
        );

    \I__5325\ : InMux
    port map (
            O => \N__26078\,
            I => \N__26075\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__26075\,
            I => \N__26072\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__26072\,
            I => \N__26069\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__26069\,
            I => \N__26066\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__26066\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__26063\,
            I => \N__26060\
        );

    \I__5319\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26057\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__26057\,
            I => \N__26054\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__26054\,
            I => \N__26050\
        );

    \I__5316\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26047\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__26050\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_0\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__26047\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_0\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__26042\,
            I => \POWERLED.un1_dutycycle_172_m4_bm_rn_0_cascade_\
        );

    \I__5312\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26036\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__26036\,
            I => \POWERLED.dutycycle_RNIMUFP1Z0Z_2\
        );

    \I__5310\ : InMux
    port map (
            O => \N__26033\,
            I => \N__26023\
        );

    \I__5309\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26020\
        );

    \I__5308\ : InMux
    port map (
            O => \N__26031\,
            I => \N__26017\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__26030\,
            I => \N__26013\
        );

    \I__5306\ : CascadeMux
    port map (
            O => \N__26029\,
            I => \N__26010\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__26028\,
            I => \N__26007\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__26027\,
            I => \N__26004\
        );

    \I__5303\ : InMux
    port map (
            O => \N__26026\,
            I => \N__25997\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__26023\,
            I => \N__25992\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__26020\,
            I => \N__25992\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__25989\
        );

    \I__5299\ : InMux
    port map (
            O => \N__26016\,
            I => \N__25986\
        );

    \I__5298\ : InMux
    port map (
            O => \N__26013\,
            I => \N__25973\
        );

    \I__5297\ : InMux
    port map (
            O => \N__26010\,
            I => \N__25973\
        );

    \I__5296\ : InMux
    port map (
            O => \N__26007\,
            I => \N__25973\
        );

    \I__5295\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25973\
        );

    \I__5294\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25973\
        );

    \I__5293\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25973\
        );

    \I__5292\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25970\
        );

    \I__5291\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25967\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25964\
        );

    \I__5289\ : Span4Mux_s3_v
    port map (
            O => \N__25992\,
            I => \N__25961\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__25989\,
            I => \N__25956\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__25986\,
            I => \N__25956\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__25973\,
            I => \N__25953\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__25970\,
            I => \N__25950\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__25967\,
            I => \N__25947\
        );

    \I__5283\ : Span4Mux_s3_h
    port map (
            O => \N__25964\,
            I => \N__25944\
        );

    \I__5282\ : Span4Mux_h
    port map (
            O => \N__25961\,
            I => \N__25941\
        );

    \I__5281\ : Span4Mux_h
    port map (
            O => \N__25956\,
            I => \N__25938\
        );

    \I__5280\ : Span4Mux_h
    port map (
            O => \N__25953\,
            I => \N__25933\
        );

    \I__5279\ : Span4Mux_h
    port map (
            O => \N__25950\,
            I => \N__25933\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__25947\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__5277\ : Odrv4
    port map (
            O => \N__25944\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__25941\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__5275\ : Odrv4
    port map (
            O => \N__25938\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__5274\ : Odrv4
    port map (
            O => \N__25933\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__5273\ : IoInMux
    port map (
            O => \N__25922\,
            I => \N__25919\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25916\
        );

    \I__5271\ : IoSpan4Mux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__5270\ : Span4Mux_s3_v
    port map (
            O => \N__25913\,
            I => \N__25910\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__25910\,
            I => \G_9\
        );

    \I__5268\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__25904\,
            I => \POWERLED.un1_dutycycle_172_m4_bm_sn\
        );

    \I__5266\ : InMux
    port map (
            O => \N__25901\,
            I => \N__25895\
        );

    \I__5265\ : InMux
    port map (
            O => \N__25900\,
            I => \N__25895\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__25895\,
            I => \N__25892\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__25892\,
            I => \N__25886\
        );

    \I__5262\ : InMux
    port map (
            O => \N__25891\,
            I => \N__25883\
        );

    \I__5261\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25878\
        );

    \I__5260\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25878\
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__25886\,
            I => \POWERLED.N_20_i\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__25883\,
            I => \POWERLED.N_20_i\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__25878\,
            I => \POWERLED.N_20_i\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__25871\,
            I => \N__25866\
        );

    \I__5255\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25862\
        );

    \I__5254\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25855\
        );

    \I__5253\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25855\
        );

    \I__5252\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25855\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__25862\,
            I => \N__25851\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25848\
        );

    \I__5249\ : InMux
    port map (
            O => \N__25854\,
            I => \N__25843\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__25851\,
            I => \N__25838\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__25848\,
            I => \N__25838\
        );

    \I__5246\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25833\
        );

    \I__5245\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25833\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__25843\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__5243\ : Odrv4
    port map (
            O => \N__25838\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__25833\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__5241\ : CascadeMux
    port map (
            O => \N__25826\,
            I => \POWERLED.un1_count_off_1_sqmuxa_2_0_cascade_\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__25823\,
            I => \N__25806\
        );

    \I__5239\ : InMux
    port map (
            O => \N__25822\,
            I => \N__25802\
        );

    \I__5238\ : CascadeMux
    port map (
            O => \N__25821\,
            I => \N__25798\
        );

    \I__5237\ : CascadeMux
    port map (
            O => \N__25820\,
            I => \N__25794\
        );

    \I__5236\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25788\
        );

    \I__5235\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25788\
        );

    \I__5234\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25783\
        );

    \I__5233\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25783\
        );

    \I__5232\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25775\
        );

    \I__5231\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25775\
        );

    \I__5230\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25775\
        );

    \I__5229\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25768\
        );

    \I__5228\ : InMux
    port map (
            O => \N__25811\,
            I => \N__25768\
        );

    \I__5227\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25768\
        );

    \I__5226\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25763\
        );

    \I__5225\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25760\
        );

    \I__5224\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25753\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25750\
        );

    \I__5222\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25747\
        );

    \I__5221\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25742\
        );

    \I__5220\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25742\
        );

    \I__5219\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25739\
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__25793\,
            I => \N__25735\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__25788\,
            I => \N__25729\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__25783\,
            I => \N__25724\
        );

    \I__5215\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25719\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__25775\,
            I => \N__25712\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25712\
        );

    \I__5212\ : InMux
    port map (
            O => \N__25767\,
            I => \N__25707\
        );

    \I__5211\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25707\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__25763\,
            I => \N__25702\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__25760\,
            I => \N__25702\
        );

    \I__5208\ : InMux
    port map (
            O => \N__25759\,
            I => \N__25699\
        );

    \I__5207\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25696\
        );

    \I__5206\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25691\
        );

    \I__5205\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25691\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25680\
        );

    \I__5203\ : Span4Mux_s1_v
    port map (
            O => \N__25750\,
            I => \N__25680\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__25747\,
            I => \N__25680\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__25742\,
            I => \N__25680\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__25739\,
            I => \N__25680\
        );

    \I__5199\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25677\
        );

    \I__5198\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25668\
        );

    \I__5197\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25668\
        );

    \I__5196\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25668\
        );

    \I__5195\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25668\
        );

    \I__5194\ : Span4Mux_v
    port map (
            O => \N__25729\,
            I => \N__25665\
        );

    \I__5193\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25660\
        );

    \I__5192\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25660\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__25724\,
            I => \N__25657\
        );

    \I__5190\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25652\
        );

    \I__5189\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25652\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__25719\,
            I => \N__25649\
        );

    \I__5187\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25644\
        );

    \I__5186\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25644\
        );

    \I__5185\ : Span4Mux_v
    port map (
            O => \N__25712\,
            I => \N__25637\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__25707\,
            I => \N__25637\
        );

    \I__5183\ : Span4Mux_v
    port map (
            O => \N__25702\,
            I => \N__25637\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__25699\,
            I => \N__25628\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__25696\,
            I => \N__25628\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__25691\,
            I => \N__25628\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__25680\,
            I => \N__25628\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__25677\,
            I => \N__25623\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__25668\,
            I => \N__25623\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__25665\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__25660\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__25657\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__25652\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__25649\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__25644\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__25637\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__25628\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5168\ : Odrv12
    port map (
            O => \N__25623\,
            I => \POWERLED.func_state_RNIBVNS_0Z0Z_1\
        );

    \I__5167\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25598\
        );

    \I__5166\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25598\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__25598\,
            I => \N__25591\
        );

    \I__5164\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25588\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__25596\,
            I => \N__25585\
        );

    \I__5162\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25573\
        );

    \I__5161\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25573\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__25591\,
            I => \N__25568\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__25588\,
            I => \N__25568\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25563\
        );

    \I__5157\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25563\
        );

    \I__5156\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25556\
        );

    \I__5155\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25556\
        );

    \I__5154\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25556\
        );

    \I__5153\ : InMux
    port map (
            O => \N__25580\,
            I => \N__25553\
        );

    \I__5152\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25548\
        );

    \I__5151\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25548\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__25573\,
            I => \N__25541\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__25568\,
            I => \N__25541\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__25563\,
            I => \N__25541\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__25556\,
            I => \N__25538\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__25553\,
            I => \POWERLED.N_2171_i\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__25548\,
            I => \POWERLED.N_2171_i\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__25541\,
            I => \POWERLED.N_2171_i\
        );

    \I__5143\ : Odrv12
    port map (
            O => \N__25538\,
            I => \POWERLED.N_2171_i\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__25529\,
            I => \POWERLED.un1_dutycycle_172_m3_ns_1_cascade_\
        );

    \I__5141\ : InMux
    port map (
            O => \N__25526\,
            I => \POWERLED.un1_count_clk_2_cry_11\
        );

    \I__5140\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25519\
        );

    \I__5139\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25516\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__25519\,
            I => \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__25516\,
            I => \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\
        );

    \I__5136\ : InMux
    port map (
            O => \N__25511\,
            I => \POWERLED.un1_count_clk_2_cry_12\
        );

    \I__5135\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25504\
        );

    \I__5134\ : InMux
    port map (
            O => \N__25507\,
            I => \N__25501\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__25504\,
            I => \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__25501\,
            I => \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\
        );

    \I__5131\ : InMux
    port map (
            O => \N__25496\,
            I => \POWERLED.un1_count_clk_2_cry_13\
        );

    \I__5130\ : InMux
    port map (
            O => \N__25493\,
            I => \POWERLED.un1_count_clk_2_cry_14\
        );

    \I__5129\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25486\
        );

    \I__5128\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__25486\,
            I => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__25483\,
            I => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\
        );

    \I__5125\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25475\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__25475\,
            I => \POWERLED.count_clk_0_15\
        );

    \I__5123\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25466\
        );

    \I__5122\ : InMux
    port map (
            O => \N__25471\,
            I => \N__25466\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__5120\ : Odrv4
    port map (
            O => \N__25463\,
            I => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\
        );

    \I__5119\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25457\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__25457\,
            I => \POWERLED.count_clk_0_7\
        );

    \I__5117\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25451\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25448\
        );

    \I__5115\ : Span4Mux_v
    port map (
            O => \N__25448\,
            I => \N__25444\
        );

    \I__5114\ : InMux
    port map (
            O => \N__25447\,
            I => \N__25441\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__25444\,
            I => \POWERLED.N_392\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__25441\,
            I => \POWERLED.N_392\
        );

    \I__5111\ : CascadeMux
    port map (
            O => \N__25436\,
            I => \N__25433\
        );

    \I__5110\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25429\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__25432\,
            I => \N__25426\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__25429\,
            I => \N__25423\
        );

    \I__5107\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25420\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__25423\,
            I => \N__25417\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__25420\,
            I => \POWERLED.mult1_un40_sum_i_5\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__25417\,
            I => \POWERLED.mult1_un40_sum_i_5\
        );

    \I__5103\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25408\
        );

    \I__5102\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25405\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__25408\,
            I => \N__25402\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__25405\,
            I => \N__25399\
        );

    \I__5099\ : Span4Mux_h
    port map (
            O => \N__25402\,
            I => \N__25396\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__25399\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__25396\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__5096\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25387\
        );

    \I__5095\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25384\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__25387\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__25384\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__5092\ : InMux
    port map (
            O => \N__25379\,
            I => \POWERLED.un1_count_clk_2_cry_2\
        );

    \I__5091\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25372\
        );

    \I__5090\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25369\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__25372\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__25369\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__5087\ : InMux
    port map (
            O => \N__25364\,
            I => \POWERLED.un1_count_clk_2_cry_3\
        );

    \I__5086\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25355\
        );

    \I__5085\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25355\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__25355\,
            I => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\
        );

    \I__5083\ : InMux
    port map (
            O => \N__25352\,
            I => \POWERLED.un1_count_clk_2_cry_4\
        );

    \I__5082\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25343\
        );

    \I__5081\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25343\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__25343\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__5079\ : InMux
    port map (
            O => \N__25340\,
            I => \POWERLED.un1_count_clk_2_cry_5\
        );

    \I__5078\ : InMux
    port map (
            O => \N__25337\,
            I => \POWERLED.un1_count_clk_2_cry_6\
        );

    \I__5077\ : InMux
    port map (
            O => \N__25334\,
            I => \N__25328\
        );

    \I__5076\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25328\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__25328\,
            I => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\
        );

    \I__5074\ : InMux
    port map (
            O => \N__25325\,
            I => \POWERLED.un1_count_clk_2_cry_7_cZ0\
        );

    \I__5073\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25316\
        );

    \I__5072\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25316\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__25316\,
            I => \N__25313\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__25313\,
            I => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\
        );

    \I__5069\ : InMux
    port map (
            O => \N__25310\,
            I => \bfn_9_8_0_\
        );

    \I__5068\ : InMux
    port map (
            O => \N__25307\,
            I => \POWERLED.un1_count_clk_2_cry_9_cZ0\
        );

    \I__5067\ : InMux
    port map (
            O => \N__25304\,
            I => \POWERLED.un1_count_clk_2_cry_10_cZ0\
        );

    \I__5066\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__25298\,
            I => \POWERLED.count_clk_0_5\
        );

    \I__5064\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25292\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__25292\,
            I => \POWERLED.count_clk_0_6\
        );

    \I__5062\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25286\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__25286\,
            I => \POWERLED.count_clk_0_8\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25280\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__25280\,
            I => \POWERLED.count_clk_0_9\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__25277\,
            I => \N__25273\
        );

    \I__5057\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25270\
        );

    \I__5056\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25267\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__25270\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__25267\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__5053\ : InMux
    port map (
            O => \N__25262\,
            I => \POWERLED.un1_count_clk_2_cry_1\
        );

    \I__5052\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25256\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__25256\,
            I => \POWERLED.un34_clk_100khz_5\
        );

    \I__5050\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25250\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__25250\,
            I => \N__25244\
        );

    \I__5048\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25237\
        );

    \I__5047\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25237\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25237\
        );

    \I__5045\ : Span4Mux_h
    port map (
            O => \N__25244\,
            I => \N__25232\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__25237\,
            I => \N__25232\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__25226\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__5039\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25215\
        );

    \I__5038\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25208\
        );

    \I__5037\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25208\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__25215\,
            I => \N__25205\
        );

    \I__5035\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25200\
        );

    \I__5034\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25200\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__25208\,
            I => \N__25197\
        );

    \I__5032\ : Odrv12
    port map (
            O => \N__25205\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__25200\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__5030\ : Odrv4
    port map (
            O => \N__25197\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__5029\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25184\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__25184\,
            I => \N__25178\
        );

    \I__5026\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25175\
        );

    \I__5025\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25170\
        );

    \I__5024\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25170\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__25178\,
            I => \POWERLED.count_RNIZ0Z_15\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__25175\,
            I => \POWERLED.count_RNIZ0Z_15\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__25170\,
            I => \POWERLED.count_RNIZ0Z_15\
        );

    \I__5020\ : InMux
    port map (
            O => \N__25163\,
            I => \N__25160\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__25160\,
            I => \N__25157\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__25154\,
            I => \POWERLED.curr_state_1_0\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__25151\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1_cascade_\
        );

    \I__5015\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__25145\,
            I => \N__25142\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__25142\,
            I => \N__25137\
        );

    \I__5012\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25133\
        );

    \I__5011\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25130\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__25137\,
            I => \N__25127\
        );

    \I__5009\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25124\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__25133\,
            I => \N__25121\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__25130\,
            I => \N__25118\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__25127\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__25124\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__25121\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__5003\ : Odrv4
    port map (
            O => \N__25118\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__25106\,
            I => \N__25103\
        );

    \I__5000\ : Odrv12
    port map (
            O => \N__25103\,
            I => \POWERLED.count_0_1\
        );

    \I__4999\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25095\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__25099\,
            I => \N__25092\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__25098\,
            I => \N__25088\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25085\
        );

    \I__4995\ : InMux
    port map (
            O => \N__25092\,
            I => \N__25079\
        );

    \I__4994\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25079\
        );

    \I__4993\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25075\
        );

    \I__4992\ : Span4Mux_s3_h
    port map (
            O => \N__25085\,
            I => \N__25072\
        );

    \I__4991\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25069\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25066\
        );

    \I__4989\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25063\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__25075\,
            I => \N__25060\
        );

    \I__4987\ : Span4Mux_v
    port map (
            O => \N__25072\,
            I => \N__25051\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__25069\,
            I => \N__25051\
        );

    \I__4985\ : Span4Mux_h
    port map (
            O => \N__25066\,
            I => \N__25051\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__25063\,
            I => \N__25051\
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__25060\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__25051\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__4981\ : InMux
    port map (
            O => \N__25046\,
            I => \N__25027\
        );

    \I__4980\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25024\
        );

    \I__4979\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25021\
        );

    \I__4978\ : InMux
    port map (
            O => \N__25043\,
            I => \N__25014\
        );

    \I__4977\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25014\
        );

    \I__4976\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25014\
        );

    \I__4975\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25005\
        );

    \I__4974\ : InMux
    port map (
            O => \N__25039\,
            I => \N__25005\
        );

    \I__4973\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25005\
        );

    \I__4972\ : InMux
    port map (
            O => \N__25037\,
            I => \N__25005\
        );

    \I__4971\ : InMux
    port map (
            O => \N__25036\,
            I => \N__24998\
        );

    \I__4970\ : InMux
    port map (
            O => \N__25035\,
            I => \N__24998\
        );

    \I__4969\ : InMux
    port map (
            O => \N__25034\,
            I => \N__24998\
        );

    \I__4968\ : InMux
    port map (
            O => \N__25033\,
            I => \N__24989\
        );

    \I__4967\ : InMux
    port map (
            O => \N__25032\,
            I => \N__24989\
        );

    \I__4966\ : InMux
    port map (
            O => \N__25031\,
            I => \N__24989\
        );

    \I__4965\ : InMux
    port map (
            O => \N__25030\,
            I => \N__24989\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__25027\,
            I => \N__24986\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__25024\,
            I => \N__24981\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__25021\,
            I => \N__24981\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__25014\,
            I => \N__24972\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__24972\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__24998\,
            I => \N__24972\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24972\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__24986\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__4956\ : Odrv12
    port map (
            O => \N__24981\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__24972\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__4954\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24962\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__4952\ : Odrv12
    port map (
            O => \N__24959\,
            I => \POWERLED.count_0_0\
        );

    \I__4951\ : CascadeMux
    port map (
            O => \N__24956\,
            I => \N__24947\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__24955\,
            I => \N__24943\
        );

    \I__4949\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24935\
        );

    \I__4948\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24935\
        );

    \I__4947\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24935\
        );

    \I__4946\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24930\
        );

    \I__4945\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24930\
        );

    \I__4944\ : InMux
    port map (
            O => \N__24947\,
            I => \N__24923\
        );

    \I__4943\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24923\
        );

    \I__4942\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24923\
        );

    \I__4941\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24919\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__24935\,
            I => \N__24916\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__24930\,
            I => \N__24911\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__24923\,
            I => \N__24911\
        );

    \I__4937\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24908\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24903\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__24916\,
            I => \N__24900\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__24911\,
            I => \N__24895\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__24908\,
            I => \N__24895\
        );

    \I__4932\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24890\
        );

    \I__4931\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24890\
        );

    \I__4930\ : Span4Mux_v
    port map (
            O => \N__24903\,
            I => \N__24887\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__24900\,
            I => \N__24882\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__24895\,
            I => \N__24882\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__24890\,
            I => \N__24879\
        );

    \I__4926\ : Sp12to4
    port map (
            O => \N__24887\,
            I => \N__24876\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__24882\,
            I => \N__24873\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__24879\,
            I => \N__24870\
        );

    \I__4923\ : Span12Mux_s8_h
    port map (
            O => \N__24876\,
            I => \N__24867\
        );

    \I__4922\ : Span4Mux_v
    port map (
            O => \N__24873\,
            I => \N__24862\
        );

    \I__4921\ : Span4Mux_v
    port map (
            O => \N__24870\,
            I => \N__24862\
        );

    \I__4920\ : Odrv12
    port map (
            O => \N__24867\,
            I => slp_s4n
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__24862\,
            I => slp_s4n
        );

    \I__4918\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24854\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__24854\,
            I => \N__24850\
        );

    \I__4916\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24846\
        );

    \I__4915\ : Span4Mux_h
    port map (
            O => \N__24850\,
            I => \N__24841\
        );

    \I__4914\ : InMux
    port map (
            O => \N__24849\,
            I => \N__24838\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__24846\,
            I => \N__24835\
        );

    \I__4912\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24832\
        );

    \I__4911\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24829\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__24841\,
            I => \N__24826\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__24838\,
            I => \N__24821\
        );

    \I__4908\ : Span4Mux_v
    port map (
            O => \N__24835\,
            I => \N__24821\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__24832\,
            I => \N__24816\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24816\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__24826\,
            I => \RSMRST_PWRGD_RSMRSTn_2_fast\
        );

    \I__4904\ : Odrv4
    port map (
            O => \N__24821\,
            I => \RSMRST_PWRGD_RSMRSTn_2_fast\
        );

    \I__4903\ : Odrv12
    port map (
            O => \N__24816\,
            I => \RSMRST_PWRGD_RSMRSTn_2_fast\
        );

    \I__4902\ : InMux
    port map (
            O => \N__24809\,
            I => \N__24804\
        );

    \I__4901\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24801\
        );

    \I__4900\ : InMux
    port map (
            O => \N__24807\,
            I => \N__24798\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__24804\,
            I => \N__24791\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__24801\,
            I => \N__24791\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__24798\,
            I => \N__24791\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__24791\,
            I => \POWERLED.N_150_i\
        );

    \I__4895\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__24785\,
            I => \N__24782\
        );

    \I__4893\ : Span4Mux_h
    port map (
            O => \N__24782\,
            I => \N__24774\
        );

    \I__4892\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24771\
        );

    \I__4891\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24768\
        );

    \I__4890\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24765\
        );

    \I__4889\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24762\
        );

    \I__4888\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24759\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__24774\,
            I => \POWERLED.N_154\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__24771\,
            I => \POWERLED.N_154\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__24768\,
            I => \POWERLED.N_154\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__24765\,
            I => \POWERLED.N_154\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__24762\,
            I => \POWERLED.N_154\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__24759\,
            I => \POWERLED.N_154\
        );

    \I__4881\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24743\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__24743\,
            I => \POWERLED.N_389\
        );

    \I__4879\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24737\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__24737\,
            I => \POWERLED.count_off_0_10\
        );

    \I__4877\ : InMux
    port map (
            O => \N__24734\,
            I => \N__24728\
        );

    \I__4876\ : InMux
    port map (
            O => \N__24733\,
            I => \N__24728\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__24728\,
            I => \POWERLED.count_off_1_9\
        );

    \I__4874\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24719\
        );

    \I__4873\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24719\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__24719\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__24716\,
            I => \POWERLED.count_offZ0Z_10_cascade_\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__24713\,
            I => \POWERLED.un34_clk_100khz_4_cascade_\
        );

    \I__4869\ : InMux
    port map (
            O => \N__24710\,
            I => \N__24706\
        );

    \I__4868\ : InMux
    port map (
            O => \N__24709\,
            I => \N__24703\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__24706\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__24703\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__4865\ : InMux
    port map (
            O => \N__24698\,
            I => \HDA_STRAP.un1_count_1_cry_12\
        );

    \I__4864\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24691\
        );

    \I__4863\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24688\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__24691\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__24688\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__4860\ : InMux
    port map (
            O => \N__24683\,
            I => \HDA_STRAP.un1_count_1_cry_13\
        );

    \I__4859\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24676\
        );

    \I__4858\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24673\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__24676\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__24673\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__4855\ : InMux
    port map (
            O => \N__24668\,
            I => \HDA_STRAP.un1_count_1_cry_14\
        );

    \I__4854\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24661\
        );

    \I__4853\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24658\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__24661\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__24658\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__4850\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24650\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__24650\,
            I => \HDA_STRAP.count_RNO_0Z0Z_16\
        );

    \I__4848\ : InMux
    port map (
            O => \N__24647\,
            I => \bfn_9_3_0_\
        );

    \I__4847\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__24638\,
            I => \N__24634\
        );

    \I__4844\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24631\
        );

    \I__4843\ : Odrv4
    port map (
            O => \N__24634\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__24631\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__4841\ : InMux
    port map (
            O => \N__24626\,
            I => \HDA_STRAP.un1_count_1_cry_16\
        );

    \I__4840\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24620\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__4838\ : Span4Mux_s2_v
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__24614\,
            I => \HDA_STRAP.count_RNO_0Z0Z_17\
        );

    \I__4836\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__24605\,
            I => \POWERLED.un1_func_state25_6_0_a2_1\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__24602\,
            I => \POWERLED.un1_func_state25_6_0_o_N_305_N_cascade_\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__24599\,
            I => \POWERLED.un1_func_state25_6_0_0_cascade_\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__24596\,
            I => \N__24593\
        );

    \I__4830\ : InMux
    port map (
            O => \N__24593\,
            I => \N__24590\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__24590\,
            I => \POWERLED.un1_func_state25_6_0_1\
        );

    \I__4828\ : InMux
    port map (
            O => \N__24587\,
            I => \HDA_STRAP.un1_count_1_cry_3\
        );

    \I__4827\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24580\
        );

    \I__4826\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24577\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__24580\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__24577\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__4823\ : InMux
    port map (
            O => \N__24572\,
            I => \HDA_STRAP.un1_count_1_cry_4\
        );

    \I__4822\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24565\
        );

    \I__4821\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24562\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__24565\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__24562\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__4818\ : CascadeMux
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__4817\ : InMux
    port map (
            O => \N__24554\,
            I => \N__24551\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__24551\,
            I => \HDA_STRAP.count_RNO_0Z0Z_6\
        );

    \I__4815\ : InMux
    port map (
            O => \N__24548\,
            I => \HDA_STRAP.un1_count_1_cry_5\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__24545\,
            I => \N__24542\
        );

    \I__4813\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__24539\,
            I => \N__24535\
        );

    \I__4811\ : InMux
    port map (
            O => \N__24538\,
            I => \N__24532\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__24535\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__24532\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__4808\ : InMux
    port map (
            O => \N__24527\,
            I => \HDA_STRAP.un1_count_1_cry_6\
        );

    \I__4807\ : CascadeMux
    port map (
            O => \N__24524\,
            I => \N__24521\
        );

    \I__4806\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24517\
        );

    \I__4805\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24514\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__24517\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__24514\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__4802\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24506\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__24506\,
            I => \HDA_STRAP.count_RNO_0Z0Z_8\
        );

    \I__4800\ : InMux
    port map (
            O => \N__24503\,
            I => \bfn_9_2_0_\
        );

    \I__4799\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24496\
        );

    \I__4798\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24493\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__24496\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__24493\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__4795\ : InMux
    port map (
            O => \N__24488\,
            I => \HDA_STRAP.un1_count_1_cry_8\
        );

    \I__4794\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24481\
        );

    \I__4793\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__24481\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__24478\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__24473\,
            I => \N__24470\
        );

    \I__4789\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__24467\,
            I => \HDA_STRAP.count_RNO_0Z0Z_10\
        );

    \I__4787\ : InMux
    port map (
            O => \N__24464\,
            I => \HDA_STRAP.un1_count_1_cry_9\
        );

    \I__4786\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24457\
        );

    \I__4785\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24454\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__24457\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__24454\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__4782\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__24446\,
            I => \HDA_STRAP.count_RNO_0Z0Z_11\
        );

    \I__4780\ : InMux
    port map (
            O => \N__24443\,
            I => \HDA_STRAP.un1_count_1_cry_10\
        );

    \I__4779\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24436\
        );

    \I__4778\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24433\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__24436\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__24433\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__4775\ : InMux
    port map (
            O => \N__24428\,
            I => \HDA_STRAP.un1_count_1_cry_11\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__24425\,
            I => \N__24417\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__24424\,
            I => \N__24410\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__24423\,
            I => \N__24407\
        );

    \I__4771\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24403\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__24421\,
            I => \N__24399\
        );

    \I__4769\ : CascadeMux
    port map (
            O => \N__24420\,
            I => \N__24395\
        );

    \I__4768\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24389\
        );

    \I__4767\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24389\
        );

    \I__4766\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24383\
        );

    \I__4765\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24378\
        );

    \I__4764\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24378\
        );

    \I__4763\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24373\
        );

    \I__4762\ : InMux
    port map (
            O => \N__24407\,
            I => \N__24373\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__24406\,
            I => \N__24370\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__24403\,
            I => \N__24367\
        );

    \I__4759\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24358\
        );

    \I__4758\ : InMux
    port map (
            O => \N__24399\,
            I => \N__24358\
        );

    \I__4757\ : InMux
    port map (
            O => \N__24398\,
            I => \N__24358\
        );

    \I__4756\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24358\
        );

    \I__4755\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24353\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__24389\,
            I => \N__24350\
        );

    \I__4753\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24345\
        );

    \I__4752\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24345\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__24386\,
            I => \N__24339\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__24383\,
            I => \N__24334\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__24378\,
            I => \N__24334\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__24373\,
            I => \N__24331\
        );

    \I__4747\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24328\
        );

    \I__4746\ : Span4Mux_v
    port map (
            O => \N__24367\,
            I => \N__24323\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24323\
        );

    \I__4744\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24318\
        );

    \I__4743\ : InMux
    port map (
            O => \N__24356\,
            I => \N__24318\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__24353\,
            I => \N__24311\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__24350\,
            I => \N__24311\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24311\
        );

    \I__4739\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24302\
        );

    \I__4738\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24302\
        );

    \I__4737\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24302\
        );

    \I__4736\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24302\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__24334\,
            I => \N__24295\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__24331\,
            I => \N__24295\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__24328\,
            I => \N__24295\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__24323\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__24318\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__24311\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__24302\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__24295\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__4727\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24276\
        );

    \I__4726\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24271\
        );

    \I__4725\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24271\
        );

    \I__4724\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24260\
        );

    \I__4723\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24255\
        );

    \I__4722\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24255\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__24276\,
            I => \N__24250\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__24271\,
            I => \N__24250\
        );

    \I__4719\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24241\
        );

    \I__4718\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24241\
        );

    \I__4717\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24241\
        );

    \I__4716\ : InMux
    port map (
            O => \N__24267\,
            I => \N__24238\
        );

    \I__4715\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24235\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__24265\,
            I => \N__24232\
        );

    \I__4713\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24229\
        );

    \I__4712\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24226\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__24260\,
            I => \N__24223\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__24255\,
            I => \N__24218\
        );

    \I__4709\ : Span4Mux_v
    port map (
            O => \N__24250\,
            I => \N__24218\
        );

    \I__4708\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24213\
        );

    \I__4707\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24213\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__24241\,
            I => \N__24206\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__24238\,
            I => \N__24206\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__24235\,
            I => \N__24206\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24203\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__24229\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__24226\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__24223\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__24218\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__24213\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__24206\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__24203\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__24188\,
            I => \POWERLED.g0_i_a6_0_1_cascade_\
        );

    \I__4694\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24182\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__24182\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_12\
        );

    \I__4692\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24172\
        );

    \I__4690\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24169\
        );

    \I__4689\ : Span4Mux_s2_v
    port map (
            O => \N__24172\,
            I => \N__24164\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__24169\,
            I => \N__24161\
        );

    \I__4687\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24153\
        );

    \I__4686\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24149\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__24164\,
            I => \N__24146\
        );

    \I__4684\ : Span4Mux_h
    port map (
            O => \N__24161\,
            I => \N__24143\
        );

    \I__4683\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24136\
        );

    \I__4682\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24136\
        );

    \I__4681\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24136\
        );

    \I__4680\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24131\
        );

    \I__4679\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24131\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__24153\,
            I => \N__24128\
        );

    \I__4677\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24125\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__24149\,
            I => \N__24122\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__24146\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__24143\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__24136\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__24131\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__4671\ : Odrv12
    port map (
            O => \N__24128\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__24125\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__4669\ : Odrv4
    port map (
            O => \N__24122\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__24107\,
            I => \N__24101\
        );

    \I__4667\ : InMux
    port map (
            O => \N__24106\,
            I => \N__24094\
        );

    \I__4666\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24094\
        );

    \I__4665\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24091\
        );

    \I__4664\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24088\
        );

    \I__4663\ : CascadeMux
    port map (
            O => \N__24100\,
            I => \N__24084\
        );

    \I__4662\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24077\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__24094\,
            I => \N__24074\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__24091\,
            I => \N__24069\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__24088\,
            I => \N__24069\
        );

    \I__4658\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24066\
        );

    \I__4657\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24063\
        );

    \I__4656\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24056\
        );

    \I__4655\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24056\
        );

    \I__4654\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24056\
        );

    \I__4653\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24053\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__24077\,
            I => \N__24050\
        );

    \I__4651\ : Span4Mux_s3_v
    port map (
            O => \N__24074\,
            I => \N__24047\
        );

    \I__4650\ : Span12Mux_s7_h
    port map (
            O => \N__24069\,
            I => \N__24036\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__24066\,
            I => \N__24036\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24036\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__24056\,
            I => \N__24036\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__24053\,
            I => \N__24036\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__24050\,
            I => \N__24033\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__24047\,
            I => \N__24030\
        );

    \I__4643\ : Span12Mux_s5_v
    port map (
            O => \N__24036\,
            I => \N__24027\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__24033\,
            I => \POWERLED.func_state_RNIC4OR2Z0Z_0\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__24030\,
            I => \POWERLED.func_state_RNIC4OR2Z0Z_0\
        );

    \I__4640\ : Odrv12
    port map (
            O => \N__24027\,
            I => \POWERLED.func_state_RNIC4OR2Z0Z_0\
        );

    \I__4639\ : InMux
    port map (
            O => \N__24020\,
            I => \N__24014\
        );

    \I__4638\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24014\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__24014\,
            I => \N__24005\
        );

    \I__4636\ : InMux
    port map (
            O => \N__24013\,
            I => \N__24001\
        );

    \I__4635\ : InMux
    port map (
            O => \N__24012\,
            I => \N__23996\
        );

    \I__4634\ : InMux
    port map (
            O => \N__24011\,
            I => \N__23996\
        );

    \I__4633\ : InMux
    port map (
            O => \N__24010\,
            I => \N__23989\
        );

    \I__4632\ : InMux
    port map (
            O => \N__24009\,
            I => \N__23989\
        );

    \I__4631\ : InMux
    port map (
            O => \N__24008\,
            I => \N__23989\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__24005\,
            I => \N__23986\
        );

    \I__4629\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23983\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__24001\,
            I => \N__23976\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__23996\,
            I => \N__23976\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23976\
        );

    \I__4625\ : Span4Mux_h
    port map (
            O => \N__23986\,
            I => \N__23971\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23966\
        );

    \I__4623\ : Span4Mux_v
    port map (
            O => \N__23976\,
            I => \N__23966\
        );

    \I__4622\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23961\
        );

    \I__4621\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23961\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__23971\,
            I => \POWERLED.N_390\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__23966\,
            I => \POWERLED.N_390\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__23961\,
            I => \POWERLED.N_390\
        );

    \I__4617\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23941\
        );

    \I__4616\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23938\
        );

    \I__4615\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23935\
        );

    \I__4614\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23932\
        );

    \I__4613\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23929\
        );

    \I__4612\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23926\
        );

    \I__4611\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23923\
        );

    \I__4610\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23916\
        );

    \I__4609\ : InMux
    port map (
            O => \N__23946\,
            I => \N__23916\
        );

    \I__4608\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23916\
        );

    \I__4607\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23913\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__23941\,
            I => \N__23910\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__23938\,
            I => \N__23905\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23905\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__23932\,
            I => \N__23900\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23897\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__23926\,
            I => \N__23894\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__23923\,
            I => \N__23888\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__23916\,
            I => \N__23885\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__23913\,
            I => \N__23879\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__23910\,
            I => \N__23874\
        );

    \I__4596\ : Span4Mux_v
    port map (
            O => \N__23905\,
            I => \N__23874\
        );

    \I__4595\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23871\
        );

    \I__4594\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23868\
        );

    \I__4593\ : Span4Mux_h
    port map (
            O => \N__23900\,
            I => \N__23863\
        );

    \I__4592\ : Span4Mux_s2_v
    port map (
            O => \N__23897\,
            I => \N__23863\
        );

    \I__4591\ : Span4Mux_v
    port map (
            O => \N__23894\,
            I => \N__23860\
        );

    \I__4590\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23857\
        );

    \I__4589\ : InMux
    port map (
            O => \N__23892\,
            I => \N__23852\
        );

    \I__4588\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23852\
        );

    \I__4587\ : Span4Mux_h
    port map (
            O => \N__23888\,
            I => \N__23847\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__23885\,
            I => \N__23847\
        );

    \I__4585\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23840\
        );

    \I__4584\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23840\
        );

    \I__4583\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23840\
        );

    \I__4582\ : Span4Mux_v
    port map (
            O => \N__23879\,
            I => \N__23829\
        );

    \I__4581\ : Span4Mux_v
    port map (
            O => \N__23874\,
            I => \N__23829\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__23871\,
            I => \N__23829\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__23868\,
            I => \N__23829\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__23863\,
            I => \N__23829\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__23860\,
            I => \POWERLED.N_209\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__23857\,
            I => \POWERLED.N_209\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__23852\,
            I => \POWERLED.N_209\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__23847\,
            I => \POWERLED.N_209\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__23840\,
            I => \POWERLED.N_209\
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__23829\,
            I => \POWERLED.N_209\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__23816\,
            I => \POWERLED.N_145_N_cascade_\
        );

    \I__4570\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23801\
        );

    \I__4569\ : InMux
    port map (
            O => \N__23812\,
            I => \N__23798\
        );

    \I__4568\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23793\
        );

    \I__4567\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23793\
        );

    \I__4566\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23790\
        );

    \I__4565\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23784\
        );

    \I__4564\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23784\
        );

    \I__4563\ : IoInMux
    port map (
            O => \N__23806\,
            I => \N__23781\
        );

    \I__4562\ : InMux
    port map (
            O => \N__23805\,
            I => \N__23772\
        );

    \I__4561\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23772\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23765\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23765\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__23793\,
            I => \N__23765\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__23790\,
            I => \N__23762\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__23789\,
            I => \N__23759\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23752\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__23781\,
            I => \N__23752\
        );

    \I__4553\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23743\
        );

    \I__4552\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23743\
        );

    \I__4551\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23743\
        );

    \I__4550\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23743\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23734\
        );

    \I__4548\ : Span4Mux_s3_v
    port map (
            O => \N__23765\,
            I => \N__23729\
        );

    \I__4547\ : Span4Mux_s3_v
    port map (
            O => \N__23762\,
            I => \N__23729\
        );

    \I__4546\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23722\
        );

    \I__4545\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23722\
        );

    \I__4544\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23722\
        );

    \I__4543\ : Span4Mux_s3_h
    port map (
            O => \N__23752\,
            I => \N__23717\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__23743\,
            I => \N__23717\
        );

    \I__4541\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23712\
        );

    \I__4540\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23712\
        );

    \I__4539\ : InMux
    port map (
            O => \N__23740\,
            I => \N__23707\
        );

    \I__4538\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23707\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__23738\,
            I => \N__23704\
        );

    \I__4536\ : InMux
    port map (
            O => \N__23737\,
            I => \N__23700\
        );

    \I__4535\ : Span4Mux_v
    port map (
            O => \N__23734\,
            I => \N__23696\
        );

    \I__4534\ : Span4Mux_v
    port map (
            O => \N__23729\,
            I => \N__23688\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__23722\,
            I => \N__23688\
        );

    \I__4532\ : Span4Mux_h
    port map (
            O => \N__23717\,
            I => \N__23688\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__23712\,
            I => \N__23683\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__23707\,
            I => \N__23683\
        );

    \I__4529\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23678\
        );

    \I__4528\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23678\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23675\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__23699\,
            I => \N__23672\
        );

    \I__4525\ : Span4Mux_v
    port map (
            O => \N__23696\,
            I => \N__23669\
        );

    \I__4524\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23666\
        );

    \I__4523\ : Span4Mux_v
    port map (
            O => \N__23688\,
            I => \N__23663\
        );

    \I__4522\ : Sp12to4
    port map (
            O => \N__23683\,
            I => \N__23656\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__23678\,
            I => \N__23656\
        );

    \I__4520\ : Span12Mux_s3_v
    port map (
            O => \N__23675\,
            I => \N__23656\
        );

    \I__4519\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23653\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__23669\,
            I => \G_154\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__23666\,
            I => \G_154\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__23663\,
            I => \G_154\
        );

    \I__4515\ : Odrv12
    port map (
            O => \N__23656\,
            I => \G_154\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23653\,
            I => \G_154\
        );

    \I__4513\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__23636\,
            I => \N__23632\
        );

    \I__4510\ : InMux
    port map (
            O => \N__23635\,
            I => \N__23629\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__23632\,
            I => \POWERLED.dutycycle_en_9\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__23629\,
            I => \POWERLED.dutycycle_en_9\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__4506\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23617\
        );

    \I__4505\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23614\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__23617\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__23614\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__4502\ : CascadeMux
    port map (
            O => \N__23609\,
            I => \N__23605\
        );

    \I__4501\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23602\
        );

    \I__4500\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23599\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__23602\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_1\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__23599\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_1\
        );

    \I__4497\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23591\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__23591\,
            I => \HDA_STRAP.count_RNO_0Z0Z_0\
        );

    \I__4495\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23584\
        );

    \I__4494\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23581\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23584\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__23581\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__4491\ : InMux
    port map (
            O => \N__23576\,
            I => \HDA_STRAP.un1_count_1_cry_0\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__4489\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23566\
        );

    \I__4488\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23563\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__23566\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__23563\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__4485\ : InMux
    port map (
            O => \N__23558\,
            I => \HDA_STRAP.un1_count_1_cry_1\
        );

    \I__4484\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23551\
        );

    \I__4483\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__23551\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__23548\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__4480\ : InMux
    port map (
            O => \N__23543\,
            I => \HDA_STRAP.un1_count_1_cry_2\
        );

    \I__4479\ : InMux
    port map (
            O => \N__23540\,
            I => \N__23536\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23539\,
            I => \N__23533\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__23536\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__23533\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__23528\,
            I => \POWERLED.count_clk_RNIBVNSZ0Z_4_cascade_\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__23525\,
            I => \N__23522\
        );

    \I__4473\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23516\
        );

    \I__4472\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23516\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__23516\,
            I => \POWERLED.dutycycle_eena_2\
        );

    \I__4470\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23509\
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__23512\,
            I => \N__23506\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__23509\,
            I => \N__23503\
        );

    \I__4467\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23500\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__23503\,
            I => \N__23497\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__23500\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__23497\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__4463\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23489\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23485\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__23488\,
            I => \N__23482\
        );

    \I__4460\ : Span4Mux_h
    port map (
            O => \N__23485\,
            I => \N__23479\
        );

    \I__4459\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23476\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__23479\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__23476\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\
        );

    \I__4456\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23462\
        );

    \I__4455\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23457\
        );

    \I__4454\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23457\
        );

    \I__4453\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23454\
        );

    \I__4452\ : InMux
    port map (
            O => \N__23467\,
            I => \N__23450\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__23466\,
            I => \N__23446\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__23465\,
            I => \N__23443\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__23462\,
            I => \N__23435\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23435\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23435\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__23453\,
            I => \N__23430\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23427\
        );

    \I__4444\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23422\
        );

    \I__4443\ : InMux
    port map (
            O => \N__23446\,
            I => \N__23422\
        );

    \I__4442\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23417\
        );

    \I__4441\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23417\
        );

    \I__4440\ : Span4Mux_h
    port map (
            O => \N__23435\,
            I => \N__23414\
        );

    \I__4439\ : InMux
    port map (
            O => \N__23434\,
            I => \N__23409\
        );

    \I__4438\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23409\
        );

    \I__4437\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23406\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__23427\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__23422\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__23417\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__23414\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__23409\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__23406\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__23393\,
            I => \POWERLED.dutycycleZ0Z_7_cascade_\
        );

    \I__4429\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__23387\,
            I => \POWERLED.un1_dutycycle_53_50_3\
        );

    \I__4427\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23375\
        );

    \I__4425\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23372\
        );

    \I__4424\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23368\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__23378\,
            I => \N__23363\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__23375\,
            I => \N__23358\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__23372\,
            I => \N__23358\
        );

    \I__4420\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23355\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__23368\,
            I => \N__23352\
        );

    \I__4418\ : InMux
    port map (
            O => \N__23367\,
            I => \N__23349\
        );

    \I__4417\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23344\
        );

    \I__4416\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23344\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__23358\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__23355\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__4413\ : Odrv12
    port map (
            O => \N__23352\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__23349\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__23344\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__23333\,
            I => \POWERLED.un1_dutycycle_53_51_0_cascade_\
        );

    \I__4409\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__4407\ : Span4Mux_h
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__23321\,
            I => \POWERLED.un1_dutycycle_53_50_4\
        );

    \I__4405\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__4403\ : Span4Mux_h
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__23309\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_15\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__4400\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23294\
        );

    \I__4398\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23289\
        );

    \I__4397\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23289\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__23297\,
            I => \N__23286\
        );

    \I__4395\ : Span4Mux_s3_v
    port map (
            O => \N__23294\,
            I => \N__23283\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__23289\,
            I => \N__23280\
        );

    \I__4393\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23277\
        );

    \I__4392\ : Span4Mux_v
    port map (
            O => \N__23283\,
            I => \N__23274\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__23280\,
            I => \N__23269\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__23277\,
            I => \N__23269\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__23274\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_1\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__23269\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_1\
        );

    \I__4387\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23251\
        );

    \I__4385\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23246\
        );

    \I__4384\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23237\
        );

    \I__4383\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23237\
        );

    \I__4382\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23237\
        );

    \I__4381\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23232\
        );

    \I__4380\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23232\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__23254\,
            I => \N__23225\
        );

    \I__4378\ : Span4Mux_v
    port map (
            O => \N__23251\,
            I => \N__23222\
        );

    \I__4377\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23217\
        );

    \I__4376\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23217\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23214\
        );

    \I__4374\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23209\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23209\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__23237\,
            I => \N__23204\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__23232\,
            I => \N__23204\
        );

    \I__4370\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23201\
        );

    \I__4369\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23194\
        );

    \I__4368\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23194\
        );

    \I__4367\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23194\
        );

    \I__4366\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23191\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__23222\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__23217\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__23214\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__23209\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__23204\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__23201\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__23194\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__23191\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__4357\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__23171\,
            I => \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_1\
        );

    \I__4355\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23165\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__23165\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_7\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__4352\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__23156\,
            I => \POWERLED.N_8_1\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__23153\,
            I => \N__23150\
        );

    \I__4349\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__23147\,
            I => \N__23144\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__23141\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__23138\,
            I => \N__23135\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23135\,
            I => \N__23121\
        );

    \I__4343\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23121\
        );

    \I__4342\ : InMux
    port map (
            O => \N__23133\,
            I => \N__23121\
        );

    \I__4341\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23112\
        );

    \I__4340\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23112\
        );

    \I__4339\ : InMux
    port map (
            O => \N__23130\,
            I => \N__23112\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__23129\,
            I => \N__23109\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__23128\,
            I => \N__23101\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__23121\,
            I => \N__23096\
        );

    \I__4335\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23091\
        );

    \I__4334\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23091\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__23112\,
            I => \N__23088\
        );

    \I__4332\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23085\
        );

    \I__4331\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23082\
        );

    \I__4330\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23073\
        );

    \I__4329\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23073\
        );

    \I__4328\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23073\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23073\
        );

    \I__4326\ : InMux
    port map (
            O => \N__23101\,
            I => \N__23066\
        );

    \I__4325\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23066\
        );

    \I__4324\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23066\
        );

    \I__4323\ : Span4Mux_h
    port map (
            O => \N__23096\,
            I => \N__23057\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__23091\,
            I => \N__23057\
        );

    \I__4321\ : Span4Mux_h
    port map (
            O => \N__23088\,
            I => \N__23057\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__23085\,
            I => \N__23057\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__23082\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__23073\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__23066\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__23057\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__23048\,
            I => \POWERLED.dutycycleZ0Z_9_cascade_\
        );

    \I__4314\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23041\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__23044\,
            I => \N__23037\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__23041\,
            I => \N__23031\
        );

    \I__4311\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23028\
        );

    \I__4310\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23023\
        );

    \I__4309\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23023\
        );

    \I__4308\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23017\
        );

    \I__4307\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23014\
        );

    \I__4306\ : Span4Mux_h
    port map (
            O => \N__23031\,
            I => \N__23009\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__23028\,
            I => \N__23009\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__23023\,
            I => \N__23006\
        );

    \I__4303\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23001\
        );

    \I__4302\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23001\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__23020\,
            I => \N__22998\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__22993\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__23014\,
            I => \N__22993\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__23009\,
            I => \N__22986\
        );

    \I__4297\ : Span4Mux_h
    port map (
            O => \N__23006\,
            I => \N__22986\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__23001\,
            I => \N__22986\
        );

    \I__4295\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22983\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__22993\,
            I => \N__22980\
        );

    \I__4293\ : Sp12to4
    port map (
            O => \N__22986\,
            I => \N__22975\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__22983\,
            I => \N__22975\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__22980\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4290\ : Odrv12
    port map (
            O => \N__22975\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4289\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22966\
        );

    \I__4288\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22963\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22960\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__22963\,
            I => \N__22957\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__22960\,
            I => \N__22954\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__22957\,
            I => \POWERLED.dutycycle_RNI_11Z0Z_7\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__22954\,
            I => \POWERLED.dutycycle_RNI_11Z0Z_7\
        );

    \I__4282\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22946\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__22946\,
            I => \POWERLED.un1_dutycycle_53_50_a0_1\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__22943\,
            I => \POWERLED.un1_dutycycle_53_2_1_cascade_\
        );

    \I__4279\ : InMux
    port map (
            O => \N__22940\,
            I => \N__22934\
        );

    \I__4278\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22934\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__4276\ : Span4Mux_h
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__4275\ : Odrv4
    port map (
            O => \N__22928\,
            I => \POWERLED.dutycycle_RNIZ0Z_8\
        );

    \I__4274\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22919\
        );

    \I__4273\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22919\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__22919\,
            I => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\
        );

    \I__4271\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22910\
        );

    \I__4270\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22910\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__22910\,
            I => \POWERLED.dutycycleZ1Z_11\
        );

    \I__4268\ : SRMux
    port map (
            O => \N__22907\,
            I => \N__22897\
        );

    \I__4267\ : SRMux
    port map (
            O => \N__22906\,
            I => \N__22894\
        );

    \I__4266\ : SRMux
    port map (
            O => \N__22905\,
            I => \N__22891\
        );

    \I__4265\ : SRMux
    port map (
            O => \N__22904\,
            I => \N__22888\
        );

    \I__4264\ : SRMux
    port map (
            O => \N__22903\,
            I => \N__22885\
        );

    \I__4263\ : SRMux
    port map (
            O => \N__22902\,
            I => \N__22881\
        );

    \I__4262\ : SRMux
    port map (
            O => \N__22901\,
            I => \N__22875\
        );

    \I__4261\ : SRMux
    port map (
            O => \N__22900\,
            I => \N__22872\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22869\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22865\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__22891\,
            I => \N__22862\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__22888\,
            I => \N__22859\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__22885\,
            I => \N__22856\
        );

    \I__4255\ : SRMux
    port map (
            O => \N__22884\,
            I => \N__22853\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__22881\,
            I => \N__22850\
        );

    \I__4253\ : SRMux
    port map (
            O => \N__22880\,
            I => \N__22847\
        );

    \I__4252\ : SRMux
    port map (
            O => \N__22879\,
            I => \N__22844\
        );

    \I__4251\ : SRMux
    port map (
            O => \N__22878\,
            I => \N__22841\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__22875\,
            I => \N__22838\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__22872\,
            I => \N__22835\
        );

    \I__4248\ : Span4Mux_s2_v
    port map (
            O => \N__22869\,
            I => \N__22832\
        );

    \I__4247\ : SRMux
    port map (
            O => \N__22868\,
            I => \N__22829\
        );

    \I__4246\ : Span4Mux_h
    port map (
            O => \N__22865\,
            I => \N__22824\
        );

    \I__4245\ : Span4Mux_h
    port map (
            O => \N__22862\,
            I => \N__22824\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__22859\,
            I => \N__22821\
        );

    \I__4243\ : Span4Mux_h
    port map (
            O => \N__22856\,
            I => \N__22818\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__22853\,
            I => \N__22813\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__22850\,
            I => \N__22813\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__22847\,
            I => \N__22810\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__22844\,
            I => \N__22807\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__22841\,
            I => \N__22804\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__22838\,
            I => \N__22801\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__22835\,
            I => \N__22798\
        );

    \I__4235\ : Sp12to4
    port map (
            O => \N__22832\,
            I => \N__22793\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__22829\,
            I => \N__22793\
        );

    \I__4233\ : Span4Mux_h
    port map (
            O => \N__22824\,
            I => \N__22790\
        );

    \I__4232\ : Span4Mux_h
    port map (
            O => \N__22821\,
            I => \N__22783\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__22818\,
            I => \N__22783\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__22813\,
            I => \N__22783\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__22810\,
            I => \N__22778\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__22807\,
            I => \N__22778\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__22804\,
            I => \N__22775\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__22801\,
            I => \N__22770\
        );

    \I__4225\ : Span4Mux_h
    port map (
            O => \N__22798\,
            I => \N__22770\
        );

    \I__4224\ : Span12Mux_s10_v
    port map (
            O => \N__22793\,
            I => \N__22767\
        );

    \I__4223\ : Span4Mux_v
    port map (
            O => \N__22790\,
            I => \N__22764\
        );

    \I__4222\ : Sp12to4
    port map (
            O => \N__22783\,
            I => \N__22761\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__22778\,
            I => \N__22758\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__22775\,
            I => \POWERLED.N_209_iZ0\
        );

    \I__4219\ : Odrv4
    port map (
            O => \N__22770\,
            I => \POWERLED.N_209_iZ0\
        );

    \I__4218\ : Odrv12
    port map (
            O => \N__22767\,
            I => \POWERLED.N_209_iZ0\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__22764\,
            I => \POWERLED.N_209_iZ0\
        );

    \I__4216\ : Odrv12
    port map (
            O => \N__22761\,
            I => \POWERLED.N_209_iZ0\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__22758\,
            I => \POWERLED.N_209_iZ0\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__22745\,
            I => \N__22742\
        );

    \I__4213\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22738\
        );

    \I__4212\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22735\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__22738\,
            I => \POWERLED.un1_dutycycle_53_31_a7_0\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__22735\,
            I => \POWERLED.un1_dutycycle_53_31_a7_0\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__22730\,
            I => \POWERLED.N_144_N_cascade_\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__22727\,
            I => \N__22724\
        );

    \I__4207\ : InMux
    port map (
            O => \N__22724\,
            I => \N__22721\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__22721\,
            I => \N__22717\
        );

    \I__4205\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22714\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__22717\,
            I => \POWERLED.dutycycle_en_7\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__22714\,
            I => \POWERLED.dutycycle_en_7\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \N__22705\
        );

    \I__4201\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22701\
        );

    \I__4200\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22696\
        );

    \I__4199\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22696\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__22701\,
            I => \N__22691\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__22696\,
            I => \N__22691\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__22691\,
            I => \POWERLED.dutycycle_eena_3_0_1\
        );

    \I__4195\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22679\
        );

    \I__4194\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22679\
        );

    \I__4193\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22679\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__22676\,
            I => \POWERLED.dutycycle_eena_3_d_0\
        );

    \I__4190\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22669\
        );

    \I__4189\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22666\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__22669\,
            I => \N__22663\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__22666\,
            I => \N__22660\
        );

    \I__4186\ : Span4Mux_s1_v
    port map (
            O => \N__22663\,
            I => \N__22655\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__22660\,
            I => \N__22655\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__22655\,
            I => \POWERLED.dutycycle_en_3\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__22652\,
            I => \POWERLED.un1_dutycycle_53_10_1_0_1_cascade_\
        );

    \I__4182\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__4180\ : Odrv12
    port map (
            O => \N__22643\,
            I => \POWERLED.un1_dutycycle_53_10_1_0\
        );

    \I__4179\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__22637\,
            I => \N__22634\
        );

    \I__4177\ : Odrv12
    port map (
            O => \N__22634\,
            I => \POWERLED.un2_count_clk_17_0_a2_4\
        );

    \I__4176\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22625\
        );

    \I__4175\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22625\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__22625\,
            I => \N__22622\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__22622\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \N__22615\
        );

    \I__4171\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22610\
        );

    \I__4170\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22610\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__22610\,
            I => \POWERLED.dutycycle_RNI4VJH7Z0Z_4\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__22607\,
            I => \N__22604\
        );

    \I__4167\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22598\
        );

    \I__4166\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22598\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__22598\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__4164\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22591\
        );

    \I__4163\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22588\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__22591\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__22588\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__22583\,
            I => \N__22579\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__22582\,
            I => \N__22576\
        );

    \I__4158\ : InMux
    port map (
            O => \N__22579\,
            I => \N__22573\
        );

    \I__4157\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22570\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__22573\,
            I => \N__22567\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__22570\,
            I => \POWERLED.dutycycleZ1Z_3\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__22567\,
            I => \POWERLED.dutycycleZ1Z_3\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__22562\,
            I => \POWERLED.dutycycleZ0Z_8_cascade_\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__22559\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_\
        );

    \I__4151\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22550\
        );

    \I__4150\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22550\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__22550\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_0\
        );

    \I__4148\ : InMux
    port map (
            O => \N__22547\,
            I => \N__22544\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__22544\,
            I => \N__22540\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__22543\,
            I => \N__22537\
        );

    \I__4145\ : Span4Mux_h
    port map (
            O => \N__22540\,
            I => \N__22534\
        );

    \I__4144\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22531\
        );

    \I__4143\ : Span4Mux_s3_h
    port map (
            O => \N__22534\,
            I => \N__22528\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22525\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__22528\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_3\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__22525\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_3\
        );

    \I__4139\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22514\
        );

    \I__4138\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22514\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__22514\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_3\
        );

    \I__4136\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__22508\,
            I => \POWERLED.un1_dutycycle_53_13_2\
        );

    \I__4134\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__22502\,
            I => \POWERLED.un1_dutycycle_53_31_4_1\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22493\
        );

    \I__4131\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22493\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__22493\,
            I => \POWERLED.dutycycle_en_8\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__22490\,
            I => \N__22486\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22481\
        );

    \I__4127\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22476\
        );

    \I__4126\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22476\
        );

    \I__4125\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22469\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__22481\,
            I => \N__22466\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__22476\,
            I => \N__22461\
        );

    \I__4122\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22456\
        );

    \I__4121\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22456\
        );

    \I__4120\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22451\
        );

    \I__4119\ : InMux
    port map (
            O => \N__22472\,
            I => \N__22451\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__22469\,
            I => \N__22448\
        );

    \I__4117\ : Span4Mux_v
    port map (
            O => \N__22466\,
            I => \N__22445\
        );

    \I__4116\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22440\
        );

    \I__4115\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22440\
        );

    \I__4114\ : Span4Mux_h
    port map (
            O => \N__22461\,
            I => \N__22437\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__22456\,
            I => \N__22432\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__22451\,
            I => \N__22432\
        );

    \I__4111\ : Span4Mux_v
    port map (
            O => \N__22448\,
            I => \N__22429\
        );

    \I__4110\ : Sp12to4
    port map (
            O => \N__22445\,
            I => \N__22424\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__22440\,
            I => \N__22424\
        );

    \I__4108\ : Sp12to4
    port map (
            O => \N__22437\,
            I => \N__22419\
        );

    \I__4107\ : Span12Mux_s10_h
    port map (
            O => \N__22432\,
            I => \N__22419\
        );

    \I__4106\ : Span4Mux_h
    port map (
            O => \N__22429\,
            I => \N__22416\
        );

    \I__4105\ : Span12Mux_s10_h
    port map (
            O => \N__22424\,
            I => \N__22413\
        );

    \I__4104\ : Odrv12
    port map (
            O => \N__22419\,
            I => slp_s3n
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__22416\,
            I => slp_s3n
        );

    \I__4102\ : Odrv12
    port map (
            O => \N__22413\,
            I => slp_s3n
        );

    \I__4101\ : IoInMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__4099\ : IoSpan4Mux
    port map (
            O => \N__22400\,
            I => \N__22396\
        );

    \I__4098\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22393\
        );

    \I__4097\ : Span4Mux_s0_v
    port map (
            O => \N__22396\,
            I => \N__22388\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22381\
        );

    \I__4095\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22376\
        );

    \I__4094\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22376\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__22388\,
            I => \N__22373\
        );

    \I__4092\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22370\
        );

    \I__4091\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22367\
        );

    \I__4090\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22362\
        );

    \I__4089\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22362\
        );

    \I__4088\ : Span4Mux_v
    port map (
            O => \N__22381\,
            I => \N__22359\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__22376\,
            I => \N__22356\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__22373\,
            I => \N__22351\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22351\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22346\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__22362\,
            I => \N__22346\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__22359\,
            I => \N__22341\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__22356\,
            I => \N__22341\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__22351\,
            I => rsmrstn
        );

    \I__4079\ : Odrv12
    port map (
            O => \N__22346\,
            I => rsmrstn
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__22341\,
            I => rsmrstn
        );

    \I__4077\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__22331\,
            I => \POWERLED.N_222\
        );

    \I__4075\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__22325\,
            I => \POWERLED.un1_dutycycle_172_sm3\
        );

    \I__4073\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__22319\,
            I => \POWERLED.un1_clk_100khz_52_and_i_m2_1\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \POWERLED.un1_dutycycle_172_m4_cascade_\
        );

    \I__4070\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__4068\ : Odrv12
    port map (
            O => \N__22307\,
            I => \POWERLED.un1_clk_100khz_52_and_i_0Z0Z_0\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__22304\,
            I => \POWERLED.N_225_cascade_\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__22301\,
            I => \POWERLED.dutycycle_eena_14_cascade_\
        );

    \I__4065\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__22289\,
            I => \POWERLED.dutycycle_eena_14\
        );

    \I__4061\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22280\
        );

    \I__4060\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22280\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__4058\ : Span4Mux_v
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__22274\,
            I => \POWERLED.dutycycle_set_1\
        );

    \I__4056\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22265\
        );

    \I__4055\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22265\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__22265\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__4053\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__22259\,
            I => \POWERLED.count_clk_0_3\
        );

    \I__4051\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__22253\,
            I => \POWERLED.count_clk_0_4\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__22250\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__22247\,
            I => \N__22239\
        );

    \I__4047\ : InMux
    port map (
            O => \N__22246\,
            I => \N__22234\
        );

    \I__4046\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22234\
        );

    \I__4045\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22231\
        );

    \I__4044\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22223\
        );

    \I__4043\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22223\
        );

    \I__4042\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22223\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__22234\,
            I => \N__22216\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22216\
        );

    \I__4039\ : InMux
    port map (
            O => \N__22230\,
            I => \N__22213\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__22223\,
            I => \N__22210\
        );

    \I__4037\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22207\
        );

    \I__4036\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22204\
        );

    \I__4035\ : Span4Mux_v
    port map (
            O => \N__22216\,
            I => \N__22201\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__22213\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__22210\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__22207\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__22204\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__22201\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4029\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22180\
        );

    \I__4026\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22177\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__22180\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_0\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__22177\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_0\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__22172\,
            I => \N__22166\
        );

    \I__4022\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22161\
        );

    \I__4021\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22161\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__22169\,
            I => \N__22158\
        );

    \I__4019\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22155\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__22161\,
            I => \N__22152\
        );

    \I__4017\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22149\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__22155\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_0\
        );

    \I__4015\ : Odrv12
    port map (
            O => \N__22152\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_0\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__22149\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_0\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__22142\,
            I => \N__22137\
        );

    \I__4012\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22133\
        );

    \I__4011\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22128\
        );

    \I__4010\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22123\
        );

    \I__4009\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22123\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__22133\,
            I => \N__22119\
        );

    \I__4007\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22114\
        );

    \I__4006\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22114\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22111\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__22123\,
            I => \N__22108\
        );

    \I__4003\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22105\
        );

    \I__4002\ : Span4Mux_v
    port map (
            O => \N__22119\,
            I => \N__22100\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__22114\,
            I => \N__22100\
        );

    \I__4000\ : Span4Mux_h
    port map (
            O => \N__22111\,
            I => \N__22097\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__22108\,
            I => \N__22092\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__22105\,
            I => \N__22092\
        );

    \I__3997\ : Span4Mux_v
    port map (
            O => \N__22100\,
            I => \N__22089\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__22097\,
            I => \N__22086\
        );

    \I__3995\ : Span4Mux_v
    port map (
            O => \N__22092\,
            I => \N__22083\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__22089\,
            I => \POWERLED.N_337\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__22086\,
            I => \POWERLED.N_337\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__22083\,
            I => \POWERLED.N_337\
        );

    \I__3991\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22073\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22069\
        );

    \I__3989\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22065\
        );

    \I__3988\ : Span4Mux_h
    port map (
            O => \N__22069\,
            I => \N__22062\
        );

    \I__3987\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22059\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__22065\,
            I => \SUSWARN_N_fast\
        );

    \I__3985\ : Odrv4
    port map (
            O => \N__22062\,
            I => \SUSWARN_N_fast\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__22059\,
            I => \SUSWARN_N_fast\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__22052\,
            I => \POWERLED.N_390_cascade_\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__22049\,
            I => \N__22045\
        );

    \I__3981\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22042\
        );

    \I__3980\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22037\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__22042\,
            I => \N__22034\
        );

    \I__3978\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22031\
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__22040\,
            I => \N__22026\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__22037\,
            I => \N__22023\
        );

    \I__3975\ : Sp12to4
    port map (
            O => \N__22034\,
            I => \N__22018\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__22031\,
            I => \N__22018\
        );

    \I__3973\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22015\
        );

    \I__3972\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22010\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22010\
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__22023\,
            I => \SUSWARN_N_rep1\
        );

    \I__3969\ : Odrv12
    port map (
            O => \N__22018\,
            I => \SUSWARN_N_rep1\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__22015\,
            I => \SUSWARN_N_rep1\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__22010\,
            I => \SUSWARN_N_rep1\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__22001\,
            I => \POWERLED.dutycycle_eena_3_0_0_sx_cascade_\
        );

    \I__3965\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__21995\,
            I => \N__21991\
        );

    \I__3963\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21987\
        );

    \I__3962\ : Span4Mux_v
    port map (
            O => \N__21991\,
            I => \N__21984\
        );

    \I__3961\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21981\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21978\
        );

    \I__3959\ : Span4Mux_h
    port map (
            O => \N__21984\,
            I => \N__21973\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__21981\,
            I => \N__21973\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__21978\,
            I => \N__21970\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__21973\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__21970\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__3953\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21956\
        );

    \I__3952\ : InMux
    port map (
            O => \N__21961\,
            I => \N__21956\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__21953\,
            I => \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7\
        );

    \I__3949\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__21947\,
            I => \POWERLED.count_0_12\
        );

    \I__3947\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__21941\,
            I => \POWERLED.count_clk_0_2\
        );

    \I__3945\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__21935\,
            I => \POWERLED.count_clk_0_13\
        );

    \I__3943\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__21926\,
            I => \POWERLED.count_clk_0_14\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__21923\,
            I => \POWERLED.un1_clk_100khz_48_and_i_o2_2_0_cascade_\
        );

    \I__3939\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__21917\,
            I => \POWERLED.un1_clk_100khz_48_and_i_o2_3_0\
        );

    \I__3937\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21910\
        );

    \I__3936\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21907\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__21910\,
            I => \POWERLED.N_197\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__21907\,
            I => \POWERLED.N_197\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__21902\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\
        );

    \I__3932\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__3930\ : Span4Mux_h
    port map (
            O => \N__21893\,
            I => \N__21888\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__21892\,
            I => \N__21885\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__21891\,
            I => \N__21882\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__21888\,
            I => \N__21877\
        );

    \I__3926\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21874\
        );

    \I__3925\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21871\
        );

    \I__3924\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21868\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21865\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__21877\,
            I => \N__21862\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__21874\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__21871\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__21868\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__21865\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__21862\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__21851\,
            I => \N__21848\
        );

    \I__3915\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__3913\ : Span4Mux_v
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__3912\ : Span4Mux_h
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__21836\,
            I => \POWERLED.un85_clk_100khz_10\
        );

    \I__3910\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__21830\,
            I => \POWERLED.un1_func_state25_6_0_o_N_287_N\
        );

    \I__3908\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__21824\,
            I => \POWERLED.func_state_RNI_1Z0Z_0\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__21821\,
            I => \POWERLED.func_state_RNI_1Z0Z_0_cascade_\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__3904\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N__21807\
        );

    \I__3902\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21804\
        );

    \I__3901\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21801\
        );

    \I__3900\ : Odrv12
    port map (
            O => \N__21807\,
            I => \POWERLED.func_state_RNIBK1UZ0Z_0\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__21804\,
            I => \POWERLED.func_state_RNIBK1UZ0Z_0\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__21801\,
            I => \POWERLED.func_state_RNIBK1UZ0Z_0\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__21794\,
            I => \N__21790\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__21793\,
            I => \N__21787\
        );

    \I__3895\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21783\
        );

    \I__3894\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21780\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__21786\,
            I => \N__21777\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__21783\,
            I => \N__21772\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__21780\,
            I => \N__21769\
        );

    \I__3890\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21764\
        );

    \I__3889\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21764\
        );

    \I__3888\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21760\
        );

    \I__3887\ : Span4Mux_v
    port map (
            O => \N__21772\,
            I => \N__21755\
        );

    \I__3886\ : Span4Mux_v
    port map (
            O => \N__21769\,
            I => \N__21755\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__21764\,
            I => \N__21752\
        );

    \I__3884\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21748\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__21760\,
            I => \N__21745\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__21755\,
            I => \N__21740\
        );

    \I__3881\ : Span4Mux_v
    port map (
            O => \N__21752\,
            I => \N__21740\
        );

    \I__3880\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21737\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__21748\,
            I => \POWERLED.N_326_0\
        );

    \I__3878\ : Odrv12
    port map (
            O => \N__21745\,
            I => \POWERLED.N_326_0\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__21740\,
            I => \POWERLED.N_326_0\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__21737\,
            I => \POWERLED.N_326_0\
        );

    \I__3875\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__21722\,
            I => \N__21718\
        );

    \I__3872\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21715\
        );

    \I__3871\ : Span4Mux_h
    port map (
            O => \N__21718\,
            I => \N__21712\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__21715\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__21712\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__3868\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21704\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__3864\ : Span4Mux_h
    port map (
            O => \N__21695\,
            I => \N__21691\
        );

    \I__3863\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21688\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__21691\,
            I => \POWERLED.func_state_RNIB74H7Z0Z_1\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__21688\,
            I => \POWERLED.func_state_RNIB74H7Z0Z_1\
        );

    \I__3860\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__3858\ : Odrv12
    port map (
            O => \N__21677\,
            I => \POWERLED.func_state_RNI6RANZ0Z_1\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__21674\,
            I => \POWERLED.func_stateZ0Z_0_cascade_\
        );

    \I__3856\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__3854\ : Span4Mux_v
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__21662\,
            I => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__21659\,
            I => \POWERLED.N_275_cascade_\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__21656\,
            I => \POWERLED.count_off_RNIZ0Z_11_cascade_\
        );

    \I__3850\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__21650\,
            I => \POWERLED.N_310\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__21647\,
            I => \POWERLED.N_314_cascade_\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__3846\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21636\
        );

    \I__3845\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21631\
        );

    \I__3844\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21631\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__21636\,
            I => \N__21624\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__21631\,
            I => \N__21624\
        );

    \I__3841\ : InMux
    port map (
            O => \N__21630\,
            I => \N__21621\
        );

    \I__3840\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21618\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__21624\,
            I => \POWERLED.count_off_RNIZ0Z_11\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__21621\,
            I => \POWERLED.count_off_RNIZ0Z_11\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__21618\,
            I => \POWERLED.count_off_RNIZ0Z_11\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__21611\,
            I => \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_\
        );

    \I__3835\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21605\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__21605\,
            I => \POWERLED.func_state_RNIHDGK3_0Z0Z_1\
        );

    \I__3833\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21595\
        );

    \I__3831\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21592\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__21595\,
            I => \POWERLED.N_67\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__21592\,
            I => \POWERLED.N_67\
        );

    \I__3828\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__21584\,
            I => \POWERLED.func_state_1_m0_0\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__21581\,
            I => \POWERLED.func_state_RNIHDGK3_0Z0Z_1_cascade_\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__21578\,
            I => \N__21566\
        );

    \I__3824\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21548\
        );

    \I__3823\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21548\
        );

    \I__3822\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21548\
        );

    \I__3821\ : InMux
    port map (
            O => \N__21574\,
            I => \N__21548\
        );

    \I__3820\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21548\
        );

    \I__3819\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21548\
        );

    \I__3818\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21548\
        );

    \I__3817\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21537\
        );

    \I__3816\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21537\
        );

    \I__3815\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21537\
        );

    \I__3814\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21537\
        );

    \I__3813\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21537\
        );

    \I__3812\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21534\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__21548\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__21537\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__21534\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__21527\,
            I => \N__21519\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \N__21515\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__21525\,
            I => \N__21512\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__21524\,
            I => \N__21509\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__21523\,
            I => \N__21500\
        );

    \I__3803\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21496\
        );

    \I__3802\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21493\
        );

    \I__3801\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21480\
        );

    \I__3800\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21480\
        );

    \I__3799\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21480\
        );

    \I__3798\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21480\
        );

    \I__3797\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21480\
        );

    \I__3796\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21480\
        );

    \I__3795\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21473\
        );

    \I__3794\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21473\
        );

    \I__3793\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21473\
        );

    \I__3792\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21466\
        );

    \I__3791\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21466\
        );

    \I__3790\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21466\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21463\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__21493\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__21480\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__21473\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__21466\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__21463\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3783\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21428\
        );

    \I__3782\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21428\
        );

    \I__3781\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21428\
        );

    \I__3780\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21428\
        );

    \I__3779\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21428\
        );

    \I__3778\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21428\
        );

    \I__3777\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21428\
        );

    \I__3776\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21421\
        );

    \I__3775\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21421\
        );

    \I__3774\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21421\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__21428\,
            I => \HDA_STRAP.un4_count\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__21421\,
            I => \HDA_STRAP.un4_count\
        );

    \I__3771\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__21413\,
            I => \POWERLED.func_state_1_m2s2_i_0\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__21410\,
            I => \POWERLED.func_state_1_m2s2_i_1_cascade_\
        );

    \I__3768\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21404\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__3766\ : Span4Mux_s3_v
    port map (
            O => \N__21401\,
            I => \N__21398\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__21398\,
            I => \POWERLED.func_state_1_m0_0_1_0\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__21395\,
            I => \HDA_STRAP.un4_count_9_cascade_\
        );

    \I__3763\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__21389\,
            I => \HDA_STRAP.un4_count_13\
        );

    \I__3761\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21383\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__21383\,
            I => \HDA_STRAP.un4_count_11\
        );

    \I__3759\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21377\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__21377\,
            I => \HDA_STRAP.un4_count_10\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__21374\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_0_0_cascade_\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__3755\ : InMux
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__21365\,
            I => \POWERLED.dutycycle_RNIEB706Z0Z_7\
        );

    \I__3753\ : InMux
    port map (
            O => \N__21362\,
            I => \N__21356\
        );

    \I__3752\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21356\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__21356\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__21353\,
            I => \POWERLED.dutycycle_RNIEB706Z0Z_7_cascade_\
        );

    \I__3749\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21344\
        );

    \I__3748\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21344\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__21341\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__21338\,
            I => \POWERLED.dutycycleZ1Z_6_cascade_\
        );

    \I__3744\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__21332\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_d_0\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__21329\,
            I => \POWERLED.N_143_N_cascade_\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__21326\,
            I => \N__21322\
        );

    \I__3740\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21317\
        );

    \I__3739\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21317\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__21317\,
            I => \N__21314\
        );

    \I__3737\ : Span4Mux_h
    port map (
            O => \N__21314\,
            I => \N__21311\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__21311\,
            I => \POWERLED.dutycycle_en_4\
        );

    \I__3735\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21301\
        );

    \I__3733\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21298\
        );

    \I__3732\ : Span4Mux_s1_v
    port map (
            O => \N__21301\,
            I => \N__21293\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21293\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__21293\,
            I => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \N__21287\
        );

    \I__3728\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21283\
        );

    \I__3727\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21280\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__21283\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__21280\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__3723\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21269\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__21269\,
            I => \HDA_STRAP.un4_count_12\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__21266\,
            I => \POWERLED.g0_i_1_cascade_\
        );

    \I__3720\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__21260\,
            I => \POWERLED.g0_i_0\
        );

    \I__3718\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__3716\ : Span4Mux_v
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__21248\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_13\
        );

    \I__3714\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21239\
        );

    \I__3713\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21239\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__21236\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__21233\,
            I => \N__21229\
        );

    \I__3709\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21224\
        );

    \I__3708\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21224\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__21224\,
            I => \POWERLED.dutycycle_rst_1\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__21221\,
            I => \POWERLED.dutycycleZ0Z_4_cascade_\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__21218\,
            I => \POWERLED.g0_1_cascade_\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__3703\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21206\
        );

    \I__3702\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21206\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__21206\,
            I => \N__21201\
        );

    \I__3700\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21196\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__21204\,
            I => \N__21193\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__21201\,
            I => \N__21190\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__21200\,
            I => \N__21186\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__21199\,
            I => \N__21183\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21179\
        );

    \I__3694\ : InMux
    port map (
            O => \N__21193\,
            I => \N__21176\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__21190\,
            I => \N__21173\
        );

    \I__3692\ : InMux
    port map (
            O => \N__21189\,
            I => \N__21168\
        );

    \I__3691\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21168\
        );

    \I__3690\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21163\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21163\
        );

    \I__3688\ : Span4Mux_s3_v
    port map (
            O => \N__21179\,
            I => \N__21158\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__21176\,
            I => \N__21158\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__21173\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__21168\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__21163\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__21158\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__21149\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__3680\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__3678\ : Span4Mux_h
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__21134\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_14\
        );

    \I__3676\ : InMux
    port map (
            O => \N__21131\,
            I => \POWERLED.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__3675\ : InMux
    port map (
            O => \N__21128\,
            I => \bfn_7_13_0_\
        );

    \I__3674\ : InMux
    port map (
            O => \N__21125\,
            I => \POWERLED.un1_dutycycle_94_cry_8_cZ0\
        );

    \I__3673\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21116\
        );

    \I__3672\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21116\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__21116\,
            I => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\
        );

    \I__3670\ : InMux
    port map (
            O => \N__21113\,
            I => \POWERLED.un1_dutycycle_94_cry_9\
        );

    \I__3669\ : InMux
    port map (
            O => \N__21110\,
            I => \POWERLED.un1_dutycycle_94_cry_10\
        );

    \I__3668\ : InMux
    port map (
            O => \N__21107\,
            I => \POWERLED.un1_dutycycle_94_cry_11\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21098\
        );

    \I__3666\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21098\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__21098\,
            I => \N__21095\
        );

    \I__3664\ : Odrv12
    port map (
            O => \N__21095\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\
        );

    \I__3663\ : InMux
    port map (
            O => \N__21092\,
            I => \POWERLED.un1_dutycycle_94_cry_12\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__21089\,
            I => \N__21085\
        );

    \I__3661\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21080\
        );

    \I__3660\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21080\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__21077\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\
        );

    \I__3657\ : InMux
    port map (
            O => \N__21074\,
            I => \POWERLED.un1_dutycycle_94_cry_13\
        );

    \I__3656\ : InMux
    port map (
            O => \N__21071\,
            I => \POWERLED.un1_dutycycle_94_cry_14\
        );

    \I__3655\ : InMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__21065\,
            I => \N__21062\
        );

    \I__3653\ : Span4Mux_h
    port map (
            O => \N__21062\,
            I => \N__21058\
        );

    \I__3652\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21055\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__21058\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__21055\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\
        );

    \I__3649\ : CascadeMux
    port map (
            O => \N__21050\,
            I => \POWERLED.un1_dutycycle_53_13_4_cascade_\
        );

    \I__3648\ : InMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__3646\ : Span4Mux_v
    port map (
            O => \N__21041\,
            I => \N__21038\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__21038\,
            I => \POWERLED.un1_dutycycle_53_13_3\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__21035\,
            I => \N__21032\
        );

    \I__3643\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__3641\ : Span4Mux_h
    port map (
            O => \N__21026\,
            I => \N__21023\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__21023\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_11\
        );

    \I__3639\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21014\
        );

    \I__3638\ : InMux
    port map (
            O => \N__21019\,
            I => \N__21014\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__21014\,
            I => \POWERLED.g0_0_1\
        );

    \I__3636\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__3634\ : Odrv12
    port map (
            O => \N__21005\,
            I => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\
        );

    \I__3633\ : InMux
    port map (
            O => \N__21002\,
            I => \POWERLED.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__3632\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20996\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__3630\ : Odrv12
    port map (
            O => \N__20993\,
            I => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\
        );

    \I__3629\ : InMux
    port map (
            O => \N__20990\,
            I => \POWERLED.un1_dutycycle_94_cry_1\
        );

    \I__3628\ : InMux
    port map (
            O => \N__20987\,
            I => \POWERLED.un1_dutycycle_94_cry_2_cZ0\
        );

    \I__3627\ : InMux
    port map (
            O => \N__20984\,
            I => \POWERLED.un1_dutycycle_94_cry_3_cZ0\
        );

    \I__3626\ : InMux
    port map (
            O => \N__20981\,
            I => \POWERLED.un1_dutycycle_94_cry_4_cZ0\
        );

    \I__3625\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__20972\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\
        );

    \I__3622\ : InMux
    port map (
            O => \N__20969\,
            I => \POWERLED.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__20966\,
            I => \POWERLED.d_i3_mux_cascade_\
        );

    \I__3620\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__20960\,
            I => \N__20957\
        );

    \I__3618\ : Span4Mux_h
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__20954\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_5\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__20951\,
            I => \N__20948\
        );

    \I__3615\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__3613\ : Odrv12
    port map (
            O => \N__20942\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_0\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__20939\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__20936\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_9_cascade_\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__20933\,
            I => \N__20930\
        );

    \I__3609\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__20924\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_7\
        );

    \I__3606\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__20918\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__3604\ : InMux
    port map (
            O => \N__20915\,
            I => \N__20912\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__20909\,
            I => \POWERLED.dutycycle_RNIZ0Z_5\
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__3600\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__3598\ : Span4Mux_v
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__20894\,
            I => \POWERLED.un1_dutycycle_53_13_4_1\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__20891\,
            I => \POWERLED.func_state_RNIBVNS_1Z0Z_0_cascade_\
        );

    \I__3595\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__20885\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_ns_1\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__20882\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\
        );

    \I__3592\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20873\
        );

    \I__3591\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20873\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__20873\,
            I => \POWERLED.N_171\
        );

    \I__3589\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__20867\,
            I => \POWERLED.N_283\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__3586\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__20855\,
            I => \N__20852\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__20852\,
            I => \POWERLED.N_275_0\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__3581\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__20843\,
            I => \POWERLED.dutycycle_set_0_0\
        );

    \I__3579\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20834\
        );

    \I__3578\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20834\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__20834\,
            I => \POWERLED.dutycycle_eena_13_0\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__20831\,
            I => \POWERLED.dutycycle_set_0_0_cascade_\
        );

    \I__3575\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20822\
        );

    \I__3574\ : InMux
    port map (
            O => \N__20827\,
            I => \N__20822\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__20822\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__20819\,
            I => \POWERLED.dutycycleZ0Z_6_cascade_\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__3570\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__3568\ : Sp12to4
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__3567\ : Span12Mux_s9_v
    port map (
            O => \N__20804\,
            I => \N__20800\
        );

    \I__3566\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20797\
        );

    \I__3565\ : Odrv12
    port map (
            O => \N__20800\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_0\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__20797\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_0\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__20792\,
            I => \POWERLED.dutycycle_en_10_cascade_\
        );

    \I__3562\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20783\
        );

    \I__3561\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20783\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__20783\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3559\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__20774\,
            I => \POWERLED.un1_func_state25_4_i_a2_1\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__20771\,
            I => \POWERLED.N_301_cascade_\
        );

    \I__3555\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__3553\ : Span4Mux_v
    port map (
            O => \N__20762\,
            I => \N__20758\
        );

    \I__3552\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20755\
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__20758\,
            I => \POWERLED.N_341\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__20755\,
            I => \POWERLED.N_341\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__20750\,
            I => \POWERLED.count_clk_en_1_0_cascade_\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__20747\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__20744\,
            I => \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_cascade_\
        );

    \I__3546\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__3544\ : Span4Mux_v
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__3543\ : Span4Mux_h
    port map (
            O => \N__20732\,
            I => \N__20727\
        );

    \I__3542\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20724\
        );

    \I__3541\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20721\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__20727\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__20724\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__20721\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__3536\ : InMux
    port map (
            O => \N__20711\,
            I => \N__20705\
        );

    \I__3535\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20705\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__20705\,
            I => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\
        );

    \I__3533\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__20699\,
            I => \POWERLED.count_0_5\
        );

    \I__3531\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__20693\,
            I => \N__20690\
        );

    \I__3529\ : Span4Mux_v
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__20687\,
            I => \N__20682\
        );

    \I__3527\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20679\
        );

    \I__3526\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20676\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__20682\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__20679\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__20676\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__20669\,
            I => \N__20666\
        );

    \I__3521\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20660\
        );

    \I__3520\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20660\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__20660\,
            I => \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\
        );

    \I__3518\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__20654\,
            I => \POWERLED.count_0_14\
        );

    \I__3516\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20648\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__3514\ : Span4Mux_v
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__20642\,
            I => \N__20637\
        );

    \I__3512\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20634\
        );

    \I__3511\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20631\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__20637\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__20634\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__20631\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__20624\,
            I => \N__20621\
        );

    \I__3506\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20615\
        );

    \I__3505\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20615\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__20615\,
            I => \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49\
        );

    \I__3503\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__20609\,
            I => \POWERLED.count_0_6\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__20606\,
            I => \POWERLED.dutycycleZ0Z_11_cascade_\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__20603\,
            I => \POWERLED.N_148_N_cascade_\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__3498\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20594\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__20594\,
            I => \POWERLED.dutycycle_en_10\
        );

    \I__3496\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20588\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__20588\,
            I => \POWERLED.dutycycle_1_0_0\
        );

    \I__3494\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20581\
        );

    \I__3493\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20578\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__20581\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__20578\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__20573\,
            I => \POWERLED.dutycycle_1_0_0_cascade_\
        );

    \I__3489\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20564\
        );

    \I__3488\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20564\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__20564\,
            I => \N__20561\
        );

    \I__3486\ : Span4Mux_h
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__20558\,
            I => \POWERLED.dutycycle_eena\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__3483\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__3481\ : Span4Mux_h
    port map (
            O => \N__20546\,
            I => \N__20542\
        );

    \I__3480\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20539\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__20542\,
            I => \N__20536\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__20539\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__20536\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3476\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__3474\ : Span12Mux_s6_h
    port map (
            O => \N__20525\,
            I => \N__20521\
        );

    \I__3473\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__3472\ : Odrv12
    port map (
            O => \N__20521\,
            I => \POWERLED.func_state_RNIG5G37Z0Z_1\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__20518\,
            I => \POWERLED.func_state_RNIG5G37Z0Z_1\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__20513\,
            I => \POWERLED.func_state_cascade_\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__20510\,
            I => \N__20507\
        );

    \I__3468\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20504\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20500\
        );

    \I__3466\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20497\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__20497\,
            I => \N__20491\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__20494\,
            I => \POWERLED.dutycycle_1_0_1\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__20491\,
            I => \POWERLED.dutycycle_1_0_1\
        );

    \I__3461\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__3459\ : Span4Mux_v
    port map (
            O => \N__20480\,
            I => \N__20477\
        );

    \I__3458\ : Span4Mux_h
    port map (
            O => \N__20477\,
            I => \N__20472\
        );

    \I__3457\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20469\
        );

    \I__3456\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20466\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__20472\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__20469\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__20466\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__20459\,
            I => \N__20456\
        );

    \I__3451\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20450\
        );

    \I__3450\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20450\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__20450\,
            I => \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7\
        );

    \I__3448\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__20444\,
            I => \POWERLED.count_0_13\
        );

    \I__3446\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__3444\ : Sp12to4
    port map (
            O => \N__20435\,
            I => \N__20432\
        );

    \I__3443\ : Odrv12
    port map (
            O => \N__20432\,
            I => \POWERLED.func_state_RNIMQ0FZ0Z_1\
        );

    \I__3442\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__20426\,
            I => \POWERLED.N_309\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__20423\,
            I => \POWERLED.func_state_1_m0_1_cascade_\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__20420\,
            I => \POWERLED.count_RNI_0_1_cascade_\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__20417\,
            I => \POWERLED.dutycycle_1_0_iv_i_a3_1_0_2_cascade_\
        );

    \I__3437\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20408\
        );

    \I__3436\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20408\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__20402\,
            I => \POWERLED.N_64\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__20399\,
            I => \POWERLED.g0_0_a3_1_cascade_\
        );

    \I__3431\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__3429\ : Span4Mux_v
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__20387\,
            I => \POWERLED.g0_3_1\
        );

    \I__3427\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__20381\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_2\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__20378\,
            I => \HDA_STRAP.N_14_cascade_\
        );

    \I__3424\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20369\
        );

    \I__3423\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20369\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__20369\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__3421\ : IoInMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__3419\ : IoSpan4Mux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__3418\ : Span4Mux_s2_h
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__3417\ : Span4Mux_h
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__20351\,
            I => hda_sdo_atp
        );

    \I__3415\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__3413\ : Span4Mux_h
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__20339\,
            I => gpio_fpga_soc_1
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__20336\,
            I => \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_\
        );

    \I__3410\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20327\
        );

    \I__3409\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20327\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20323\
        );

    \I__3407\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20320\
        );

    \I__3406\ : Odrv12
    port map (
            O => \N__20323\,
            I => \PCH_PWRGD_delayed_vccin_ok\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__20320\,
            I => \PCH_PWRGD_delayed_vccin_ok\
        );

    \I__3404\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__20312\,
            I => \HDA_STRAP.curr_state_RNO_0Z0Z_0\
        );

    \I__3402\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20306\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__20306\,
            I => \HDA_STRAP.N_5_0\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__20303\,
            I => \POWERLED.N_341_cascade_\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__20300\,
            I => \POWERLED.dutycycle_RNI_11Z0Z_7_cascade_\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__20297\,
            I => \N__20294\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__20288\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_12\
        );

    \I__3394\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__20282\,
            I => \POWERLED.un1_dutycycle_53_4_1\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__20279\,
            I => \POWERLED.dutycycleZ0Z_3_cascade_\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__3390\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20270\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__20270\,
            I => \POWERLED.un1_dutycycle_53_45_a0_1\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__20267\,
            I => \POWERLED.un1_dutycycle_53_45_a0_1_cascade_\
        );

    \I__3387\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20261\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__20261\,
            I => \N__20258\
        );

    \I__3385\ : Span4Mux_v
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__20255\,
            I => \POWERLED.un1_dutycycle_53_10_1\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__3382\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20246\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__20246\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__3380\ : InMux
    port map (
            O => \N__20243\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__3378\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__20234\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__3375\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__20225\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__3373\ : InMux
    port map (
            O => \N__20222\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__3372\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__20216\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__3370\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__20210\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__3368\ : InMux
    port map (
            O => \N__20207\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__3367\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20200\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__20203\,
            I => \N__20196\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__20200\,
            I => \N__20192\
        );

    \I__3364\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20187\
        );

    \I__3363\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20187\
        );

    \I__3362\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20184\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__20192\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__20187\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__20184\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__3357\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__20171\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__3355\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__20165\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__3353\ : InMux
    port map (
            O => \N__20162\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__3352\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__20156\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__20153\,
            I => \N__20149\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__20152\,
            I => \N__20145\
        );

    \I__3348\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20138\
        );

    \I__3347\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20138\
        );

    \I__3346\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20138\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__20138\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__3343\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__20129\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__3341\ : InMux
    port map (
            O => \N__20126\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__20123\,
            I => \N__20120\
        );

    \I__3339\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__20117\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__3337\ : InMux
    port map (
            O => \N__20114\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__3336\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__20108\,
            I => \N__20104\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__20107\,
            I => \N__20100\
        );

    \I__3333\ : Span4Mux_h
    port map (
            O => \N__20104\,
            I => \N__20095\
        );

    \I__3332\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20092\
        );

    \I__3331\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20085\
        );

    \I__3330\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20085\
        );

    \I__3329\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20085\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__20095\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__20092\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__20085\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3325\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__20075\,
            I => \N__20071\
        );

    \I__3323\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20068\
        );

    \I__3322\ : Span4Mux_v
    port map (
            O => \N__20071\,
            I => \N__20065\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__20068\,
            I => \N__20062\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__20065\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__3319\ : Odrv12
    port map (
            O => \N__20062\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__3318\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__20054\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__3316\ : InMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__20048\,
            I => \N__20043\
        );

    \I__3314\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20040\
        );

    \I__3313\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20037\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__20043\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__20040\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__20037\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20030\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__3307\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__3305\ : Odrv4
    port map (
            O => \N__20018\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__3304\ : InMux
    port map (
            O => \N__20015\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__3302\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20006\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__20006\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__3299\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__19994\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__3296\ : InMux
    port map (
            O => \N__19991\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__3295\ : InMux
    port map (
            O => \N__19988\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__3293\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__19979\,
            I => \POWERLED.un1_dutycycle_53_i_29\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__19976\,
            I => \N__19971\
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__19975\,
            I => \N__19967\
        );

    \I__3289\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19962\
        );

    \I__3288\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19962\
        );

    \I__3287\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19957\
        );

    \I__3286\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19957\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__19962\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__19957\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__3283\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19945\
        );

    \I__3282\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19945\
        );

    \I__3281\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19942\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__19945\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__19942\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__3277\ : InMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__19931\,
            I => \POWERLED.mult1_un47_sum_s_4_sf\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19924\
        );

    \I__3274\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19921\
        );

    \I__3273\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19918\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__19921\,
            I => \N__19915\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__19918\,
            I => \N__19912\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__19915\,
            I => \N__19909\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__19912\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__19909\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \N__19900\
        );

    \I__3266\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19897\
        );

    \I__3265\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19894\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19891\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19888\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__19891\,
            I => \N__19885\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__19888\,
            I => \POWERLED.dutycycle_en_12\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__19885\,
            I => \POWERLED.dutycycle_en_12\
        );

    \I__3259\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19876\
        );

    \I__3258\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19873\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__19876\,
            I => \N__19870\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__19873\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__19870\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__19865\,
            I => \POWERLED.un1_dutycycle_53_axb_10_1_cascade_\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__19862\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__3251\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__19853\,
            I => \POWERLED.dutycycle_RNIZ0Z_13\
        );

    \I__3249\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19844\
        );

    \I__3248\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19844\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__19844\,
            I => \POWERLED.dutycycleZ1Z_10\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__19841\,
            I => \POWERLED.dutycycleZ0Z_2_cascade_\
        );

    \I__3245\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__19835\,
            I => \POWERLED.dutycycle_RNIZ0Z_10\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__19832\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_9_cascade_\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__19829\,
            I => \N__19825\
        );

    \I__3241\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19822\
        );

    \I__3240\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19819\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__19822\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__19819\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__3237\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__19811\,
            I => \POWERLED.N_353_0\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__19808\,
            I => \POWERLED.dutycycleZ0Z_10_cascade_\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__3233\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__19796\,
            I => \POWERLED.dutycycle_RNIZ0Z_14\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__19793\,
            I => \POWERLED.N_86_f0_cascade_\
        );

    \I__3229\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__19787\,
            I => \POWERLED.dutycycle_en_11\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__19784\,
            I => \POWERLED.dutycycle_en_11_cascade_\
        );

    \I__3226\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__19778\,
            I => \N__19774\
        );

    \I__3224\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19771\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__19774\,
            I => \N__19768\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__19771\,
            I => \POWERLED.dutycycleZ1Z_14\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__19768\,
            I => \POWERLED.dutycycleZ1Z_14\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__3219\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__19757\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_15\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__19754\,
            I => \N__19750\
        );

    \I__3216\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19747\
        );

    \I__3215\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19744\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__19747\,
            I => \N__19741\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19738\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__19741\,
            I => \N__19735\
        );

    \I__3211\ : Span12Mux_s10_h
    port map (
            O => \N__19738\,
            I => \N__19732\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__19735\,
            I => \POWERLED.N_2215_i\
        );

    \I__3209\ : Odrv12
    port map (
            O => \N__19732\,
            I => \POWERLED.N_2215_i\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__19727\,
            I => \POWERLED.N_84_f0_cascade_\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__19724\,
            I => \POWERLED.N_108_f0_1_cascade_\
        );

    \I__3206\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__19718\,
            I => \POWERLED.dutycycle_eena_0\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__19715\,
            I => \POWERLED.dutycycle_eena_0_cascade_\
        );

    \I__3203\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19706\
        );

    \I__3202\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19706\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__19706\,
            I => \POWERLED.dutycycleZ1Z_1\
        );

    \I__3200\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__19700\,
            I => \POWERLED.dutycycle_eena_1\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__3197\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19690\
        );

    \I__3196\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19687\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__19690\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__19687\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__19682\,
            I => \POWERLED.func_state_0_sqmuxa_0_o2_xZ0Z1_cascade_\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__19679\,
            I => \POWERLED.g1_1_cascade_\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__19676\,
            I => \POWERLED.N_300_N_0_cascade_\
        );

    \I__3190\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__19670\,
            I => \POWERLED.N_4548_0\
        );

    \I__3188\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__19664\,
            I => \POWERLED.N_217_N_0\
        );

    \I__3186\ : InMux
    port map (
            O => \N__19661\,
            I => \POWERLED.un1_count_cry_12\
        );

    \I__3185\ : InMux
    port map (
            O => \N__19658\,
            I => \POWERLED.un1_count_cry_13\
        );

    \I__3184\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__19652\,
            I => \N__19647\
        );

    \I__3182\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19644\
        );

    \I__3181\ : InMux
    port map (
            O => \N__19650\,
            I => \N__19641\
        );

    \I__3180\ : Span4Mux_v
    port map (
            O => \N__19647\,
            I => \N__19638\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__19644\,
            I => \N__19633\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__19641\,
            I => \N__19633\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__19638\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__19633\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__3175\ : InMux
    port map (
            O => \N__19628\,
            I => \POWERLED.un1_count_cry_14\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__3173\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19616\
        );

    \I__3172\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19616\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__19616\,
            I => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\
        );

    \I__3170\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__19610\,
            I => \POWERLED.count_0_9\
        );

    \I__3168\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19603\
        );

    \I__3167\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19600\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__19603\,
            I => \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__19600\,
            I => \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79\
        );

    \I__3164\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__19592\,
            I => \N__19588\
        );

    \I__3162\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19584\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__19588\,
            I => \N__19581\
        );

    \I__3160\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19578\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__19584\,
            I => \N__19575\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__19581\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__19578\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__19575\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \POWERLED.dutycycle_eena_1_cascade_\
        );

    \I__3154\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__19562\,
            I => \POWERLED.N_108_f0_1\
        );

    \I__3152\ : InMux
    port map (
            O => \N__19559\,
            I => \POWERLED.un1_count_cry_4\
        );

    \I__3151\ : InMux
    port map (
            O => \N__19556\,
            I => \POWERLED.un1_count_cry_5\
        );

    \I__3150\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__19550\,
            I => \N__19545\
        );

    \I__3148\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19542\
        );

    \I__3147\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19539\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__19545\,
            I => \N__19532\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__19542\,
            I => \N__19532\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__19539\,
            I => \N__19532\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__19532\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__19529\,
            I => \N__19526\
        );

    \I__3141\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19520\
        );

    \I__3140\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19520\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__19520\,
            I => \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59\
        );

    \I__3138\ : InMux
    port map (
            O => \N__19517\,
            I => \POWERLED.un1_count_cry_6\
        );

    \I__3137\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19510\
        );

    \I__3136\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19507\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__19510\,
            I => \N__19503\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__19507\,
            I => \N__19500\
        );

    \I__3133\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19497\
        );

    \I__3132\ : Span4Mux_h
    port map (
            O => \N__19503\,
            I => \N__19492\
        );

    \I__3131\ : Span4Mux_h
    port map (
            O => \N__19500\,
            I => \N__19492\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__19497\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__19492\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__3127\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19478\
        );

    \I__3126\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19478\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__19478\,
            I => \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69\
        );

    \I__3124\ : InMux
    port map (
            O => \N__19475\,
            I => \POWERLED.un1_count_cry_7\
        );

    \I__3123\ : InMux
    port map (
            O => \N__19472\,
            I => \bfn_6_8_0_\
        );

    \I__3122\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19466\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__19466\,
            I => \N__19461\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__19465\,
            I => \N__19458\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__19464\,
            I => \N__19455\
        );

    \I__3118\ : Span4Mux_v
    port map (
            O => \N__19461\,
            I => \N__19452\
        );

    \I__3117\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19449\
        );

    \I__3116\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19446\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__19452\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__19449\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__19446\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__19439\,
            I => \N__19435\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__3110\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__3109\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__19429\,
            I => \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__19426\,
            I => \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\
        );

    \I__3106\ : InMux
    port map (
            O => \N__19421\,
            I => \POWERLED.un1_count_cry_9\
        );

    \I__3105\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__3103\ : Span4Mux_v
    port map (
            O => \N__19412\,
            I => \N__19407\
        );

    \I__3102\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19404\
        );

    \I__3101\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19401\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__19407\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__19404\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__19401\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__19394\,
            I => \N__19390\
        );

    \I__3096\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19385\
        );

    \I__3095\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19385\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__19385\,
            I => \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7\
        );

    \I__3093\ : InMux
    port map (
            O => \N__19382\,
            I => \POWERLED.un1_count_cry_10\
        );

    \I__3092\ : InMux
    port map (
            O => \N__19379\,
            I => \POWERLED.un1_count_cry_11\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \POWERLED.un79_clk_100khzlt15_0_cascade_\
        );

    \I__3090\ : SRMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__3088\ : Span4Mux_v
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__3087\ : Span4Mux_s2_v
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__19361\,
            I => \POWERLED.pwm_out_1_sqmuxa\
        );

    \I__3085\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__19355\,
            I => \POWERLED.un79_clk_100khzlto15_5\
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__19352\,
            I => \POWERLED.un79_clk_100khzlto15_6_cascade_\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__19349\,
            I => \POWERLED.count_RNIZ0Z_15_cascade_\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__3080\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19337\
        );

    \I__3079\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19337\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__19337\,
            I => \POWERLED.N_8\
        );

    \I__3077\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__3075\ : Span4Mux_v
    port map (
            O => \N__19328\,
            I => \N__19323\
        );

    \I__3074\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19320\
        );

    \I__3073\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19317\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__19323\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__19320\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__19317\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__3068\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19301\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19301\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__19301\,
            I => \POWERLED.un1_count_cry_1_c_RNIBZ0Z209\
        );

    \I__3065\ : InMux
    port map (
            O => \N__19298\,
            I => \POWERLED.un1_count_cry_1\
        );

    \I__3064\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__3062\ : Span4Mux_v
    port map (
            O => \N__19289\,
            I => \N__19284\
        );

    \I__3061\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19281\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19278\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__19284\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__19281\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__19278\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__3055\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19262\
        );

    \I__3054\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19262\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__19262\,
            I => \POWERLED.un1_count_cry_2_c_RNICZ0Z419\
        );

    \I__3052\ : InMux
    port map (
            O => \N__19259\,
            I => \POWERLED.un1_count_cry_2\
        );

    \I__3051\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19249\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__19252\,
            I => \N__19245\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__19249\,
            I => \N__19242\
        );

    \I__3047\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19239\
        );

    \I__3046\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19236\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__19242\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__19239\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__19236\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__3042\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__19223\,
            I => \N__19219\
        );

    \I__3039\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19216\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__19219\,
            I => \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__19216\,
            I => \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\
        );

    \I__3036\ : InMux
    port map (
            O => \N__19211\,
            I => \POWERLED.un1_count_cry_3\
        );

    \I__3035\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19204\
        );

    \I__3034\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19201\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__19204\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__19201\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__3031\ : InMux
    port map (
            O => \N__19196\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__19193\,
            I => \N__19189\
        );

    \I__3029\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19186\
        );

    \I__3028\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19183\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__19186\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__19183\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__3025\ : InMux
    port map (
            O => \N__19178\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__19175\,
            I => \N__19171\
        );

    \I__3023\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19168\
        );

    \I__3022\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19165\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__19168\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__19165\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__3019\ : InMux
    port map (
            O => \N__19160\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__3018\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19153\
        );

    \I__3017\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19150\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__19153\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__19150\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__3014\ : InMux
    port map (
            O => \N__19145\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__3013\ : InMux
    port map (
            O => \N__19142\,
            I => \bfn_6_5_0_\
        );

    \I__3012\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19135\
        );

    \I__3011\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19132\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__19135\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__19132\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__3008\ : CEMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__19118\,
            I => \RSMRST_PWRGD.N_27_2\
        );

    \I__3004\ : SRMux
    port map (
            O => \N__19115\,
            I => \N__19111\
        );

    \I__3003\ : SRMux
    port map (
            O => \N__19114\,
            I => \N__19108\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__19111\,
            I => \N__19105\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19101\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__19105\,
            I => \N__19098\
        );

    \I__2999\ : SRMux
    port map (
            O => \N__19104\,
            I => \N__19095\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__19101\,
            I => \G_11\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__19098\,
            I => \G_11\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__19095\,
            I => \G_11\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__19088\,
            I => \POWERLED.un79_clk_100khzlto4_0_cascade_\
        );

    \I__2994\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19081\
        );

    \I__2993\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__19081\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__19078\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__2990\ : InMux
    port map (
            O => \N__19073\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__19070\,
            I => \N__19066\
        );

    \I__2988\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19063\
        );

    \I__2987\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19060\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__19063\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__19060\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__2984\ : InMux
    port map (
            O => \N__19055\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__2983\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19048\
        );

    \I__2982\ : InMux
    port map (
            O => \N__19051\,
            I => \N__19045\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__19048\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__19045\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__2979\ : InMux
    port map (
            O => \N__19040\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__2978\ : InMux
    port map (
            O => \N__19037\,
            I => \N__19033\
        );

    \I__2977\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__19033\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__19030\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__2974\ : InMux
    port map (
            O => \N__19025\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__2973\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19018\
        );

    \I__2972\ : InMux
    port map (
            O => \N__19021\,
            I => \N__19015\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__19018\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__19015\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__2969\ : InMux
    port map (
            O => \N__19010\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__2968\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19003\
        );

    \I__2967\ : InMux
    port map (
            O => \N__19006\,
            I => \N__19000\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__19003\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__19000\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__2964\ : InMux
    port map (
            O => \N__18995\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__18992\,
            I => \N__18988\
        );

    \I__2962\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18985\
        );

    \I__2961\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18982\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__18985\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__18982\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__2958\ : InMux
    port map (
            O => \N__18977\,
            I => \bfn_6_4_0_\
        );

    \I__2957\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18970\
        );

    \I__2956\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18967\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__18970\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__18967\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__2953\ : InMux
    port map (
            O => \N__18962\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__2952\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18955\
        );

    \I__2951\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18952\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__18955\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__18952\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__2948\ : InMux
    port map (
            O => \N__18947\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__2947\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__18941\,
            I => \PCH_PWRGD.un2_count_1_axb_2\
        );

    \I__2945\ : SRMux
    port map (
            O => \N__18938\,
            I => \N__18932\
        );

    \I__2944\ : SRMux
    port map (
            O => \N__18937\,
            I => \N__18929\
        );

    \I__2943\ : SRMux
    port map (
            O => \N__18936\,
            I => \N__18923\
        );

    \I__2942\ : SRMux
    port map (
            O => \N__18935\,
            I => \N__18920\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18917\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__18929\,
            I => \N__18914\
        );

    \I__2939\ : SRMux
    port map (
            O => \N__18928\,
            I => \N__18910\
        );

    \I__2938\ : SRMux
    port map (
            O => \N__18927\,
            I => \N__18907\
        );

    \I__2937\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18904\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__18923\,
            I => \N__18901\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__18920\,
            I => \N__18898\
        );

    \I__2934\ : IoSpan4Mux
    port map (
            O => \N__18917\,
            I => \N__18893\
        );

    \I__2933\ : Span4Mux_v
    port map (
            O => \N__18914\,
            I => \N__18893\
        );

    \I__2932\ : SRMux
    port map (
            O => \N__18913\,
            I => \N__18890\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__18910\,
            I => \N__18883\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18883\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__18904\,
            I => \N__18883\
        );

    \I__2928\ : Span4Mux_s1_v
    port map (
            O => \N__18901\,
            I => \N__18876\
        );

    \I__2927\ : Span4Mux_h
    port map (
            O => \N__18898\,
            I => \N__18867\
        );

    \I__2926\ : Span4Mux_s1_v
    port map (
            O => \N__18893\,
            I => \N__18867\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18867\
        );

    \I__2924\ : Span4Mux_v
    port map (
            O => \N__18883\,
            I => \N__18867\
        );

    \I__2923\ : InMux
    port map (
            O => \N__18882\,
            I => \N__18860\
        );

    \I__2922\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18860\
        );

    \I__2921\ : InMux
    port map (
            O => \N__18880\,
            I => \N__18860\
        );

    \I__2920\ : SRMux
    port map (
            O => \N__18879\,
            I => \N__18857\
        );

    \I__2919\ : Sp12to4
    port map (
            O => \N__18876\,
            I => \N__18850\
        );

    \I__2918\ : Sp12to4
    port map (
            O => \N__18867\,
            I => \N__18850\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__18860\,
            I => \N__18850\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__18857\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__2915\ : Odrv12
    port map (
            O => \N__18850\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__2913\ : InMux
    port map (
            O => \N__18842\,
            I => \N__18833\
        );

    \I__2912\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18833\
        );

    \I__2911\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18833\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__18833\,
            I => \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSCZ0\
        );

    \I__2909\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18824\
        );

    \I__2908\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18824\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__18824\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__18821\,
            I => \PCH_PWRGD.count_rst_12_cascade_\
        );

    \I__2905\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__18815\,
            I => \N__18811\
        );

    \I__2903\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18808\
        );

    \I__2902\ : Span4Mux_s1_v
    port map (
            O => \N__18811\,
            I => \N__18805\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__18808\,
            I => \N__18802\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__18805\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__18802\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__2898\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__2896\ : Span4Mux_v
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__18788\,
            I => \PCH_PWRGD.un12_clk_100khz_3\
        );

    \I__2894\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__18782\,
            I => \PCH_PWRGD.count_0_12\
        );

    \I__2892\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__18776\,
            I => \N__18772\
        );

    \I__2890\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18769\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__18772\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__18769\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__2887\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__18761\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__2885\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18751\
        );

    \I__2884\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18751\
        );

    \I__2883\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18748\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__18751\,
            I => \N__18745\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__18748\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__2880\ : Odrv12
    port map (
            O => \N__18745\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__2879\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18733\
        );

    \I__2877\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18730\
        );

    \I__2876\ : Span4Mux_s1_v
    port map (
            O => \N__18733\,
            I => \N__18727\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__18730\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__18727\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__18722\,
            I => \PCH_PWRGD.countZ0Z_12_cascade_\
        );

    \I__2872\ : CEMux
    port map (
            O => \N__18719\,
            I => \N__18710\
        );

    \I__2871\ : CEMux
    port map (
            O => \N__18718\,
            I => \N__18707\
        );

    \I__2870\ : CEMux
    port map (
            O => \N__18717\,
            I => \N__18704\
        );

    \I__2869\ : CEMux
    port map (
            O => \N__18716\,
            I => \N__18698\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__18715\,
            I => \N__18694\
        );

    \I__2867\ : CEMux
    port map (
            O => \N__18714\,
            I => \N__18685\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__18713\,
            I => \N__18682\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__18710\,
            I => \N__18673\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__18707\,
            I => \N__18670\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__18704\,
            I => \N__18667\
        );

    \I__2862\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18658\
        );

    \I__2861\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18658\
        );

    \I__2860\ : CEMux
    port map (
            O => \N__18701\,
            I => \N__18655\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__18698\,
            I => \N__18652\
        );

    \I__2858\ : CEMux
    port map (
            O => \N__18697\,
            I => \N__18647\
        );

    \I__2857\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18647\
        );

    \I__2856\ : InMux
    port map (
            O => \N__18693\,
            I => \N__18642\
        );

    \I__2855\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18642\
        );

    \I__2854\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18637\
        );

    \I__2853\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18637\
        );

    \I__2852\ : InMux
    port map (
            O => \N__18689\,
            I => \N__18629\
        );

    \I__2851\ : InMux
    port map (
            O => \N__18688\,
            I => \N__18629\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__18685\,
            I => \N__18626\
        );

    \I__2849\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18623\
        );

    \I__2848\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18618\
        );

    \I__2847\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18618\
        );

    \I__2846\ : InMux
    port map (
            O => \N__18679\,
            I => \N__18609\
        );

    \I__2845\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18609\
        );

    \I__2844\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18609\
        );

    \I__2843\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18609\
        );

    \I__2842\ : Span4Mux_s3_v
    port map (
            O => \N__18673\,
            I => \N__18606\
        );

    \I__2841\ : Span4Mux_v
    port map (
            O => \N__18670\,
            I => \N__18601\
        );

    \I__2840\ : Span4Mux_s3_v
    port map (
            O => \N__18667\,
            I => \N__18601\
        );

    \I__2839\ : CEMux
    port map (
            O => \N__18666\,
            I => \N__18592\
        );

    \I__2838\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18592\
        );

    \I__2837\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18592\
        );

    \I__2836\ : InMux
    port map (
            O => \N__18663\,
            I => \N__18592\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__18658\,
            I => \N__18589\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__18655\,
            I => \N__18586\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__18652\,
            I => \N__18577\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18577\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__18642\,
            I => \N__18577\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18577\
        );

    \I__2829\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18570\
        );

    \I__2828\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18570\
        );

    \I__2827\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18570\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__18629\,
            I => \N__18567\
        );

    \I__2825\ : Span4Mux_s1_v
    port map (
            O => \N__18626\,
            I => \N__18560\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__18623\,
            I => \N__18560\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__18618\,
            I => \N__18560\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__18609\,
            I => \N__18557\
        );

    \I__2821\ : Span4Mux_h
    port map (
            O => \N__18606\,
            I => \N__18554\
        );

    \I__2820\ : Span4Mux_h
    port map (
            O => \N__18601\,
            I => \N__18547\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__18592\,
            I => \N__18547\
        );

    \I__2818\ : Span4Mux_s3_v
    port map (
            O => \N__18589\,
            I => \N__18547\
        );

    \I__2817\ : Span4Mux_s0_v
    port map (
            O => \N__18586\,
            I => \N__18542\
        );

    \I__2816\ : Span4Mux_h
    port map (
            O => \N__18577\,
            I => \N__18542\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__18570\,
            I => \N__18539\
        );

    \I__2814\ : Span4Mux_h
    port map (
            O => \N__18567\,
            I => \N__18532\
        );

    \I__2813\ : Span4Mux_h
    port map (
            O => \N__18560\,
            I => \N__18532\
        );

    \I__2812\ : Span4Mux_h
    port map (
            O => \N__18557\,
            I => \N__18532\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__18554\,
            I => \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__18547\,
            I => \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__18542\,
            I => \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0\
        );

    \I__2808\ : Odrv4
    port map (
            O => \N__18539\,
            I => \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__18532\,
            I => \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0\
        );

    \I__2806\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__2804\ : Span4Mux_h
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__2803\ : Odrv4
    port map (
            O => \N__18512\,
            I => \PCH_PWRGD.un12_clk_100khz_2\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__18509\,
            I => \N__18505\
        );

    \I__2801\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18502\
        );

    \I__2800\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18499\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__18502\,
            I => \N__18494\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__18499\,
            I => \N__18494\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__18491\,
            I => \RSMRST_PWRGD.N_256_i\
        );

    \I__2795\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18484\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18481\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__18484\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__18481\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__2791\ : InMux
    port map (
            O => \N__18476\,
            I => \N__18472\
        );

    \I__2790\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18469\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__18472\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__18469\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__2787\ : InMux
    port map (
            O => \N__18464\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__2786\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__18455\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__2782\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__18446\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__2780\ : InMux
    port map (
            O => \N__18443\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__2778\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__18434\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__2776\ : InMux
    port map (
            O => \N__18431\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__2775\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__18425\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__2773\ : InMux
    port map (
            O => \N__18422\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__2772\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__18416\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__2770\ : InMux
    port map (
            O => \N__18413\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__18410\,
            I => \N__18407\
        );

    \I__2768\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__18404\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__2766\ : InMux
    port map (
            O => \N__18401\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__2765\ : InMux
    port map (
            O => \N__18398\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__2764\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__18392\,
            I => \N__18388\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__18391\,
            I => \N__18384\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__18388\,
            I => \N__18379\
        );

    \I__2760\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18376\
        );

    \I__2759\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18369\
        );

    \I__2758\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18369\
        );

    \I__2757\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18369\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__18379\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__18376\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__18369\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__18362\,
            I => \N__18358\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__18361\,
            I => \N__18354\
        );

    \I__2751\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18347\
        );

    \I__2750\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18347\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18347\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__18347\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__2747\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__18341\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__2745\ : InMux
    port map (
            O => \N__18338\,
            I => \POWERLED.mult1_un68_sum_cry_2_c\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__2743\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__18329\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__2741\ : InMux
    port map (
            O => \N__18326\,
            I => \POWERLED.mult1_un68_sum_cry_3_c\
        );

    \I__2740\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__18320\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__2738\ : InMux
    port map (
            O => \N__18317\,
            I => \POWERLED.mult1_un68_sum_cry_4_c\
        );

    \I__2737\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18310\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__18313\,
            I => \N__18306\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__18310\,
            I => \N__18302\
        );

    \I__2734\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18297\
        );

    \I__2733\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18297\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18294\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__18302\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__18297\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__18294\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__2727\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18281\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__2725\ : InMux
    port map (
            O => \N__18278\,
            I => \POWERLED.mult1_un68_sum_cry_5_c\
        );

    \I__2724\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__18272\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__18269\,
            I => \N__18265\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__18268\,
            I => \N__18261\
        );

    \I__2720\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18254\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18254\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18254\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__18254\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__2716\ : InMux
    port map (
            O => \N__18251\,
            I => \POWERLED.mult1_un68_sum_cry_6_c\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__18248\,
            I => \N__18245\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__18242\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__2712\ : InMux
    port map (
            O => \N__18239\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \POWERLED.mult1_un68_sum_s_8_cascade_\
        );

    \I__2710\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18229\
        );

    \I__2709\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18226\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__18229\,
            I => \N__18223\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__18226\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2706\ : Odrv12
    port map (
            O => \N__18223\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2705\ : InMux
    port map (
            O => \N__18218\,
            I => \POWERLED.un1_dutycycle_53_cry_14\
        );

    \I__2704\ : InMux
    port map (
            O => \N__18215\,
            I => \bfn_5_13_0_\
        );

    \I__2703\ : InMux
    port map (
            O => \N__18212\,
            I => \POWERLED.CO2\
        );

    \I__2702\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__2700\ : Span4Mux_s3_v
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__18200\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__2697\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18191\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__18191\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__2695\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18184\
        );

    \I__2694\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18181\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__18184\,
            I => \N__18178\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__18181\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__18178\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__2689\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18164\
        );

    \I__2688\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18164\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__18164\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__2686\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18157\
        );

    \I__2685\ : InMux
    port map (
            O => \N__18160\,
            I => \N__18154\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__18157\,
            I => \N__18151\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__18154\,
            I => \N__18148\
        );

    \I__2682\ : Span4Mux_s2_v
    port map (
            O => \N__18151\,
            I => \N__18145\
        );

    \I__2681\ : Span4Mux_s1_v
    port map (
            O => \N__18148\,
            I => \N__18142\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__18145\,
            I => \N__18139\
        );

    \I__2679\ : Span4Mux_v
    port map (
            O => \N__18142\,
            I => \N__18136\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__18139\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__18136\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__2676\ : InMux
    port map (
            O => \N__18131\,
            I => \POWERLED.un1_dutycycle_53_cry_5_cZ0\
        );

    \I__2675\ : InMux
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__18125\,
            I => \N__18121\
        );

    \I__2673\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18118\
        );

    \I__2672\ : Span4Mux_s1_v
    port map (
            O => \N__18121\,
            I => \N__18113\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__18118\,
            I => \N__18113\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__18113\,
            I => \N__18110\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__18110\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__2668\ : InMux
    port map (
            O => \N__18107\,
            I => \POWERLED.un1_dutycycle_53_cry_6_cZ0\
        );

    \I__2667\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__18101\,
            I => \N__18097\
        );

    \I__2665\ : InMux
    port map (
            O => \N__18100\,
            I => \N__18094\
        );

    \I__2664\ : Span4Mux_h
    port map (
            O => \N__18097\,
            I => \N__18089\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__18094\,
            I => \N__18089\
        );

    \I__2662\ : Span4Mux_s2_v
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__18086\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__2660\ : InMux
    port map (
            O => \N__18083\,
            I => \bfn_5_12_0_\
        );

    \I__2659\ : InMux
    port map (
            O => \N__18080\,
            I => \POWERLED.un1_dutycycle_53_cry_8_cZ0\
        );

    \I__2658\ : InMux
    port map (
            O => \N__18077\,
            I => \POWERLED.un1_dutycycle_53_cry_9_cZ0\
        );

    \I__2657\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__18071\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_14\
        );

    \I__2655\ : InMux
    port map (
            O => \N__18068\,
            I => \POWERLED.un1_dutycycle_53_cry_10\
        );

    \I__2654\ : InMux
    port map (
            O => \N__18065\,
            I => \POWERLED.un1_dutycycle_53_cry_11\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__18062\,
            I => \N__18058\
        );

    \I__2652\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18055\
        );

    \I__2651\ : InMux
    port map (
            O => \N__18058\,
            I => \N__18052\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__18055\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__18052\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__2648\ : InMux
    port map (
            O => \N__18047\,
            I => \POWERLED.un1_dutycycle_53_cry_12\
        );

    \I__2647\ : InMux
    port map (
            O => \N__18044\,
            I => \POWERLED.un1_dutycycle_53_cry_13\
        );

    \I__2646\ : InMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__2644\ : Odrv12
    port map (
            O => \N__18035\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__2643\ : InMux
    port map (
            O => \N__18032\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__18029\,
            I => \N__18024\
        );

    \I__2641\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18017\
        );

    \I__2640\ : InMux
    port map (
            O => \N__18027\,
            I => \N__18017\
        );

    \I__2639\ : InMux
    port map (
            O => \N__18024\,
            I => \N__18012\
        );

    \I__2638\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18012\
        );

    \I__2637\ : InMux
    port map (
            O => \N__18022\,
            I => \N__18009\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__18017\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__18012\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__18009\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__2633\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__17993\,
            I => \N__17989\
        );

    \I__2629\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17986\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__17989\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__17986\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__2626\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__17978\,
            I => \N__17974\
        );

    \I__2624\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17971\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__17974\,
            I => \N__17968\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__17971\,
            I => \N__17965\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__17968\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__17965\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__2619\ : InMux
    port map (
            O => \N__17960\,
            I => \POWERLED.un1_dutycycle_53_cry_0_cZ0\
        );

    \I__2618\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__17954\,
            I => \N__17950\
        );

    \I__2616\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17947\
        );

    \I__2615\ : Span4Mux_v
    port map (
            O => \N__17950\,
            I => \N__17942\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__17947\,
            I => \N__17942\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__17942\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__2612\ : InMux
    port map (
            O => \N__17939\,
            I => \POWERLED.un1_dutycycle_53_cry_1_cZ0\
        );

    \I__2611\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17932\
        );

    \I__2610\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17929\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__17932\,
            I => \N__17924\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__17929\,
            I => \N__17924\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__17921\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__2605\ : InMux
    port map (
            O => \N__17918\,
            I => \POWERLED.un1_dutycycle_53_cry_2_cZ0\
        );

    \I__2604\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17911\
        );

    \I__2603\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17908\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__17911\,
            I => \N__17905\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__17908\,
            I => \N__17902\
        );

    \I__2600\ : Span4Mux_v
    port map (
            O => \N__17905\,
            I => \N__17899\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__17902\,
            I => \N__17896\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__17899\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__17896\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__2596\ : InMux
    port map (
            O => \N__17891\,
            I => \POWERLED.un1_dutycycle_53_cry_3_cZ0\
        );

    \I__2595\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__17885\,
            I => \N__17881\
        );

    \I__2593\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17878\
        );

    \I__2592\ : Span4Mux_s2_h
    port map (
            O => \N__17881\,
            I => \N__17873\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__17878\,
            I => \N__17873\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__17873\,
            I => \N__17870\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__17870\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__2588\ : InMux
    port map (
            O => \N__17867\,
            I => \POWERLED.un1_dutycycle_53_cry_4_cZ0\
        );

    \I__2587\ : InMux
    port map (
            O => \N__17864\,
            I => \N__17861\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__17861\,
            I => \POWERLED.count_0_8\
        );

    \I__2585\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__17852\,
            I => \POWERLED.count_0_10\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__2581\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__17843\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__2579\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__17837\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__2577\ : InMux
    port map (
            O => \N__17834\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__2576\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__2574\ : Odrv12
    port map (
            O => \N__17825\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__2572\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__17813\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__2569\ : InMux
    port map (
            O => \N__17810\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__2568\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__2566\ : Odrv12
    port map (
            O => \N__17801\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__2565\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17795\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__17795\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__2563\ : InMux
    port map (
            O => \N__17792\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__17789\,
            I => \N__17785\
        );

    \I__2561\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17780\
        );

    \I__2560\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17780\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__17780\,
            I => \N__17774\
        );

    \I__2558\ : InMux
    port map (
            O => \N__17779\,
            I => \N__17769\
        );

    \I__2557\ : InMux
    port map (
            O => \N__17778\,
            I => \N__17769\
        );

    \I__2556\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17766\
        );

    \I__2555\ : Odrv12
    port map (
            O => \N__17774\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__17769\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__17766\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__17759\,
            I => \N__17756\
        );

    \I__2551\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__2549\ : Odrv12
    port map (
            O => \N__17750\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__17747\,
            I => \N__17744\
        );

    \I__2547\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17738\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__17738\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__2544\ : InMux
    port map (
            O => \N__17735\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__17732\,
            I => \N__17728\
        );

    \I__2542\ : InMux
    port map (
            O => \N__17731\,
            I => \N__17720\
        );

    \I__2541\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17720\
        );

    \I__2540\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17720\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__17720\,
            I => \N__17717\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__17714\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__2535\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17705\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__17705\,
            I => \N__17702\
        );

    \I__2533\ : Odrv12
    port map (
            O => \N__17702\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__2532\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__17696\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__2530\ : InMux
    port map (
            O => \N__17693\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__2529\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__17687\,
            I => \POWERLED.count_0_11\
        );

    \I__2527\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__17681\,
            I => \POWERLED.count_0_3\
        );

    \I__2525\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__17675\,
            I => \POWERLED.count_0_15\
        );

    \I__2523\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__17669\,
            I => \POWERLED.count_0_7\
        );

    \I__2521\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17663\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__17663\,
            I => \PCH_PWRGD.count_0_6\
        );

    \I__2519\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__17654\,
            I => \PCH_PWRGD.un2_count_1_axb_10\
        );

    \I__2516\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17647\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__17650\,
            I => \N__17643\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17637\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17626\
        );

    \I__2512\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17626\
        );

    \I__2511\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17626\
        );

    \I__2510\ : InMux
    port map (
            O => \N__17641\,
            I => \N__17626\
        );

    \I__2509\ : InMux
    port map (
            O => \N__17640\,
            I => \N__17626\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__17637\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__17626\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__2506\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__17618\,
            I => \N_187\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__17615\,
            I => \G_11_cascade_\
        );

    \I__2503\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__17609\,
            I => \POWERLED.count_0_4\
        );

    \I__2501\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__17603\,
            I => \POWERLED.count_0_2\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__17600\,
            I => \POWERLED.g0_i_o3_0_cascade_\
        );

    \I__2498\ : InMux
    port map (
            O => \N__17597\,
            I => \N__17591\
        );

    \I__2497\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17591\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__17591\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__2495\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__17585\,
            I => \POWERLED.g0_i_o3_0\
        );

    \I__2493\ : IoInMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__2491\ : Span4Mux_s3_v
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__17567\,
            I => pwrbtn_led
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__17564\,
            I => \POWERLED.curr_state_3_0_cascade_\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__17561\,
            I => \POWERLED.curr_stateZ0Z_0_cascade_\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__17558\,
            I => \POWERLED.count_0_sqmuxa_i_cascade_\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__17555\,
            I => \POWERLED.count_RNIZ0Z_0_cascade_\
        );

    \I__2483\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17546\
        );

    \I__2482\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17546\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__2480\ : Odrv12
    port map (
            O => \N__17543\,
            I => \PCH_PWRGD.count_rst_8\
        );

    \I__2479\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17536\
        );

    \I__2478\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17533\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__17536\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__17533\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__17528\,
            I => \N__17524\
        );

    \I__2474\ : InMux
    port map (
            O => \N__17527\,
            I => \N__17519\
        );

    \I__2473\ : InMux
    port map (
            O => \N__17524\,
            I => \N__17519\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__17519\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__2471\ : InMux
    port map (
            O => \N__17516\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__2470\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17510\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17507\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__17507\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__2467\ : InMux
    port map (
            O => \N__17504\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__2466\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17495\
        );

    \I__2465\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17495\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__17495\,
            I => \PCH_PWRGD.count_rst\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__17492\,
            I => \N__17489\
        );

    \I__2462\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17467\
        );

    \I__2461\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17467\
        );

    \I__2460\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17467\
        );

    \I__2459\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17467\
        );

    \I__2458\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17467\
        );

    \I__2457\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17460\
        );

    \I__2456\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17460\
        );

    \I__2455\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17460\
        );

    \I__2454\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17456\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__17480\,
            I => \N__17453\
        );

    \I__2452\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17450\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__17478\,
            I => \N__17443\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__17467\,
            I => \N__17440\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__17460\,
            I => \N__17437\
        );

    \I__2448\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17434\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__17456\,
            I => \N__17431\
        );

    \I__2446\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17428\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__17450\,
            I => \N__17425\
        );

    \I__2444\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17414\
        );

    \I__2443\ : InMux
    port map (
            O => \N__17448\,
            I => \N__17414\
        );

    \I__2442\ : InMux
    port map (
            O => \N__17447\,
            I => \N__17414\
        );

    \I__2441\ : InMux
    port map (
            O => \N__17446\,
            I => \N__17414\
        );

    \I__2440\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17414\
        );

    \I__2439\ : Span4Mux_h
    port map (
            O => \N__17440\,
            I => \N__17409\
        );

    \I__2438\ : Span4Mux_s3_h
    port map (
            O => \N__17437\,
            I => \N__17409\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__17434\,
            I => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\
        );

    \I__2436\ : Odrv4
    port map (
            O => \N__17431\,
            I => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__17428\,
            I => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__17425\,
            I => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__17414\,
            I => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__17409\,
            I => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\
        );

    \I__2431\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17370\
        );

    \I__2430\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17370\
        );

    \I__2429\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17370\
        );

    \I__2428\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17367\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17364\
        );

    \I__2426\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17359\
        );

    \I__2425\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17359\
        );

    \I__2424\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17356\
        );

    \I__2423\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17347\
        );

    \I__2422\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17347\
        );

    \I__2421\ : InMux
    port map (
            O => \N__17386\,
            I => \N__17347\
        );

    \I__2420\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17347\
        );

    \I__2419\ : InMux
    port map (
            O => \N__17384\,
            I => \N__17336\
        );

    \I__2418\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17336\
        );

    \I__2417\ : InMux
    port map (
            O => \N__17382\,
            I => \N__17336\
        );

    \I__2416\ : InMux
    port map (
            O => \N__17381\,
            I => \N__17336\
        );

    \I__2415\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17336\
        );

    \I__2414\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17323\
        );

    \I__2413\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17323\
        );

    \I__2412\ : InMux
    port map (
            O => \N__17377\,
            I => \N__17323\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__17370\,
            I => \N__17320\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__17367\,
            I => \N__17307\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__17364\,
            I => \N__17307\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17307\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17307\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__17347\,
            I => \N__17307\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__17336\,
            I => \N__17307\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17335\,
            I => \N__17295\
        );

    \I__2403\ : InMux
    port map (
            O => \N__17334\,
            I => \N__17295\
        );

    \I__2402\ : InMux
    port map (
            O => \N__17333\,
            I => \N__17295\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17332\,
            I => \N__17295\
        );

    \I__2400\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17295\
        );

    \I__2399\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17292\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__17323\,
            I => \N__17285\
        );

    \I__2397\ : Span4Mux_h
    port map (
            O => \N__17320\,
            I => \N__17285\
        );

    \I__2396\ : Span4Mux_s2_v
    port map (
            O => \N__17307\,
            I => \N__17285\
        );

    \I__2395\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17282\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__17295\,
            I => \N__17279\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__17292\,
            I => \PCH_PWRGD.N_386\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__17285\,
            I => \PCH_PWRGD.N_386\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__17282\,
            I => \PCH_PWRGD.N_386\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__17279\,
            I => \PCH_PWRGD.N_386\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__2388\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17260\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17260\
        );

    \I__2386\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17257\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__17260\,
            I => \N__17254\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__17257\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__17254\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__2382\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17246\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__17246\,
            I => \N__17242\
        );

    \I__2380\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17239\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__17242\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__17239\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__2377\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17231\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__17228\,
            I => \PCH_PWRGD.count_rst_5\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__17225\,
            I => \RSMRST_PWRGD.un4_count_9_cascade_\
        );

    \I__2373\ : InMux
    port map (
            O => \N__17222\,
            I => \N__17218\
        );

    \I__2372\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17215\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__17218\,
            I => \RSMRST_PWRGD.N_1_i\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__17215\,
            I => \RSMRST_PWRGD.N_1_i\
        );

    \I__2369\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__17207\,
            I => \RSMRST_PWRGD.un4_count_8\
        );

    \I__2367\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17201\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__17201\,
            I => \RSMRST_PWRGD.un4_count_10\
        );

    \I__2365\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__17195\,
            I => \RSMRST_PWRGD.un4_count_11\
        );

    \I__2363\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17186\
        );

    \I__2362\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17186\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__17186\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__2360\ : InMux
    port map (
            O => \N__17183\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__2359\ : InMux
    port map (
            O => \N__17180\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__2358\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17170\
        );

    \I__2357\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17175\,
            I => \N__17167\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__17170\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__17167\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__17162\,
            I => \N__17158\
        );

    \I__2352\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17155\
        );

    \I__2351\ : InMux
    port map (
            O => \N__17158\,
            I => \N__17152\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__17155\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__17152\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__2348\ : InMux
    port map (
            O => \N__17147\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__2347\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17139\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__17143\,
            I => \N__17136\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__17142\,
            I => \N__17133\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__17139\,
            I => \N__17130\
        );

    \I__2343\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17125\
        );

    \I__2342\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17125\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__17130\,
            I => \N__17122\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__17125\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__17122\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__2338\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17111\
        );

    \I__2337\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17111\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__2335\ : Span4Mux_s1_v
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__17105\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__2333\ : InMux
    port map (
            O => \N__17102\,
            I => \PCH_PWRGD.un2_count_1_cry_7\
        );

    \I__2332\ : InMux
    port map (
            O => \N__17099\,
            I => \bfn_5_3_0_\
        );

    \I__2331\ : InMux
    port map (
            O => \N__17096\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__2330\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17089\
        );

    \I__2329\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__17089\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__17086\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__2326\ : InMux
    port map (
            O => \N__17081\,
            I => \N__17075\
        );

    \I__2325\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17075\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__17075\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__2323\ : InMux
    port map (
            O => \N__17072\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__2322\ : InMux
    port map (
            O => \N__17069\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__2321\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17062\
        );

    \I__2320\ : InMux
    port map (
            O => \N__17065\,
            I => \N__17059\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__17062\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__17059\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__2317\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17048\
        );

    \I__2316\ : InMux
    port map (
            O => \N__17053\,
            I => \N__17048\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__17048\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__2314\ : InMux
    port map (
            O => \N__17045\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__17042\,
            I => \PCH_PWRGD.count_rst_7_cascade_\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__17039\,
            I => \PCH_PWRGD.countZ0Z_7_cascade_\
        );

    \I__2311\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__17033\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__2309\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17027\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__17024\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__2306\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17017\
        );

    \I__2305\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17014\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__17017\,
            I => \N__17010\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__17014\,
            I => \N__17007\
        );

    \I__2302\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17004\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__17010\,
            I => \N__17001\
        );

    \I__2300\ : Span4Mux_h
    port map (
            O => \N__17007\,
            I => \N__16998\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__17004\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__17001\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__16998\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__16991\,
            I => \N__16986\
        );

    \I__2295\ : InMux
    port map (
            O => \N__16990\,
            I => \N__16983\
        );

    \I__2294\ : InMux
    port map (
            O => \N__16989\,
            I => \N__16980\
        );

    \I__2293\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16977\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__16983\,
            I => \N__16973\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__16980\,
            I => \N__16970\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__16977\,
            I => \N__16967\
        );

    \I__2289\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16964\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__16973\,
            I => \N__16961\
        );

    \I__2287\ : Span4Mux_h
    port map (
            O => \N__16970\,
            I => \N__16958\
        );

    \I__2286\ : Span4Mux_v
    port map (
            O => \N__16967\,
            I => \N__16955\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__16964\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__16961\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__16958\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__16955\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__2281\ : InMux
    port map (
            O => \N__16946\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \I__2280\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16939\
        );

    \I__2279\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__16939\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__16936\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__2276\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__16928\,
            I => \N__16924\
        );

    \I__2274\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16921\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__16924\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__16921\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__2271\ : InMux
    port map (
            O => \N__16916\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__16913\,
            I => \N__16910\
        );

    \I__2269\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16905\
        );

    \I__2268\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16902\
        );

    \I__2267\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16899\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__16905\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__16902\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__16899\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__2263\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16886\
        );

    \I__2262\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16886\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__16886\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__2260\ : InMux
    port map (
            O => \N__16883\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \N__16877\
        );

    \I__2258\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16873\
        );

    \I__2257\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16870\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__16873\,
            I => \PCH_PWRGD.un2_count_1_axb_5\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__16870\,
            I => \PCH_PWRGD.un2_count_1_axb_5\
        );

    \I__2254\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__16862\,
            I => \N__16859\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__16859\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__2251\ : InMux
    port map (
            O => \N__16856\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__2250\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16850\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__16850\,
            I => \N__16847\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__16847\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__2247\ : InMux
    port map (
            O => \N__16844\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__2246\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__16835\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__2243\ : InMux
    port map (
            O => \N__16832\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__2242\ : InMux
    port map (
            O => \N__16829\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__2241\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16819\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__16822\,
            I => \N__16816\
        );

    \I__2238\ : Span4Mux_h
    port map (
            O => \N__16819\,
            I => \N__16810\
        );

    \I__2237\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16803\
        );

    \I__2236\ : InMux
    port map (
            O => \N__16815\,
            I => \N__16803\
        );

    \I__2235\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16803\
        );

    \I__2234\ : InMux
    port map (
            O => \N__16813\,
            I => \N__16800\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__16810\,
            I => \N__16795\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__16803\,
            I => \N__16795\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__16800\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__16795\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__16790\,
            I => \N__16786\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__16789\,
            I => \N__16782\
        );

    \I__2227\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16775\
        );

    \I__2226\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16775\
        );

    \I__2225\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16775\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__16775\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__16772\,
            I => \PCH_PWRGD.un2_count_1_axb_5_cascade_\
        );

    \I__2222\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16763\
        );

    \I__2221\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16763\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__16763\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__2219\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__16751\,
            I => \PCH_PWRGD.un12_clk_100khz_6\
        );

    \I__2215\ : InMux
    port map (
            O => \N__16748\,
            I => \N__16742\
        );

    \I__2214\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16742\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__16742\,
            I => \PCH_PWRGD.count_rst_9\
        );

    \I__2212\ : InMux
    port map (
            O => \N__16739\,
            I => \N__16736\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__16736\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__2210\ : InMux
    port map (
            O => \N__16733\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__16730\,
            I => \N__16726\
        );

    \I__2208\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16720\
        );

    \I__2207\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16720\
        );

    \I__2206\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16717\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__16720\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__16717\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__2202\ : InMux
    port map (
            O => \N__16709\,
            I => \N__16706\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__16706\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__2200\ : InMux
    port map (
            O => \N__16703\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__2199\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16697\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__16697\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__16694\,
            I => \N__16690\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__16693\,
            I => \N__16686\
        );

    \I__2195\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16679\
        );

    \I__2194\ : InMux
    port map (
            O => \N__16689\,
            I => \N__16679\
        );

    \I__2193\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16679\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__16679\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16676\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__2189\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__16667\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__2187\ : InMux
    port map (
            O => \N__16664\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__16661\,
            I => \POWERLED.mult1_un61_sum_s_8_cascade_\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__2184\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__16649\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__2181\ : InMux
    port map (
            O => \N__16646\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__2179\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16637\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__2177\ : Odrv12
    port map (
            O => \N__16634\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__2176\ : InMux
    port map (
            O => \N__16631\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__2175\ : InMux
    port map (
            O => \N__16628\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16625\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__2173\ : InMux
    port map (
            O => \N__16622\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__2172\ : InMux
    port map (
            O => \N__16619\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__2171\ : InMux
    port map (
            O => \N__16616\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__16613\,
            I => \POWERLED.mult1_un54_sum_s_8_cascade_\
        );

    \I__2169\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16607\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__16604\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__2166\ : InMux
    port map (
            O => \N__16601\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__2164\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__16592\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__2162\ : InMux
    port map (
            O => \N__16589\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__16586\,
            I => \POWERLED.un2_count_clk_17_0_a2_5_cascade_\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \POWERLED.un1_dutycycle_53_46_0_cascade_\
        );

    \I__2159\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__16577\,
            I => \N__16574\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__16574\,
            I => \POWERLED.mult1_un47_sum_i\
        );

    \I__2156\ : InMux
    port map (
            O => \N__16571\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__16568\,
            I => \N__16565\
        );

    \I__2154\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16562\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__16562\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__2152\ : InMux
    port map (
            O => \N__16559\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16553\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__16553\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__2149\ : InMux
    port map (
            O => \N__16550\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__2148\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16544\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__16544\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__2146\ : InMux
    port map (
            O => \N__16541\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__2145\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__16535\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__2143\ : InMux
    port map (
            O => \N__16532\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__2142\ : InMux
    port map (
            O => \N__16529\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__2141\ : InMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__16523\,
            I => \N__16519\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__16522\,
            I => \N__16516\
        );

    \I__2138\ : Span4Mux_v
    port map (
            O => \N__16519\,
            I => \N__16510\
        );

    \I__2137\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16503\
        );

    \I__2136\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16503\
        );

    \I__2135\ : InMux
    port map (
            O => \N__16514\,
            I => \N__16503\
        );

    \I__2134\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16500\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__16510\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__16503\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__16500\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__2129\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__16487\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__16484\,
            I => \N__16480\
        );

    \I__2126\ : InMux
    port map (
            O => \N__16483\,
            I => \N__16472\
        );

    \I__2125\ : InMux
    port map (
            O => \N__16480\,
            I => \N__16472\
        );

    \I__2124\ : InMux
    port map (
            O => \N__16479\,
            I => \N__16472\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__16472\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__2121\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__16457\,
            I => \N__16454\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__16454\,
            I => \POWERLED.un85_clk_100khz_2\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__16451\,
            I => \N__16447\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__16450\,
            I => \N__16443\
        );

    \I__2114\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16436\
        );

    \I__2113\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16436\
        );

    \I__2112\ : InMux
    port map (
            O => \N__16443\,
            I => \N__16436\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__16436\,
            I => \G_2121\
        );

    \I__2110\ : InMux
    port map (
            O => \N__16433\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__16430\,
            I => \N__16427\
        );

    \I__2108\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16424\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__16424\,
            I => \N__16421\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__16421\,
            I => \POWERLED.un85_clk_100khz_0\
        );

    \I__2105\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16415\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__16415\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__16412\,
            I => \N__16409\
        );

    \I__2102\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__16406\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__2100\ : InMux
    port map (
            O => \N__16403\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__2098\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__16394\,
            I => \N__16391\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__16391\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__2094\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__16382\,
            I => \N__16379\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__16379\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__16376\,
            I => \N__16373\
        );

    \I__2090\ : InMux
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__16370\,
            I => \N__16367\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__16367\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__2087\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__16358\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__2083\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16349\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__16349\,
            I => \N__16346\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__16346\,
            I => \N__16343\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__16343\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__2079\ : InMux
    port map (
            O => \N__16340\,
            I => \bfn_4_8_0_\
        );

    \I__2078\ : IoInMux
    port map (
            O => \N__16337\,
            I => \N__16334\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__16334\,
            I => \N__16330\
        );

    \I__2076\ : IoInMux
    port map (
            O => \N__16333\,
            I => \N__16327\
        );

    \I__2075\ : Span4Mux_s2_h
    port map (
            O => \N__16330\,
            I => \N__16324\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__16327\,
            I => \N__16321\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__16324\,
            I => \N__16318\
        );

    \I__2072\ : Span4Mux_s3_h
    port map (
            O => \N__16321\,
            I => \N__16315\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__16318\,
            I => v5s_enn
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__16315\,
            I => v5s_enn
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__16310\,
            I => \N_187_cascade_\
        );

    \I__2068\ : IoInMux
    port map (
            O => \N__16307\,
            I => \N__16303\
        );

    \I__2067\ : IoInMux
    port map (
            O => \N__16306\,
            I => \N__16300\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__16303\,
            I => \N__16297\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__16300\,
            I => \N__16293\
        );

    \I__2064\ : Span4Mux_s3_h
    port map (
            O => \N__16297\,
            I => \N__16290\
        );

    \I__2063\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16287\
        );

    \I__2062\ : IoSpan4Mux
    port map (
            O => \N__16293\,
            I => \N__16284\
        );

    \I__2061\ : Sp12to4
    port map (
            O => \N__16290\,
            I => \N__16279\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__16287\,
            I => \N__16279\
        );

    \I__2059\ : IoSpan4Mux
    port map (
            O => \N__16284\,
            I => \N__16276\
        );

    \I__2058\ : Span12Mux_v
    port map (
            O => \N__16279\,
            I => \N__16273\
        );

    \I__2057\ : IoSpan4Mux
    port map (
            O => \N__16276\,
            I => \N__16270\
        );

    \I__2056\ : Odrv12
    port map (
            O => \N__16273\,
            I => v33a_ok
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__16270\,
            I => v33a_ok
        );

    \I__2054\ : InMux
    port map (
            O => \N__16265\,
            I => \N__16262\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__16262\,
            I => \N__16259\
        );

    \I__2052\ : Odrv12
    port map (
            O => \N__16259\,
            I => v5a_ok
        );

    \I__2051\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16252\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__16255\,
            I => \N__16249\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__16252\,
            I => \N__16246\
        );

    \I__2048\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16243\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__16246\,
            I => \N__16240\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__16243\,
            I => \N__16237\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__16240\,
            I => \N__16234\
        );

    \I__2044\ : Span12Mux_s8_h
    port map (
            O => \N__16237\,
            I => \N__16231\
        );

    \I__2043\ : Span4Mux_h
    port map (
            O => \N__16234\,
            I => \N__16228\
        );

    \I__2042\ : Odrv12
    port map (
            O => \N__16231\,
            I => slp_susn
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__16228\,
            I => slp_susn
        );

    \I__2040\ : IoInMux
    port map (
            O => \N__16223\,
            I => \N__16220\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__16220\,
            I => \N__16216\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16213\
        );

    \I__2037\ : Span4Mux_s2_h
    port map (
            O => \N__16216\,
            I => \N__16210\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__16213\,
            I => \N__16207\
        );

    \I__2035\ : Sp12to4
    port map (
            O => \N__16210\,
            I => \N__16204\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__16207\,
            I => \N__16201\
        );

    \I__2033\ : Span12Mux_s11_v
    port map (
            O => \N__16204\,
            I => \N__16198\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__16201\,
            I => \N__16195\
        );

    \I__2031\ : Odrv12
    port map (
            O => \N__16198\,
            I => v1p8a_ok
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__16195\,
            I => v1p8a_ok
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__16190\,
            I => \rsmrst_pwrgd_signal_cascade_\
        );

    \I__2028\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16177\
        );

    \I__2027\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16177\
        );

    \I__2026\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16168\
        );

    \I__2025\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16168\
        );

    \I__2024\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16168\
        );

    \I__2023\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16168\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__16177\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__16168\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__16163\,
            I => \N__16160\
        );

    \I__2019\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16157\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16154\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__16151\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__16148\,
            I => \N__16145\
        );

    \I__2014\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16142\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__16142\,
            I => \N__16139\
        );

    \I__2012\ : Span4Mux_h
    port map (
            O => \N__16139\,
            I => \N__16136\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__16136\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__16133\,
            I => \N__16130\
        );

    \I__2009\ : InMux
    port map (
            O => \N__16130\,
            I => \N__16127\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__16124\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__2006\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16113\
        );

    \I__2005\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16110\
        );

    \I__2004\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16107\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16104\
        );

    \I__2002\ : InMux
    port map (
            O => \N__16117\,
            I => \N__16099\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16099\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__16113\,
            I => \N__16092\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__16110\,
            I => \N__16092\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__16107\,
            I => \N__16092\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__16104\,
            I => \N__16089\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__16099\,
            I => \N__16084\
        );

    \I__1995\ : Span4Mux_v
    port map (
            O => \N__16092\,
            I => \N__16084\
        );

    \I__1994\ : Odrv12
    port map (
            O => \N__16089\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__16084\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__1992\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16076\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__16076\,
            I => \N__16072\
        );

    \I__1990\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16069\
        );

    \I__1989\ : Span4Mux_h
    port map (
            O => \N__16072\,
            I => \N__16062\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__16069\,
            I => \N__16062\
        );

    \I__1987\ : InMux
    port map (
            O => \N__16068\,
            I => \N__16057\
        );

    \I__1986\ : InMux
    port map (
            O => \N__16067\,
            I => \N__16057\
        );

    \I__1985\ : Span4Mux_s3_h
    port map (
            O => \N__16062\,
            I => \N__16054\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__16057\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__16054\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__16049\,
            I => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2_cascade_\
        );

    \I__1981\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__16043\,
            I => \N__16040\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__16040\,
            I => \PCH_PWRGD.curr_state_7_1\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__16037\,
            I => \PCH_PWRGD.countZ0Z_15_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16031\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__16031\,
            I => \PCH_PWRGD.un12_clk_100khz_8\
        );

    \I__1975\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__16025\,
            I => \PCH_PWRGD.count_0_14\
        );

    \I__1973\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__16019\,
            I => \PCH_PWRGD.count_0_13\
        );

    \I__1971\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16013\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__16013\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__1967\ : Span4Mux_s1_v
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__16001\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__15998\,
            I => \PCH_PWRGD.count_rst_3_cascade_\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__15995\,
            I => \PCH_PWRGD.un2_count_1_axb_11_cascade_\
        );

    \I__1963\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15989\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__15989\,
            I => \PCH_PWRGD.count_rst_3\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__1960\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15977\
        );

    \I__1959\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15977\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__15977\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__1957\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__15971\,
            I => \PCH_PWRGD.un12_clk_100khz_7\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__15968\,
            I => \PCH_PWRGD.un12_clk_100khz_4_cascade_\
        );

    \I__1954\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15962\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__15959\,
            I => \PCH_PWRGD.un12_clk_100khz_5\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__15956\,
            I => \PCH_PWRGD.un12_clk_100khz_13_cascade_\
        );

    \I__1950\ : InMux
    port map (
            O => \N__15953\,
            I => \N__15947\
        );

    \I__1949\ : InMux
    port map (
            O => \N__15952\,
            I => \N__15947\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__15944\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__15941\,
            I => \PCH_PWRGD.N_1_i_cascade_\
        );

    \I__1945\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15935\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__15935\,
            I => \N__15931\
        );

    \I__1943\ : InMux
    port map (
            O => \N__15934\,
            I => \N__15928\
        );

    \I__1942\ : Odrv12
    port map (
            O => \N__15931\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__15928\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__15923\,
            I => \PCH_PWRGD.countZ0Z_9_cascade_\
        );

    \I__1939\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15917\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__15917\,
            I => \N__15914\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__15914\,
            I => \PCH_PWRGD.count_rst_6\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__15911\,
            I => \N__15907\
        );

    \I__1935\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15902\
        );

    \I__1934\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15902\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__1932\ : Span4Mux_s1_v
    port map (
            O => \N__15899\,
            I => \N__15895\
        );

    \I__1931\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15892\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__15895\,
            I => \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__15892\,
            I => \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0\
        );

    \I__1928\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__15884\,
            I => \PCH_PWRGD.curr_state_0_0\
        );

    \I__1926\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15878\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__15878\,
            I => \PCH_PWRGD.count_rst_11\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__15875\,
            I => \PCH_PWRGD.count_rst_11_cascade_\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__15872\,
            I => \PCH_PWRGD.un2_count_1_axb_3_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15863\
        );

    \I__1921\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15863\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__15863\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__15860\,
            I => \PCH_PWRGD.count_rst_10_cascade_\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__15857\,
            I => \PCH_PWRGD.countZ0Z_4_cascade_\
        );

    \I__1917\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15851\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__15851\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__1915\ : InMux
    port map (
            O => \N__15848\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__15845\,
            I => \N__15841\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__15844\,
            I => \N__15837\
        );

    \I__1912\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15830\
        );

    \I__1911\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15830\
        );

    \I__1910\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15830\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__15830\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__1908\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15824\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__15824\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__15821\,
            I => \N__15817\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__15820\,
            I => \N__15813\
        );

    \I__1904\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15806\
        );

    \I__1903\ : InMux
    port map (
            O => \N__15816\,
            I => \N__15806\
        );

    \I__1902\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15806\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__15806\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__1900\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15800\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__15800\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__15797\,
            I => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__15794\,
            I => \PCH_PWRGD.m4_0_0_cascade_\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__15791\,
            I => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__1895\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15785\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__15785\,
            I => \PCH_PWRGD.curr_state_0_1\
        );

    \I__1893\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__1891\ : Odrv12
    port map (
            O => \N__15776\,
            I => \POWERLED.un85_clk_100khz_14\
        );

    \I__1890\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__1888\ : Span4Mux_s3_v
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__15764\,
            I => vpp_ok
        );

    \I__1886\ : IoInMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__15758\,
            I => \N__15755\
        );

    \I__1884\ : Span4Mux_s2_v
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__15752\,
            I => vddq_en
        );

    \I__1882\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__15743\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__1878\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15734\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__15734\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__1876\ : InMux
    port map (
            O => \N__15731\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__1875\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15725\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__15725\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__1873\ : InMux
    port map (
            O => \N__15722\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__1872\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15716\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__15716\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__1870\ : InMux
    port map (
            O => \N__15713\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__1869\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15707\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__15707\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__1867\ : InMux
    port map (
            O => \N__15704\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__1866\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15698\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__15698\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__1864\ : InMux
    port map (
            O => \N__15695\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__1862\ : InMux
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__15680\,
            I => \POWERLED.un85_clk_100khz_8\
        );

    \I__1858\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__15674\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__15671\,
            I => \N__15666\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__15670\,
            I => \N__15663\
        );

    \I__1854\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15659\
        );

    \I__1853\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15656\
        );

    \I__1852\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15653\
        );

    \I__1851\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15650\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__15659\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__15656\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__15653\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__15650\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__1845\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__15629\,
            I => \POWERLED.un85_clk_100khz_7\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__15626\,
            I => \N__15623\
        );

    \I__1840\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__15620\,
            I => \N__15617\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__15617\,
            I => \POWERLED.un85_clk_100khz_12\
        );

    \I__1837\ : InMux
    port map (
            O => \N__15614\,
            I => \N__15611\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__15611\,
            I => \N__15608\
        );

    \I__1835\ : Span4Mux_s2_h
    port map (
            O => \N__15608\,
            I => \N__15605\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__15605\,
            I => \POWERLED.mult1_un61_sum_i_8\
        );

    \I__1833\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15599\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__15599\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__1831\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15591\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__15595\,
            I => \N__15587\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__15594\,
            I => \N__15584\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__15591\,
            I => \N__15580\
        );

    \I__1827\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15577\
        );

    \I__1826\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15574\
        );

    \I__1825\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15571\
        );

    \I__1824\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15568\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__15580\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__15577\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__15574\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__15571\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__15568\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__15557\,
            I => \N__15552\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__15556\,
            I => \N__15549\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__15555\,
            I => \N__15546\
        );

    \I__1815\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15543\
        );

    \I__1814\ : InMux
    port map (
            O => \N__15549\,
            I => \N__15538\
        );

    \I__1813\ : InMux
    port map (
            O => \N__15546\,
            I => \N__15538\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__15543\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__15538\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__1810\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15530\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__15530\,
            I => \N__15524\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__15529\,
            I => \N__15521\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15518\
        );

    \I__1806\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15515\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__15524\,
            I => \N__15512\
        );

    \I__1804\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15509\
        );

    \I__1803\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15506\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__15515\,
            I => \N__15503\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__15512\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__15509\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__15506\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__15503\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__15494\,
            I => \N__15491\
        );

    \I__1796\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15488\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__15485\,
            I => \POWERLED.un85_clk_100khz_9\
        );

    \I__1793\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__15479\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__15476\,
            I => \N__15473\
        );

    \I__1790\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15470\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__15467\,
            I => \N__15464\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__15464\,
            I => \POWERLED.un85_clk_100khz_5\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__1785\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__15455\,
            I => \POWERLED.un85_clk_100khz_11\
        );

    \I__1783\ : IoInMux
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__15449\,
            I => \N__15446\
        );

    \I__1781\ : Span4Mux_s1_h
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__15443\,
            I => v33a_enn
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__15440\,
            I => \N__15435\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__15439\,
            I => \N__15432\
        );

    \I__1777\ : InMux
    port map (
            O => \N__15438\,
            I => \N__15427\
        );

    \I__1776\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15424\
        );

    \I__1775\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15421\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15418\
        );

    \I__1773\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15415\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__15427\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__15424\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__15421\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__15418\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__15415\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__15404\,
            I => \N__15399\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__15403\,
            I => \N__15396\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__15402\,
            I => \N__15393\
        );

    \I__1764\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15390\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15385\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15385\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15390\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__15385\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__1758\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15374\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__15374\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__1755\ : InMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__15365\,
            I => \N__15362\
        );

    \I__1753\ : Span4Mux_s1_h
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__15359\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__1751\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__15350\,
            I => \POWERLED.un85_clk_100khz_13\
        );

    \I__1748\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__15344\,
            I => \POWERLED.N_4535_i\
        );

    \I__1746\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15338\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__15338\,
            I => \POWERLED.N_4536_i\
        );

    \I__1744\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15332\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__15332\,
            I => \POWERLED.N_4537_i\
        );

    \I__1742\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__15326\,
            I => \POWERLED.N_4538_i\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__15323\,
            I => \N__15320\
        );

    \I__1739\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__15317\,
            I => \POWERLED.N_4539_i\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__15314\,
            I => \N__15311\
        );

    \I__1736\ : InMux
    port map (
            O => \N__15311\,
            I => \N__15308\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__15308\,
            I => \POWERLED.N_4540_i\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__1733\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15299\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15299\,
            I => \N__15296\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__15296\,
            I => \POWERLED.N_4541_i\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15293\,
            I => \bfn_2_11_0_\
        );

    \I__1729\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15287\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__15287\,
            I => \N__15284\
        );

    \I__1727\ : Odrv12
    port map (
            O => \N__15284\,
            I => \POWERLED.un85_clk_100khz_1\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__15281\,
            I => \N__15278\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15278\,
            I => \N__15275\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__15275\,
            I => \POWERLED.N_4527_i\
        );

    \I__1723\ : InMux
    port map (
            O => \N__15272\,
            I => \N__15269\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__15269\,
            I => \POWERLED.N_4528_i\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__15266\,
            I => \N__15263\
        );

    \I__1720\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__15260\,
            I => \N__15257\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__15257\,
            I => \POWERLED.un85_clk_100khz_3\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15251\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__15251\,
            I => \POWERLED.N_4529_i\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__15248\,
            I => \N__15245\
        );

    \I__1714\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__1712\ : Span12Mux_s10_v
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__1711\ : Odrv12
    port map (
            O => \N__15236\,
            I => \POWERLED.un85_clk_100khz_4\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__15230\,
            I => \POWERLED.N_4530_i\
        );

    \I__1708\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15224\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__15224\,
            I => \POWERLED.N_4531_i\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__15221\,
            I => \N__15218\
        );

    \I__1705\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15215\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__15215\,
            I => \N__15212\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__15212\,
            I => \POWERLED.un85_clk_100khz_6\
        );

    \I__1702\ : InMux
    port map (
            O => \N__15209\,
            I => \N__15206\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__15206\,
            I => \POWERLED.N_4532_i\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15203\,
            I => \N__15200\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__15200\,
            I => \POWERLED.N_4533_i\
        );

    \I__1698\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15194\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__15194\,
            I => \POWERLED.N_4534_i\
        );

    \I__1696\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15187\
        );

    \I__1695\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15184\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__15187\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__15184\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__1692\ : InMux
    port map (
            O => \N__15179\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__15176\,
            I => \N__15172\
        );

    \I__1690\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15169\
        );

    \I__1689\ : InMux
    port map (
            O => \N__15172\,
            I => \N__15166\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__15169\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__15166\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__1686\ : InMux
    port map (
            O => \N__15161\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__1685\ : InMux
    port map (
            O => \N__15158\,
            I => \N__15154\
        );

    \I__1684\ : InMux
    port map (
            O => \N__15157\,
            I => \N__15151\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__15154\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__15151\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__1681\ : InMux
    port map (
            O => \N__15146\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__15143\,
            I => \N__15139\
        );

    \I__1679\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15136\
        );

    \I__1678\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15133\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__15136\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__15133\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__1675\ : InMux
    port map (
            O => \N__15128\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__1674\ : InMux
    port map (
            O => \N__15125\,
            I => \N__15121\
        );

    \I__1673\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15118\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__15121\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__15118\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__1670\ : InMux
    port map (
            O => \N__15113\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__1669\ : InMux
    port map (
            O => \N__15110\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15103\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15100\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__15103\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__15100\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__1664\ : InMux
    port map (
            O => \N__15095\,
            I => \N__15092\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__15092\,
            I => \N__15088\
        );

    \I__1662\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15084\
        );

    \I__1661\ : Span4Mux_h
    port map (
            O => \N__15088\,
            I => \N__15081\
        );

    \I__1660\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15078\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__15084\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__15081\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__15078\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15068\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__15068\,
            I => \N__15064\
        );

    \I__1654\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15060\
        );

    \I__1653\ : Span4Mux_h
    port map (
            O => \N__15064\,
            I => \N__15057\
        );

    \I__1652\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15054\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__15060\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__15057\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__15054\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1648\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__15044\,
            I => \N__15039\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__15043\,
            I => \N__15036\
        );

    \I__1645\ : InMux
    port map (
            O => \N__15042\,
            I => \N__15033\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__15039\,
            I => \N__15030\
        );

    \I__1643\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15027\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__15033\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__1641\ : Odrv4
    port map (
            O => \N__15030\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__15027\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__1639\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15016\
        );

    \I__1638\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15013\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__15016\,
            I => \N__15010\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__15013\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__15010\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__1634\ : InMux
    port map (
            O => \N__15005\,
            I => \N__15002\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__15002\,
            I => \POWERLED.un1_count_cry_0_i\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__14999\,
            I => \N__14995\
        );

    \I__1631\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14992\
        );

    \I__1630\ : InMux
    port map (
            O => \N__14995\,
            I => \N__14989\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__14992\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__14989\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1627\ : InMux
    port map (
            O => \N__14984\,
            I => \bfn_2_7_0_\
        );

    \I__1626\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14977\
        );

    \I__1625\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14974\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__14977\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__14974\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1622\ : InMux
    port map (
            O => \N__14969\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14966\,
            I => \N__14962\
        );

    \I__1620\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14959\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__14962\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__14959\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1617\ : InMux
    port map (
            O => \N__14954\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__1616\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14947\
        );

    \I__1615\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14944\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__14947\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__14944\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__1612\ : InMux
    port map (
            O => \N__14939\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__1611\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14932\
        );

    \I__1610\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14929\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__14932\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__14929\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__1607\ : InMux
    port map (
            O => \N__14924\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__1606\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14917\
        );

    \I__1605\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14914\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__14917\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__14914\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__1602\ : InMux
    port map (
            O => \N__14909\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__14906\,
            I => \N__14902\
        );

    \I__1600\ : InMux
    port map (
            O => \N__14905\,
            I => \N__14899\
        );

    \I__1599\ : InMux
    port map (
            O => \N__14902\,
            I => \N__14896\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__14899\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__14896\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__1596\ : InMux
    port map (
            O => \N__14891\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__1595\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14884\
        );

    \I__1594\ : InMux
    port map (
            O => \N__14887\,
            I => \N__14881\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__14884\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__14881\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__1591\ : InMux
    port map (
            O => \N__14876\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__1590\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14869\
        );

    \I__1589\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14866\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__14869\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__14866\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__1586\ : InMux
    port map (
            O => \N__14861\,
            I => \bfn_2_8_0_\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__14858\,
            I => \N__14854\
        );

    \I__1584\ : InMux
    port map (
            O => \N__14857\,
            I => \N__14851\
        );

    \I__1583\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14848\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__14851\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__14848\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1580\ : InMux
    port map (
            O => \N__14843\,
            I => \bfn_2_6_0_\
        );

    \I__1579\ : InMux
    port map (
            O => \N__14840\,
            I => \N__14836\
        );

    \I__1578\ : InMux
    port map (
            O => \N__14839\,
            I => \N__14833\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__14836\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14833\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1575\ : InMux
    port map (
            O => \N__14828\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__1574\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14821\
        );

    \I__1573\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14818\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__14821\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__14818\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1570\ : InMux
    port map (
            O => \N__14813\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \N__14806\
        );

    \I__1568\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14803\
        );

    \I__1567\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14800\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__14803\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__14800\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1564\ : InMux
    port map (
            O => \N__14795\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__1563\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14788\
        );

    \I__1562\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14785\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__14788\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__14785\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1559\ : InMux
    port map (
            O => \N__14780\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__1558\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14773\
        );

    \I__1557\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14770\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__14773\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__14770\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1554\ : InMux
    port map (
            O => \N__14765\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__1553\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14758\
        );

    \I__1552\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14755\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__14758\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__14755\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1549\ : InMux
    port map (
            O => \N__14750\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__1548\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14743\
        );

    \I__1547\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14740\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__14743\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__14740\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1544\ : InMux
    port map (
            O => \N__14735\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__14732\,
            I => \N__14729\
        );

    \I__1542\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14720\
        );

    \I__1540\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14713\
        );

    \I__1539\ : InMux
    port map (
            O => \N__14724\,
            I => \N__14713\
        );

    \I__1538\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14713\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__14720\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__14713\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__1535\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__14705\,
            I => \N__14700\
        );

    \I__1533\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14695\
        );

    \I__1532\ : InMux
    port map (
            O => \N__14703\,
            I => \N__14695\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__14700\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__14695\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__1529\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14687\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__14681\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__1525\ : InMux
    port map (
            O => \N__14678\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__1524\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14671\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__14674\,
            I => \N__14667\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__14671\,
            I => \N__14664\
        );

    \I__1521\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14659\
        );

    \I__1520\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14659\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__14664\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__14659\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__1517\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__14648\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__1514\ : InMux
    port map (
            O => \N__14645\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__1513\ : InMux
    port map (
            O => \N__14642\,
            I => \N__14639\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__14639\,
            I => \N__14635\
        );

    \I__1511\ : InMux
    port map (
            O => \N__14638\,
            I => \N__14631\
        );

    \I__1510\ : Span4Mux_h
    port map (
            O => \N__14635\,
            I => \N__14628\
        );

    \I__1509\ : InMux
    port map (
            O => \N__14634\,
            I => \N__14625\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__14631\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__14628\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__14625\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1505\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__14612\,
            I => \N__14609\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__14609\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__1501\ : InMux
    port map (
            O => \N__14606\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__1500\ : InMux
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__14597\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__1497\ : InMux
    port map (
            O => \N__14594\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__1496\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14588\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__14585\,
            I => \N__14582\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__14582\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__1492\ : InMux
    port map (
            O => \N__14579\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__1491\ : InMux
    port map (
            O => \N__14576\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__1490\ : InMux
    port map (
            O => \N__14573\,
            I => \N__14569\
        );

    \I__1489\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14566\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__14569\,
            I => \N__14563\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__14566\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__14563\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1485\ : InMux
    port map (
            O => \N__14558\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14551\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14554\,
            I => \N__14548\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__14551\,
            I => \DSW_PWRGD.countZ0Z_9\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__14548\,
            I => \DSW_PWRGD.countZ0Z_9\
        );

    \I__1480\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14539\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14536\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__14539\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__14536\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__14531\,
            I => \N__14528\
        );

    \I__1475\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14524\
        );

    \I__1474\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14521\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__14524\,
            I => \N__14518\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__14521\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__14518\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__1470\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14509\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14506\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__14509\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__14506\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__14501\,
            I => \PCH_PWRGD.N_2126_i_cascade_\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__14498\,
            I => \PCH_PWRGD.N_381_cascade_\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14495\,
            I => \N__14489\
        );

    \I__1463\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14489\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__14489\,
            I => \PCH_PWRGD.N_254_0\
        );

    \I__1461\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14482\
        );

    \I__1460\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14479\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__14482\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__14479\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__1457\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14470\
        );

    \I__1456\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14467\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__14470\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__14467\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__14462\,
            I => \N__14458\
        );

    \I__1452\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14455\
        );

    \I__1451\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14452\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__14455\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__14452\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__1448\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14443\
        );

    \I__1447\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14440\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__14443\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__14440\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__1444\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14432\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__14432\,
            I => \DSW_PWRGD.un4_count_11\
        );

    \I__1442\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14426\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__14426\,
            I => \DSW_PWRGD.un4_count_10\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__14423\,
            I => \DSW_PWRGD.un4_count_8_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14417\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__14417\,
            I => \DSW_PWRGD.un4_count_9\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__14414\,
            I => \N__14409\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__14413\,
            I => \N__14406\
        );

    \I__1435\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14399\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14399\
        );

    \I__1433\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14399\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__14399\,
            I => \N__14396\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__14396\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__1430\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14390\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__14390\,
            I => \PCH_PWRGD.N_381\
        );

    \I__1428\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14383\
        );

    \I__1427\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14380\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__14383\,
            I => \PCH_PWRGD.N_2126_i\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__14380\,
            I => \PCH_PWRGD.N_2126_i\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__14375\,
            I => \N__14372\
        );

    \I__1423\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14366\
        );

    \I__1422\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14361\
        );

    \I__1421\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14361\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14358\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__14366\,
            I => \N__14351\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__14361\,
            I => \N__14351\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__14358\,
            I => \N__14351\
        );

    \I__1416\ : Span12Mux_s8_v
    port map (
            O => \N__14351\,
            I => \N__14348\
        );

    \I__1415\ : Odrv12
    port map (
            O => \N__14348\,
            I => vr_ready_vccin
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__14345\,
            I => \PCH_PWRGD.N_255_0_cascade_\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__14342\,
            I => \PCH_PWRGD.count_RNIZ0Z_1_cascade_\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__14339\,
            I => \N__14336\
        );

    \I__1411\ : InMux
    port map (
            O => \N__14336\,
            I => \N__14333\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__14333\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14330\,
            I => \N__14326\
        );

    \I__1408\ : InMux
    port map (
            O => \N__14329\,
            I => \N__14323\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__14326\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__14323\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__1405\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14314\
        );

    \I__1404\ : InMux
    port map (
            O => \N__14317\,
            I => \N__14311\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__14314\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__14311\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__14306\,
            I => \N__14302\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14299\
        );

    \I__1399\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14296\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__14299\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__14296\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__1396\ : InMux
    port map (
            O => \N__14291\,
            I => \N__14287\
        );

    \I__1395\ : InMux
    port map (
            O => \N__14290\,
            I => \N__14284\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__14287\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__14284\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14273\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14273\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14273\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__14270\,
            I => \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0_cascade_\
        );

    \I__1388\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14263\
        );

    \I__1387\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14260\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14257\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__14260\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__14257\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__1383\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14248\
        );

    \I__1382\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14245\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__14248\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__14245\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__14240\,
            I => \N__14236\
        );

    \I__1378\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14233\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14230\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__14233\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__14230\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__1374\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14221\
        );

    \I__1373\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14218\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__14221\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__14218\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__1370\ : InMux
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__14210\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__1368\ : InMux
    port map (
            O => \N__14207\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__1367\ : InMux
    port map (
            O => \N__14204\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__14201\,
            I => \POWERLED.mult1_un103_sum_s_8_cascade_\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__14198\,
            I => \N__14193\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__14197\,
            I => \N__14190\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__14196\,
            I => \N__14187\
        );

    \I__1362\ : InMux
    port map (
            O => \N__14193\,
            I => \N__14184\
        );

    \I__1361\ : InMux
    port map (
            O => \N__14190\,
            I => \N__14179\
        );

    \I__1360\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14179\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__14184\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__14179\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__14174\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__14171\,
            I => \PCH_PWRGD.count_rst_14_cascade_\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__14168\,
            I => \PCH_PWRGD.countZ0Z_0_cascade_\
        );

    \I__1354\ : InMux
    port map (
            O => \N__14165\,
            I => \N__14162\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__14162\,
            I => \PCH_PWRGD.count_RNIZ0Z_1\
        );

    \I__1352\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14156\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__14156\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__1350\ : InMux
    port map (
            O => \N__14153\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14147\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__14147\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__1347\ : InMux
    port map (
            O => \N__14144\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__1346\ : InMux
    port map (
            O => \N__14141\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__1345\ : InMux
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__14135\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__1343\ : InMux
    port map (
            O => \N__14132\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__1342\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14126\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__14126\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__1340\ : InMux
    port map (
            O => \N__14123\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14117\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__14117\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__1337\ : InMux
    port map (
            O => \N__14114\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__1336\ : InMux
    port map (
            O => \N__14111\,
            I => \N__14108\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__14108\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__1334\ : InMux
    port map (
            O => \N__14105\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14099\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__14099\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__1331\ : InMux
    port map (
            O => \N__14096\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__1330\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14090\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__14090\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__1328\ : InMux
    port map (
            O => \N__14087\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__1327\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14081\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__14081\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__1325\ : InMux
    port map (
            O => \N__14078\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__1324\ : InMux
    port map (
            O => \N__14075\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__14072\,
            I => \POWERLED.mult1_un117_sum_s_8_cascade_\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__14069\,
            I => \N__14064\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__14068\,
            I => \N__14061\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__14067\,
            I => \N__14058\
        );

    \I__1319\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14055\
        );

    \I__1318\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14050\
        );

    \I__1317\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14050\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__14055\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__14050\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__1314\ : InMux
    port map (
            O => \N__14045\,
            I => \N__14042\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__14042\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__1312\ : InMux
    port map (
            O => \N__14039\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__1311\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14033\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__14033\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__1309\ : InMux
    port map (
            O => \N__14030\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__1308\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14024\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__14024\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__1306\ : InMux
    port map (
            O => \N__14021\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__1305\ : InMux
    port map (
            O => \N__14018\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__1304\ : InMux
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__14012\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__1302\ : InMux
    port map (
            O => \N__14009\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__1301\ : InMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__14003\,
            I => \N__13999\
        );

    \I__1299\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13996\
        );

    \I__1298\ : Odrv12
    port map (
            O => \N__13999\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__13996\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__1296\ : InMux
    port map (
            O => \N__13991\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__1295\ : InMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__13985\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__1293\ : InMux
    port map (
            O => \N__13982\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__1292\ : InMux
    port map (
            O => \N__13979\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__1291\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13968\
        );

    \I__1290\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13968\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__13974\,
            I => \N__13965\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13962\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__13968\,
            I => \N__13957\
        );

    \I__1286\ : InMux
    port map (
            O => \N__13965\,
            I => \N__13954\
        );

    \I__1285\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13949\
        );

    \I__1284\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13949\
        );

    \I__1283\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13946\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__13957\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__13954\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__13949\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__13946\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \POWERLED.mult1_un124_sum_s_8_cascade_\
        );

    \I__1277\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__13931\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__1275\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13925\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__13925\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__1273\ : InMux
    port map (
            O => \N__13922\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__1272\ : InMux
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__13916\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__1270\ : InMux
    port map (
            O => \N__13913\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__1269\ : InMux
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__13907\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__1267\ : InMux
    port map (
            O => \N__13904\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__1266\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__13898\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__1264\ : InMux
    port map (
            O => \N__13895\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__1263\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__13889\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__1261\ : InMux
    port map (
            O => \N__13886\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__1259\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__13874\,
            I => \POWERLED.mult1_un131_sum_axb_7_l_fx\
        );

    \I__1256\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__13868\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__1254\ : InMux
    port map (
            O => \N__13865\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__1253\ : InMux
    port map (
            O => \N__13862\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__1251\ : InMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__13853\,
            I => \POWERLED.mult1_un131_sum_axb_4_l_fx\
        );

    \I__1249\ : InMux
    port map (
            O => \N__13850\,
            I => \N__13844\
        );

    \I__1248\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13844\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__13844\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__1246\ : InMux
    port map (
            O => \N__13841\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__1245\ : InMux
    port map (
            O => \N__13838\,
            I => \N__13835\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__13835\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__1243\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13829\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__13829\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__1241\ : InMux
    port map (
            O => \N__13826\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__1240\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__13820\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__1238\ : InMux
    port map (
            O => \N__13817\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__1237\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__13811\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__1235\ : InMux
    port map (
            O => \N__13808\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__13805\,
            I => \N__13802\
        );

    \I__1233\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13799\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__13799\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__1231\ : InMux
    port map (
            O => \N__13796\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__1230\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13790\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__13790\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__1228\ : InMux
    port map (
            O => \N__13787\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__1227\ : InMux
    port map (
            O => \N__13784\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__13781\,
            I => \N__13777\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__13780\,
            I => \N__13774\
        );

    \I__1224\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13769\
        );

    \I__1223\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13764\
        );

    \I__1222\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13764\
        );

    \I__1221\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13761\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__13769\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__13764\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__13761\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__13754\,
            I => \POWERLED.mult1_un138_sum_s_8_cascade_\
        );

    \I__1216\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13748\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__13748\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__1214\ : InMux
    port map (
            O => \N__13745\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__1213\ : InMux
    port map (
            O => \N__13742\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__1212\ : InMux
    port map (
            O => \N__13739\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__1211\ : InMux
    port map (
            O => \N__13736\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__1210\ : InMux
    port map (
            O => \N__13733\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__1209\ : InMux
    port map (
            O => \N__13730\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__1208\ : InMux
    port map (
            O => \N__13727\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__13724\,
            I => \N__13720\
        );

    \I__1206\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13712\
        );

    \I__1205\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13712\
        );

    \I__1204\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13712\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__13712\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__1202\ : InMux
    port map (
            O => \N__13709\,
            I => \bfn_1_4_0_\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__13706\,
            I => \N__13702\
        );

    \I__1200\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13699\
        );

    \I__1199\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13696\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__13699\,
            I => \N__13691\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__13696\,
            I => \N__13691\
        );

    \I__1196\ : Odrv12
    port map (
            O => \N__13691\,
            I => \DSW_PWRGD.un1_curr_state10_0\
        );

    \I__1195\ : InMux
    port map (
            O => \N__13688\,
            I => \N__13673\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13673\
        );

    \I__1193\ : InMux
    port map (
            O => \N__13686\,
            I => \N__13673\
        );

    \I__1192\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13673\
        );

    \I__1191\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13673\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__13673\,
            I => \N__13670\
        );

    \I__1189\ : IoSpan4Mux
    port map (
            O => \N__13670\,
            I => \N__13667\
        );

    \I__1188\ : IoSpan4Mux
    port map (
            O => \N__13667\,
            I => \N__13664\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__13664\,
            I => v33dsw_ok
        );

    \I__1186\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13646\
        );

    \I__1185\ : InMux
    port map (
            O => \N__13660\,
            I => \N__13646\
        );

    \I__1184\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13646\
        );

    \I__1183\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13646\
        );

    \I__1182\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13646\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__13646\,
            I => \DSW_PWRGD.curr_stateZ0Z_1\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__13643\,
            I => \N__13638\
        );

    \I__1179\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13627\
        );

    \I__1178\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13627\
        );

    \I__1177\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13627\
        );

    \I__1176\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13627\
        );

    \I__1175\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13624\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__13627\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__13624\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__13619\,
            I => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\
        );

    \I__1171\ : SRMux
    port map (
            O => \N__13616\,
            I => \N__13611\
        );

    \I__1170\ : SRMux
    port map (
            O => \N__13615\,
            I => \N__13608\
        );

    \I__1169\ : SRMux
    port map (
            O => \N__13614\,
            I => \N__13605\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__13611\,
            I => \N__13602\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__13608\,
            I => \N__13599\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__13605\,
            I => \N__13596\
        );

    \I__1165\ : Span4Mux_s3_v
    port map (
            O => \N__13602\,
            I => \N__13591\
        );

    \I__1164\ : Span4Mux_s1_h
    port map (
            O => \N__13599\,
            I => \N__13591\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__13596\,
            I => \G_27\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__13591\,
            I => \G_27\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__13586\,
            I => \G_27_cascade_\
        );

    \I__1160\ : CEMux
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13577\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__13577\,
            I => \DSW_PWRGD.N_27_1\
        );

    \I__1157\ : InMux
    port map (
            O => \N__13574\,
            I => \DSW_PWRGD.un1_count_1_cry_5\
        );

    \I__1156\ : InMux
    port map (
            O => \N__13571\,
            I => \DSW_PWRGD.un1_count_1_cry_6\
        );

    \I__1155\ : InMux
    port map (
            O => \N__13568\,
            I => \bfn_1_3_0_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__13565\,
            I => \DSW_PWRGD.un1_count_1_cry_8\
        );

    \I__1153\ : InMux
    port map (
            O => \N__13562\,
            I => \DSW_PWRGD.un1_count_1_cry_9\
        );

    \I__1152\ : InMux
    port map (
            O => \N__13559\,
            I => \DSW_PWRGD.un1_count_1_cry_10\
        );

    \I__1151\ : InMux
    port map (
            O => \N__13556\,
            I => \DSW_PWRGD.un1_count_1_cry_11\
        );

    \I__1150\ : InMux
    port map (
            O => \N__13553\,
            I => \DSW_PWRGD.un1_count_1_cry_12\
        );

    \I__1149\ : InMux
    port map (
            O => \N__13550\,
            I => \DSW_PWRGD.un1_count_1_cry_13\
        );

    \I__1148\ : InMux
    port map (
            O => \N__13547\,
            I => \DSW_PWRGD.un1_count_1_cry_0\
        );

    \I__1147\ : InMux
    port map (
            O => \N__13544\,
            I => \DSW_PWRGD.un1_count_1_cry_1\
        );

    \I__1146\ : InMux
    port map (
            O => \N__13541\,
            I => \DSW_PWRGD.un1_count_1_cry_2\
        );

    \I__1145\ : InMux
    port map (
            O => \N__13538\,
            I => \DSW_PWRGD.un1_count_1_cry_3\
        );

    \I__1144\ : InMux
    port map (
            O => \N__13535\,
            I => \DSW_PWRGD.un1_count_1_cry_4\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un3_count_off_1_cry_8\,
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_cry_8\,
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_4_8_0_\
        );

    \IN_MUX_bfv_2_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_5_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_7_cZ0\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_7\,
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_15\,
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_1_4_0_\
        );

    \N_579_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23806\,
            GLOBALBUFFEROUTPUT => \N_579_g\
        );

    \N_27_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25922\,
            GLOBALBUFFEROUTPUT => \N_27_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \DSW_PWRGD.count_0_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29557\,
            in1 => \N__14305\,
            in2 => \N__13706\,
            in3 => \N__13705\,
            lcout => \DSW_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_0\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_1_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29553\,
            in1 => \N__14291\,
            in2 => \_gnd_net_\,
            in3 => \N__13547\,
            lcout => \DSW_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_0\,
            carryout => \DSW_PWRGD.un1_count_1_cry_1\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_2_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29558\,
            in1 => \N__14513\,
            in2 => \_gnd_net_\,
            in3 => \N__13544\,
            lcout => \DSW_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_1\,
            carryout => \DSW_PWRGD.un1_count_1_cry_2\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_3_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29554\,
            in1 => \N__14330\,
            in2 => \_gnd_net_\,
            in3 => \N__13541\,
            lcout => \DSW_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_2\,
            carryout => \DSW_PWRGD.un1_count_1_cry_3\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_4_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29559\,
            in1 => \N__14318\,
            in2 => \_gnd_net_\,
            in3 => \N__13538\,
            lcout => \DSW_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_3\,
            carryout => \DSW_PWRGD.un1_count_1_cry_4\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_5_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29555\,
            in1 => \N__14225\,
            in2 => \_gnd_net_\,
            in3 => \N__13535\,
            lcout => \DSW_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_4\,
            carryout => \DSW_PWRGD.un1_count_1_cry_5\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_6_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29560\,
            in1 => \N__14239\,
            in2 => \_gnd_net_\,
            in3 => \N__13574\,
            lcout => \DSW_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_5\,
            carryout => \DSW_PWRGD.un1_count_1_cry_6\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_7_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29556\,
            in1 => \N__14543\,
            in2 => \_gnd_net_\,
            in3 => \N__13571\,
            lcout => \DSW_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_6\,
            carryout => \DSW_PWRGD.un1_count_1_cry_7\,
            clk => \N__32928\,
            ce => 'H',
            sr => \N__13616\
        );

    \DSW_PWRGD.count_8_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29574\,
            in1 => \N__14527\,
            in2 => \_gnd_net_\,
            in3 => \N__13568\,
            lcout => \DSW_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_8\,
            clk => \N__32973\,
            ce => 'H',
            sr => \N__13614\
        );

    \DSW_PWRGD.count_9_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29570\,
            in1 => \N__14555\,
            in2 => \_gnd_net_\,
            in3 => \N__13565\,
            lcout => \DSW_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_8\,
            carryout => \DSW_PWRGD.un1_count_1_cry_9\,
            clk => \N__32973\,
            ce => 'H',
            sr => \N__13614\
        );

    \DSW_PWRGD.count_10_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29571\,
            in1 => \N__14252\,
            in2 => \_gnd_net_\,
            in3 => \N__13562\,
            lcout => \DSW_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_9\,
            carryout => \DSW_PWRGD.un1_count_1_cry_10\,
            clk => \N__32973\,
            ce => 'H',
            sr => \N__13614\
        );

    \DSW_PWRGD.count_11_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29568\,
            in1 => \N__14266\,
            in2 => \_gnd_net_\,
            in3 => \N__13559\,
            lcout => \DSW_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_10\,
            carryout => \DSW_PWRGD.un1_count_1_cry_11\,
            clk => \N__32973\,
            ce => 'H',
            sr => \N__13614\
        );

    \DSW_PWRGD.count_12_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29572\,
            in1 => \N__14486\,
            in2 => \_gnd_net_\,
            in3 => \N__13556\,
            lcout => \DSW_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_11\,
            carryout => \DSW_PWRGD.un1_count_1_cry_12\,
            clk => \N__32973\,
            ce => 'H',
            sr => \N__13614\
        );

    \DSW_PWRGD.count_13_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29569\,
            in1 => \N__14474\,
            in2 => \_gnd_net_\,
            in3 => \N__13553\,
            lcout => \DSW_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_12\,
            carryout => \DSW_PWRGD.un1_count_1_cry_13\,
            clk => \N__32973\,
            ce => 'H',
            sr => \N__13614\
        );

    \DSW_PWRGD.count_14_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29573\,
            in1 => \N__14461\,
            in2 => \_gnd_net_\,
            in3 => \N__13550\,
            lcout => \DSW_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_13\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14\,
            clk => \N__32973\,
            ce => 'H',
            sr => \N__13614\
        );

    \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27470\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_14\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_15_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14447\,
            in2 => \_gnd_net_\,
            in3 => \N__13709\,
            lcout => \DSW_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32959\,
            ce => \N__13583\,
            sr => \N__13615\
        );

    \DSW_PWRGD.DSW_PWROK_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13684\,
            in1 => \N__13659\,
            in2 => \_gnd_net_\,
            in3 => \N__13641\,
            lcout => dsw_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32974\,
            ce => \N__29408\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNIADII_0_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__13658\,
            in1 => \N__13636\,
            in2 => \_gnd_net_\,
            in3 => \N__13687\,
            lcout => \DSW_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_0_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__13685\,
            in1 => \N__13660\,
            in2 => \N__14414\,
            in3 => \N__13642\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32974\,
            ce => \N__29408\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_1_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001110"
        )
    port map (
            in0 => \N__13661\,
            in1 => \N__13686\,
            in2 => \N__13643\,
            in3 => \N__14412\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32974\,
            ce => \N__29408\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNILLF15_0_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011101"
        )
    port map (
            in0 => \N__13688\,
            in1 => \N__13657\,
            in2 => \N__14413\,
            in3 => \N__13637\,
            lcout => OPEN,
            ltout => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.G_27_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13619\,
            in3 => \N__29541\,
            lcout => \G_27\,
            ltout => \G_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNO_0_15_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29542\,
            in1 => \_gnd_net_\,
            in2 => \N__13586\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.N_27_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14824\,
            in1 => \N__14839\,
            in2 => \N__14858\,
            in3 => \N__14573\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14791\,
            in1 => \N__14776\,
            in2 => \N__14810\,
            in3 => \N__14761\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14746\,
            in1 => \N__14965\,
            in2 => \N__14999\,
            in3 => \N__14980\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14935\,
            in1 => \N__14950\,
            in2 => \N__14906\,
            in3 => \N__14920\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15190\,
            in1 => \N__14872\,
            in2 => \N__15176\,
            in3 => \N__14887\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14703\,
            in1 => \N__14634\,
            in2 => \N__14674\,
            in3 => \N__14723\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__14724\,
            in1 => \_gnd_net_\,
            in2 => \N__26030\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__15042\,
            in1 => \N__26003\,
            in2 => \_gnd_net_\,
            in3 => \N__14725\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14690\,
            in2 => \N__26027\,
            in3 => \N__14704\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15157\,
            in1 => \N__15124\,
            in2 => \N__15143\,
            in3 => \N__15106\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14654\,
            in2 => \N__26028\,
            in3 => \N__14670\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__14603\,
            in1 => \N__26002\,
            in2 => \_gnd_net_\,
            in3 => \N__15067\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__14591\,
            in1 => \_gnd_net_\,
            in2 => \N__26029\,
            in3 => \N__15091\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__23807\,
            in1 => \N__20545\,
            in2 => \N__21794\,
            in3 => \N__20531\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__21721\,
            in1 => \N__23808\,
            in2 => \N__21793\,
            in3 => \N__21707\,
            lcout => \POWERLED.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__14618\,
            in1 => \N__14638\,
            in2 => \_gnd_net_\,
            in3 => \N__26026\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14006\,
            in2 => \_gnd_net_\,
            in3 => \N__13976\,
            lcout => \POWERLED.mult1_un131_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17778\,
            lcout => \POWERLED.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18002\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13719\,
            in2 => \N__15371\,
            in3 => \N__13742\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13832\,
            in2 => \N__13724\,
            in3 => \N__13739\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13823\,
            in2 => \N__13781\,
            in3 => \N__13736\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13814\,
            in2 => \N__13780\,
            in3 => \N__13733\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17777\,
            in1 => \N__13723\,
            in2 => \N__13805\,
            in3 => \N__13730\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13727\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13773\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17977\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15482\,
            in2 => \N__15402\,
            in3 => \N__13826\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13751\,
            in2 => \N__15404\,
            in3 => \N__13817\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13910\,
            in2 => \N__15439\,
            in3 => \N__13808\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13901\,
            in2 => \N__15440\,
            in3 => \N__13796\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13772\,
            in1 => \N__13892\,
            in2 => \N__15403\,
            in3 => \N__13787\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13784\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => \POWERLED.mult1_un138_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13754\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17957\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13934\,
            in2 => \N__15380\,
            in3 => \N__13745\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13850\,
            in2 => \N__13859\,
            in3 => \N__13904\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13838\,
            in2 => \N__13974\,
            in3 => \N__13895\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14015\,
            in2 => \N__13973\,
            in3 => \N__13886\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15430\,
            in1 => \N__14002\,
            in2 => \N__13883\,
            in3 => \N__13865\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13988\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13862\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__13849\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13961\,
            lcout => \POWERLED.mult1_un131_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17936\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15677\,
            in2 => \N__14067\,
            in3 => \N__13841\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13928\,
            in2 => \N__14069\,
            in3 => \N__14018\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13919\,
            in2 => \N__15670\,
            in3 => \N__14009\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14102\,
            in2 => \N__15671\,
            in3 => \N__13991\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13960\,
            in1 => \N__14093\,
            in2 => \N__14068\,
            in3 => \N__13982\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13979\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => \POWERLED.mult1_un124_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13937\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17915\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15602\,
            in2 => \N__15555\,
            in3 => \N__13922\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14045\,
            in2 => \N__15557\,
            in3 => \N__13913\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14036\,
            in2 => \N__15594\,
            in3 => \N__14096\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14027\,
            in2 => \N__15595\,
            in3 => \N__14087\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15662\,
            in1 => \N__14159\,
            in2 => \N__15556\,
            in3 => \N__14078\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14075\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => \POWERLED.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14072\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17888\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15827\,
            in2 => \N__14196\,
            in3 => \N__14039\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14138\,
            in2 => \N__14198\,
            in3 => \N__14030\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14129\,
            in2 => \N__15528\,
            in3 => \N__14021\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14120\,
            in2 => \N__15529\,
            in3 => \N__14153\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15583\,
            in1 => \N__14111\,
            in2 => \N__14197\,
            in3 => \N__14144\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14141\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18161\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15803\,
            in2 => \N__15820\,
            in3 => \N__14132\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15816\,
            in2 => \N__15740\,
            in3 => \N__14123\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15728\,
            in2 => \N__21891\,
            in3 => \N__14114\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15719\,
            in2 => \N__21892\,
            in3 => \N__14105\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15527\,
            in1 => \N__15710\,
            in2 => \N__15821\,
            in3 => \N__14207\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15701\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14204\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => \POWERLED.mult1_un103_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14201\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI8CTK3_1_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__17332\,
            in1 => \N__18635\,
            in2 => \N__14339\,
            in3 => \N__14165\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNI16MB1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__17116\,
            in1 => \N__17333\,
            in2 => \N__17142\,
            in3 => \N__17483\,
            lcout => \PCH_PWRGD.count_rst_6\,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIDC024_8_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15934\,
            in2 => \N__14174\,
            in3 => \N__18636\,
            lcout => \PCH_PWRGD.un2_count_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI3DJU_0_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__16976\,
            in1 => \N__17482\,
            in2 => \_gnd_net_\,
            in3 => \N__17331\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI7BTK3_0_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16010\,
            in2 => \N__14171\,
            in3 => \N__18634\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => \PCH_PWRGD.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI_1_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14168\,
            in3 => \N__17013\,
            lcout => \PCH_PWRGD.count_RNIZ0Z_1\,
            ltout => \PCH_PWRGD.count_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_1_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__17334\,
            in1 => \_gnd_net_\,
            in2 => \N__14342\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32844\,
            ce => \N__18701\,
            sr => \N__18879\
        );

    \PCH_PWRGD.count_8_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__17117\,
            in1 => \N__17335\,
            in2 => \N__17143\,
            in3 => \N__17484\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32844\,
            ce => \N__18701\,
            sr => \N__18879\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIB2J23_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20326\,
            in2 => \_gnd_net_\,
            in3 => \N__30585\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNI8U0P_0_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14329\,
            in1 => \N__14317\,
            in2 => \N__14306\,
            in3 => \N__14290\,
            lcout => \DSW_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__14279\,
            in1 => \N__15898\,
            in2 => \N__31802\,
            in3 => \N__14495\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17306\,
            in2 => \_gnd_net_\,
            in3 => \N__32004\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI3DJU_0_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14386\,
            in1 => \N__16120\,
            in2 => \N__14375\,
            in3 => \N__30584\,
            lcout => \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0\,
            ltout => \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIM8IJ2_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__14494\,
            in1 => \N__14278\,
            in2 => \N__14270\,
            in3 => \N__31795\,
            lcout => \PCH_PWRGD_delayed_vccin_ok\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIEFB91_5_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14267\,
            in1 => \N__14251\,
            in2 => \N__14240\,
            in3 => \N__14224\,
            lcout => \DSW_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIQG1P_2_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14554\,
            in1 => \N__14542\,
            in2 => \N__14531\,
            in3 => \N__14512\,
            lcout => \DSW_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16075\,
            lcout => \PCH_PWRGD.N_2126_i\,
            ltout => \PCH_PWRGD.N_2126_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14501\,
            in3 => \N__16119\,
            lcout => \PCH_PWRGD.N_381\,
            ltout => \PCH_PWRGD.N_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI3DJU_0_0_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__30549\,
            in1 => \_gnd_net_\,
            in2 => \N__14498\,
            in3 => \N__14371\,
            lcout => \PCH_PWRGD.N_254_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14485\,
            in1 => \N__14473\,
            in2 => \N__14462\,
            in3 => \N__14446\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.un4_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIB8TE4_0_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14435\,
            in1 => \N__14429\,
            in2 => \N__14423\,
            in3 => \N__14420\,
            lcout => \DSW_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14370\,
            in1 => \N__14393\,
            in2 => \_gnd_net_\,
            in3 => \N__30548\,
            lcout => \PCH_PWRGD.N_386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__14387\,
            in1 => \N__14369\,
            in2 => \_gnd_net_\,
            in3 => \N__30583\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.N_255_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI7EHJ2_0_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000000"
        )
    port map (
            in0 => \N__16121\,
            in1 => \N__17330\,
            in2 => \N__14345\,
            in3 => \N__31793\,
            lcout => \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15047\,
            in2 => \N__14732\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_5_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14708\,
            in2 => \_gnd_net_\,
            in3 => \N__14678\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14675\,
            in2 => \_gnd_net_\,
            in3 => \N__14645\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14642\,
            in2 => \_gnd_net_\,
            in3 => \N__14606\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15071\,
            in2 => \_gnd_net_\,
            in3 => \N__14594\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15095\,
            in2 => \_gnd_net_\,
            in3 => \N__14579\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15019\,
            in2 => \_gnd_net_\,
            in3 => \N__14576\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__33086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14572\,
            in2 => \_gnd_net_\,
            in3 => \N__14558\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__33086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14857\,
            in2 => \_gnd_net_\,
            in3 => \N__14843\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14840\,
            in2 => \_gnd_net_\,
            in3 => \N__14828\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14825\,
            in2 => \_gnd_net_\,
            in3 => \N__14813\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14809\,
            in2 => \_gnd_net_\,
            in3 => \N__14795\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14792\,
            in2 => \_gnd_net_\,
            in3 => \N__14780\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14777\,
            in2 => \_gnd_net_\,
            in3 => \N__14765\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14762\,
            in2 => \_gnd_net_\,
            in3 => \N__14750\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14747\,
            in2 => \_gnd_net_\,
            in3 => \N__14735\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__32963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14998\,
            in2 => \_gnd_net_\,
            in3 => \N__14984\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14981\,
            in2 => \_gnd_net_\,
            in3 => \N__14969\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14966\,
            in2 => \_gnd_net_\,
            in3 => \N__14954\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14951\,
            in2 => \_gnd_net_\,
            in3 => \N__14939\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14936\,
            in2 => \_gnd_net_\,
            in3 => \N__14924\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14921\,
            in2 => \_gnd_net_\,
            in3 => \N__14909\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14905\,
            in2 => \_gnd_net_\,
            in3 => \N__14891\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14888\,
            in2 => \_gnd_net_\,
            in3 => \N__14876\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__33069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14873\,
            in2 => \_gnd_net_\,
            in3 => \N__14861\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__33059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15191\,
            in2 => \_gnd_net_\,
            in3 => \N__15179\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__33059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15175\,
            in2 => \_gnd_net_\,
            in3 => \N__15161\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__33059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15158\,
            in2 => \_gnd_net_\,
            in3 => \N__15146\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__33059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15142\,
            in2 => \_gnd_net_\,
            in3 => \N__15128\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__33059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15125\,
            in2 => \_gnd_net_\,
            in3 => \N__15113\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__33059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15107\,
            in2 => \_gnd_net_\,
            in3 => \N__15110\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__15087\,
            in1 => \N__15063\,
            in2 => \N__15043\,
            in3 => \N__15020\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15005\,
            in2 => \N__16430\,
            in3 => \N__25100\,
            lcout => \POWERLED.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15290\,
            in2 => \N__15281\,
            in3 => \N__25148\,
            lcout => \POWERLED.N_4527_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_0\,
            carryout => \POWERLED.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15272\,
            in2 => \N__16469\,
            in3 => \N__19334\,
            lcout => \POWERLED.N_4528_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_1\,
            carryout => \POWERLED.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15254\,
            in2 => \N__15266\,
            in3 => \N__19295\,
            lcout => \POWERLED.N_4529_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_2\,
            carryout => \POWERLED.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15233\,
            in2 => \N__15248\,
            in3 => \N__19256\,
            lcout => \POWERLED.N_4530_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_3\,
            carryout => \POWERLED.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20741\,
            in1 => \N__15227\,
            in2 => \N__15476\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4531_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_4\,
            carryout => \POWERLED.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20651\,
            in1 => \N__15209\,
            in2 => \N__15221\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4532_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_5\,
            carryout => \POWERLED.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15203\,
            in2 => \N__15641\,
            in3 => \N__19553\,
            lcout => \POWERLED.N_4533_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_6\,
            carryout => \POWERLED.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19514\,
            in1 => \N__15197\,
            in2 => \N__15692\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4534_i\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19595\,
            in1 => \N__15347\,
            in2 => \N__15494\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4535_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_8\,
            carryout => \POWERLED.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19469\,
            in1 => \N__15341\,
            in2 => \N__21851\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4536_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_9\,
            carryout => \POWERLED.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19418\,
            in1 => \N__15335\,
            in2 => \N__15461\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4537_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_10\,
            carryout => \POWERLED.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21998\,
            in1 => \N__15329\,
            in2 => \N__15626\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4538_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_11\,
            carryout => \POWERLED.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15356\,
            in2 => \N__15323\,
            in3 => \N__20486\,
            lcout => \POWERLED.N_4539_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_12\,
            carryout => \POWERLED.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20696\,
            in1 => \N__15782\,
            in2 => \N__15314\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4540_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_13\,
            carryout => \POWERLED.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19655\,
            in1 => \N__15614\,
            in2 => \N__15305\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4541_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_14\,
            carryout => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15293\,
            lcout => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16526\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15533\,
            lcout => \POWERLED.un85_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15438\,
            lcout => \POWERLED.un85_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16826\,
            lcout => \POWERLED.un85_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_SUSn_RNIN4K9_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16256\,
            lcout => v33a_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15431\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17981\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20111\,
            lcout => \POWERLED.un85_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15596\,
            lcout => \POWERLED.un85_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17914\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23379\,
            lcout => \POWERLED.N_2215_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15669\,
            lcout => \POWERLED.un85_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18395\,
            lcout => \POWERLED.un85_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18314\,
            lcout => \POWERLED.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18104\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17884\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15590\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20204\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__15773\,
            in1 => \N__29276\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18124\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15749\,
            in2 => \N__15844\,
            in3 => \N__15731\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15840\,
            in2 => \N__16658\,
            in3 => \N__15722\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16815\,
            in2 => \N__16643\,
            in3 => \N__15713\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16865\,
            in2 => \N__16822\,
            in3 => \N__15704\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21880\,
            in1 => \N__16853\,
            in2 => \N__15845\,
            in3 => \N__15695\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16841\,
            in2 => \_gnd_net_\,
            in3 => \N__15848\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16814\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18160\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18128\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15788\,
            in1 => \N__16046\,
            in2 => \_gnd_net_\,
            in3 => \N__31959\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__15910\,
            in1 => \N__16117\,
            in2 => \N__15797\,
            in3 => \N__15953\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.m4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI09KEQ_0_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15887\,
            in2 => \N__15794\,
            in3 => \N__31960\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__16068\,
            in1 => \N__17481\,
            in2 => \N__15791\,
            in3 => \N__17393\,
            lcout => \PCH_PWRGD.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32843\,
            ce => \N__31764\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIFF124_9_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17030\,
            in1 => \N__17234\,
            in2 => \_gnd_net_\,
            in3 => \N__18692\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => \PCH_PWRGD.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIDC024_0_8_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__18693\,
            in1 => \N__15938\,
            in2 => \N__15923\,
            in3 => \N__15920\,
            lcout => \PCH_PWRGD.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__16067\,
            in1 => \N__16116\,
            in2 => \N__15911\,
            in3 => \N__15952\,
            lcout => \PCH_PWRGD.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32843\,
            ce => \N__31764\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI3TQ14_0_3_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__15881\,
            in1 => \N__15869\,
            in2 => \N__18713\,
            in3 => \N__16909\,
            lcout => \PCH_PWRGD.un12_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNISRGB1_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__16927\,
            in1 => \N__16943\,
            in2 => \N__17478\,
            in3 => \N__17380\,
            lcout => \PCH_PWRGD.count_rst_11\,
            ltout => \PCH_PWRGD.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI3TQ14_3_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18680\,
            in2 => \N__15875\,
            in3 => \N__15868\,
            lcout => \PCH_PWRGD.un2_count_1_axb_3\,
            ltout => \PCH_PWRGD.un2_count_1_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_3_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__17448\,
            in1 => \N__16931\,
            in2 => \N__15872\,
            in3 => \N__17384\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32769\,
            ce => \N__18717\,
            sr => \N__18913\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNITTHB1_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17381\,
            in1 => \N__17446\,
            in2 => \N__16913\,
            in3 => \N__16891\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI50S14_4_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18681\,
            in1 => \_gnd_net_\,
            in2 => \N__15860\,
            in3 => \N__15854\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => \PCH_PWRGD.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17382\,
            in1 => \N__17449\,
            in2 => \N__15857\,
            in3 => \N__16892\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32769\,
            ce => \N__18717\,
            sr => \N__18913\
        );

    \PCH_PWRGD.count_0_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17447\,
            in1 => \N__16990\,
            in2 => \_gnd_net_\,
            in3 => \N__17383\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32769\,
            ce => \N__18717\,
            sr => \N__18913\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNIBHA61_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__17377\,
            in1 => \N__17080\,
            in2 => \N__17480\,
            in3 => \N__17093\,
            lcout => \PCH_PWRGD.count_rst_3\,
            ltout => \PCH_PWRGD.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI14454_11_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15982\,
            in1 => \_gnd_net_\,
            in2 => \N__15998\,
            in3 => \N__18702\,
            lcout => \PCH_PWRGD.un2_count_1_axb_11\,
            ltout => \PCH_PWRGD.un2_count_1_axb_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_11_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17378\,
            in1 => \N__17459\,
            in2 => \N__15995\,
            in3 => \N__17081\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32985\,
            ce => \N__18719\,
            sr => \N__18937\
        );

    \PCH_PWRGD.count_RNI14454_0_11_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__15992\,
            in1 => \N__17021\,
            in2 => \N__15986\,
            in3 => \N__18703\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOGSAG_3_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15974\,
            in1 => \N__16760\,
            in2 => \N__15968\,
            in3 => \N__15965\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIVBLSO_2_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18797\,
            in1 => \N__16034\,
            in2 => \N__15956\,
            in3 => \N__18521\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => \PCH_PWRGD.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIVBLSO_0_2_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15941\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2\,
            ltout => \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__16118\,
            in1 => \N__16079\,
            in2 => \N__16049\,
            in3 => \N__17379\,
            lcout => \PCH_PWRGD.curr_state_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_14_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17527\,
            lcout => \PCH_PWRGD.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32819\,
            ce => \N__18666\,
            sr => \N__18927\
        );

    \PCH_PWRGD.count_RNI9G854_15_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16016\,
            in1 => \N__17500\,
            in2 => \_gnd_net_\,
            in3 => \N__18665\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => \PCH_PWRGD.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI_15_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16989\,
            in1 => \N__17540\,
            in2 => \N__16037\,
            in3 => \N__17066\,
            lcout => \PCH_PWRGD.un12_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNILIKA4_14_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__16028\,
            in1 => \_gnd_net_\,
            in2 => \N__17528\,
            in3 => \N__18664\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI5A654_13_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16022\,
            in1 => \N__18663\,
            in2 => \_gnd_net_\,
            in3 => \N__17053\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_13_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32819\,
            ce => \N__18666\,
            sr => \N__18927\
        );

    \PCH_PWRGD.count_15_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17501\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32819\,
            ce => \N__18666\,
            sr => \N__18927\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30415\,
            in1 => \N__17642\,
            in2 => \_gnd_net_\,
            in3 => \N__16185\,
            lcout => \RSMRST_PWRGD_RSMRSTn_2_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33085\,
            ce => \N__29415\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_0_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__30418\,
            in1 => \N__17640\,
            in2 => \_gnd_net_\,
            in3 => \N__16182\,
            lcout => \RSMRST_PWRGD.N_256_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000010"
        )
    port map (
            in0 => \N__16184\,
            in1 => \N__17222\,
            in2 => \N__17650\,
            in3 => \N__30416\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33085\,
            ce => \N__29415\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_o2_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30417\,
            in1 => \N__17221\,
            in2 => \_gnd_net_\,
            in3 => \N__16183\,
            lcout => \N_187\,
            ltout => \N_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__17646\,
            in1 => \_gnd_net_\,
            in2 => \N__16310\,
            in3 => \N__16187\,
            lcout => \RSMRST_PWRGD_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33085\,
            ce => \N__29415\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16296\,
            in1 => \N__16265\,
            in2 => \N__16255\,
            in3 => \N__16219\,
            lcout => rsmrst_pwrgd_signal,
            ltout => \rsmrst_pwrgd_signal_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__17641\,
            in1 => \_gnd_net_\,
            in2 => \N__16190\,
            in3 => \N__16186\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33085\,
            ce => \N__29415\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_4_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19229\,
            lcout => \POWERLED.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32964\,
            ce => \N__31765\,
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16163\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16133\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16400\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16388\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16376\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16364\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16355\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16340\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.slp_s3n_signal_i_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__22387\,
            in1 => \N__22489\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26933\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16418\,
            in2 => \N__16450\,
            in3 => \N__16514\,
            lcout => \G_2121\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16446\,
            in2 => \N__16412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16515\,
            in2 => \N__16568\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16556\,
            in2 => \N__16522\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16547\,
            in2 => \N__16451\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__16538\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16433\,
            lcout => \POWERLED.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26490\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26491\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16479\,
            in2 => \N__16493\,
            in3 => \N__16403\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17840\,
            in2 => \N__16484\,
            in3 => \N__16559\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18023\,
            in2 => \N__17822\,
            in3 => \N__16550\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17798\,
            in2 => \N__18029\,
            in3 => \N__16541\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16513\,
            in1 => \N__16483\,
            in2 => \N__17747\,
            in3 => \N__16532\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16529\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26266\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18027\,
            lcout => \POWERLED.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17992\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19828\,
            lcout => \POWERLED.mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18061\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__19903\,
            in1 => \N__25817\,
            in2 => \N__19928\,
            in3 => \N__21068\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33113\,
            ce => 'H',
            sr => \N__22884\
        );

    \POWERLED.dutycycle_12_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__23492\,
            in1 => \N__25816\,
            in2 => \N__23512\,
            in3 => \N__23642\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33113\,
            ce => 'H',
            sr => \N__22884\
        );

    \POWERLED.dutycycle_RNI_2_14_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__19753\,
            in1 => \N__23470\,
            in2 => \N__21215\,
            in3 => \N__23045\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_9_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24280\,
            in1 => \N__23264\,
            in2 => \N__16586\,
            in3 => \N__22640\,
            lcout => \POWERLED.N_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_11_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23469\,
            in2 => \_gnd_net_\,
            in3 => \N__24279\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_46_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_14_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__22649\,
            in1 => \N__21211\,
            in2 => \N__16583\,
            in3 => \N__20264\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18062\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16580\,
            in2 => \_gnd_net_\,
            in3 => \N__16571\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20051\,
            in2 => \N__18197\,
            in3 => \N__16628\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27461\,
            in2 => \N__20027\,
            in3 => \N__16625\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27469\,
            in2 => \N__20003\,
            in3 => \N__16622\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16725\,
            in1 => \N__26108\,
            in2 => \N__26081\,
            in3 => \N__16619\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25411\,
            in2 => \N__25432\,
            in3 => \N__16616\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => \POWERLED.mult1_un54_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16613\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18188\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16610\,
            in2 => \N__16693\,
            in3 => \N__16601\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16689\,
            in2 => \N__16598\,
            in3 => \N__16589\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16739\,
            in2 => \N__16730\,
            in3 => \N__16733\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16729\,
            in2 => \N__16712\,
            in3 => \N__16703\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18305\,
            in1 => \N__16700\,
            in2 => \N__16694\,
            in3 => \N__16676\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16673\,
            in3 => \N__16664\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => \POWERLED.mult1_un61_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16661\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18100\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18209\,
            in2 => \N__16789\,
            in3 => \N__16646\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16785\,
            in2 => \N__18452\,
            in3 => \N__16631\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18383\,
            in2 => \N__18440\,
            in3 => \N__16856\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18428\,
            in2 => \N__18391\,
            in3 => \N__16844\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16813\,
            in1 => \N__18419\,
            in2 => \N__16790\,
            in3 => \N__16832\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18410\,
            in3 => \N__16829\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18382\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI73T14_5_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16768\,
            in1 => \N__16747\,
            in2 => \_gnd_net_\,
            in3 => \N__18690\,
            lcout => \PCH_PWRGD.un2_count_1_axb_5\,
            ltout => \PCH_PWRGD.un2_count_1_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_5_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__17487\,
            in1 => \N__17192\,
            in2 => \N__16772\,
            in3 => \N__17388\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32693\,
            ce => \N__18697\,
            sr => \N__18938\
        );

    \PCH_PWRGD.count_RNI73T14_0_5_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__16769\,
            in1 => \N__17176\,
            in2 => \N__18715\,
            in3 => \N__16748\,
            lcout => \PCH_PWRGD.un12_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNIUVIB1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__17485\,
            in1 => \N__17191\,
            in2 => \N__16880\,
            in3 => \N__17385\,
            lcout => \PCH_PWRGD.count_rst_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNI04LB1_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17386\,
            in1 => \N__17486\,
            in2 => \N__17162\,
            in3 => \N__17177\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIB9V14_7_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18691\,
            in1 => \_gnd_net_\,
            in2 => \N__17042\,
            in3 => \N__17036\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => \PCH_PWRGD.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_7_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17387\,
            in1 => \N__17488\,
            in2 => \N__17039\,
            in3 => \N__17161\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32693\,
            ce => \N__18697\,
            sr => \N__18938\
        );

    \PCH_PWRGD.count_9_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__17392\,
            in1 => \N__17249\,
            in2 => \N__17492\,
            in3 => \N__17265\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32693\,
            ce => \N__18697\,
            sr => \N__18938\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17020\,
            in2 => \N__16991\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSC_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18944\,
            in2 => \_gnd_net_\,
            in3 => \N__16946\,
            lcout => \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSCZ0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16942\,
            in2 => \_gnd_net_\,
            in3 => \N__16916\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16908\,
            in2 => \_gnd_net_\,
            in3 => \N__16883\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16876\,
            in2 => \_gnd_net_\,
            in3 => \N__17183\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNIV1KB1_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17389\,
            in1 => \N__18814\,
            in2 => \_gnd_net_\,
            in3 => \N__17180\,
            lcout => \PCH_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17175\,
            in2 => \_gnd_net_\,
            in3 => \N__17147\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17144\,
            in2 => \_gnd_net_\,
            in3 => \N__17102\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17266\,
            in2 => \_gnd_net_\,
            in3 => \N__17099\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNI3AOB1_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17394\,
            in1 => \N__17660\,
            in2 => \_gnd_net_\,
            in3 => \N__17096\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17092\,
            in2 => \_gnd_net_\,
            in3 => \N__17072\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNICJB61_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17395\,
            in1 => \N__18764\,
            in2 => \_gnd_net_\,
            in3 => \N__17069\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNIDLC61_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17391\,
            in1 => \N__17065\,
            in2 => \_gnd_net_\,
            in3 => \N__17045\,
            lcout => \PCH_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNISSQB1_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18926\,
            in1 => \N__17539\,
            in2 => \_gnd_net_\,
            in3 => \N__17516\,
            lcout => \PCH_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNIFPE61_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__17513\,
            in1 => \N__17396\,
            in2 => \_gnd_net_\,
            in3 => \N__17504\,
            lcout => \PCH_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNI28NB1_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__17479\,
            in1 => \N__17390\,
            in2 => \N__17270\,
            in3 => \N__17245\,
            lcout => \PCH_PWRGD.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI9RLK1_3_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19021\,
            in1 => \N__19036\,
            in2 => \N__19070\,
            in3 => \N__19006\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIR8OP4_10_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17198\,
            in1 => \N__17204\,
            in2 => \N__17225\,
            in3 => \N__17210\,
            lcout => \RSMRST_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19156\,
            in1 => \N__19138\,
            in2 => \N__19193\,
            in3 => \N__19207\,
            lcout => \RSMRST_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIBFU91_13_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19084\,
            in1 => \N__18487\,
            in2 => \N__19175\,
            in3 => \N__18475\,
            lcout => \RSMRST_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIQUU91_10_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19051\,
            in1 => \N__18973\,
            in2 => \N__18992\,
            in3 => \N__18958\,
            lcout => \RSMRST_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI1KAM_0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31800\,
            in2 => \_gnd_net_\,
            in3 => \N__25213\,
            lcout => \POWERLED.g0_i_o3_0\,
            ltout => \POWERLED.g0_i_o3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__17596\,
            in1 => \N__25248\,
            in2 => \N__17600\,
            in3 => \N__19342\,
            lcout => \POWERLED.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32900\,
            ce => 'H',
            sr => \N__19373\
        );

    \POWERLED.pwm_out_RNIB7P12_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001110"
        )
    port map (
            in0 => \N__25249\,
            in1 => \N__17597\,
            in2 => \N__19346\,
            in3 => \N__17588\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__25214\,
            in1 => \N__25182\,
            in2 => \_gnd_net_\,
            in3 => \N__25247\,
            lcout => OPEN,
            ltout => \POWERLED.curr_state_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI2P6L_0_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25163\,
            in2 => \N__17564\,
            in3 => \N__31967\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => \POWERLED.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIE5D5_0_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__31968\,
            in1 => \_gnd_net_\,
            in2 => \N__17561\,
            in3 => \N__25181\,
            lcout => \POWERLED.count_0_sqmuxa_i\,
            ltout => \POWERLED.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_0_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__25084\,
            in1 => \_gnd_net_\,
            in2 => \N__17558\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.count_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIFAFE_0_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31969\,
            in1 => \_gnd_net_\,
            in2 => \N__17555\,
            in3 => \N__24965\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI96U14_6_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18688\,
            in1 => \N__17666\,
            in2 => \_gnd_net_\,
            in3 => \N__17551\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_6_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32989\,
            ce => \N__18718\,
            sr => \N__18928\
        );

    \PCH_PWRGD.count_RNIORHA4_10_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18689\,
            in1 => \N__18736\,
            in2 => \_gnd_net_\,
            in3 => \N__18757\,
            lcout => \PCH_PWRGD.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_10_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18758\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32989\,
            ce => \N__18718\,
            sr => \N__18928\
        );

    \POWERLED.G_11_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__17651\,
            in1 => \N__17621\,
            in2 => \_gnd_net_\,
            in3 => \N__29539\,
            lcout => \G_11\,
            ltout => \G_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29540\,
            in1 => \_gnd_net_\,
            in2 => \N__17615\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.N_27_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_209_i_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27890\,
            in1 => \N__28056\,
            in2 => \_gnd_net_\,
            in3 => \N__31993\,
            lcout => \POWERLED.N_209_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI0LHN_4_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31992\,
            in1 => \N__17612\,
            in2 => \_gnd_net_\,
            in3 => \N__19222\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIJKSP_10_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__17858\,
            in1 => \_gnd_net_\,
            in2 => \N__19438\,
            in3 => \N__31997\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNISEFN_2_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17606\,
            in1 => \N__31994\,
            in2 => \_gnd_net_\,
            in3 => \N__19306\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19310\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33016\,
            ce => \N__31768\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNISF4O_11_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__17690\,
            in1 => \_gnd_net_\,
            in2 => \N__19394\,
            in3 => \N__31996\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_11_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19393\,
            lcout => \POWERLED.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33016\,
            ce => \N__31768\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUHGN_3_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17684\,
            in1 => \N__31995\,
            in2 => \_gnd_net_\,
            in3 => \N__19267\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_3_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19271\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33016\,
            ce => \N__31768\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI4S8O_15_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17678\,
            in1 => \N__31989\,
            in2 => \_gnd_net_\,
            in3 => \N__19621\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_15_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19625\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33070\,
            ce => \N__31770\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI6UKN_7_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17672\,
            in1 => \N__31990\,
            in2 => \_gnd_net_\,
            in3 => \N__19525\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_7_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19529\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33070\,
            ce => \N__31770\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI81MN_8_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17864\,
            in1 => \N__31991\,
            in2 => \_gnd_net_\,
            in3 => \N__19483\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_8_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19487\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33070\,
            ce => \N__31770\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_9_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19607\,
            lcout => \POWERLED.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33070\,
            ce => \N__31770\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_10_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19439\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33078\,
            ce => \N__31769\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26241\,
            in3 => \N__26739\,
            lcout => \POWERLED.N_337\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17727\,
            in2 => \N__17849\,
            in3 => \N__17834\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17831\,
            in2 => \N__17732\,
            in3 => \N__17810\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17807\,
            in2 => \N__17789\,
            in3 => \N__17792\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17788\,
            in2 => \N__17759\,
            in3 => \N__17735\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18022\,
            in1 => \N__17731\,
            in2 => \N__17711\,
            in3 => \N__17693\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18041\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18032\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22072\,
            lcout => \SUSWARN_N_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_3_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26695\,
            in2 => \N__26942\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26937\,
            in2 => \N__20951\,
            in3 => \N__17960\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26278\,
            in2 => \N__27194\,
            in3 => \N__17939\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26804\,
            in2 => \N__26287\,
            in3 => \N__17918\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20963\,
            in2 => \N__22543\,
            in3 => \N__17891\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26194\,
            in2 => \N__23153\,
            in3 => \N__17867\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_4_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20915\,
            in2 => \N__26198\,
            in3 => \N__18131\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24263\,
            in2 => \N__20933\,
            in3 => \N__18107\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23471\,
            in2 => \N__21035\,
            in3 => \N__18083\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24175\,
            in2 => \N__20297\,
            in3 => \N__18080\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_8_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23036\,
            in2 => \N__19859\,
            in3 => \N__18077\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_9_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18074\,
            in2 => \N__21200\,
            in3 => \N__18068\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_10\,
            carryout => \POWERLED.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23318\,
            in2 => \N__23378\,
            in3 => \N__18065\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_11\,
            carryout => \POWERLED.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21257\,
            in2 => \N__23044\,
            in3 => \N__18047\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_12\,
            carryout => \POWERLED.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21189\,
            in2 => \N__21146\,
            in3 => \N__18044\,
            lcout => \POWERLED.mult1_un47_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_13\,
            carryout => \POWERLED.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23366\,
            in2 => \N__19763\,
            in3 => \N__18218\,
            lcout => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_14\,
            carryout => \POWERLED.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23367\,
            in2 => \N__19805\,
            in3 => \N__18215\,
            lcout => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18212\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18232\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__20046\,
            in1 => \N__20047\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__19952\,
            in1 => \_gnd_net_\,
            in2 => \N__18173\,
            in3 => \N__19974\,
            lcout => \POWERLED.mult1_un40_sum_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19879\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18187\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18169\,
            in2 => \N__19976\,
            in3 => \N__19951\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20074\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18344\,
            in2 => \N__18268\,
            in3 => \N__18338\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2_c\,
            carryout => \POWERLED.mult1_un68_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18264\,
            in2 => \N__18335\,
            in3 => \N__18326\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3_c\,
            carryout => \POWERLED.mult1_un68_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18323\,
            in2 => \N__18313\,
            in3 => \N__18317\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4_c\,
            carryout => \POWERLED.mult1_un68_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18309\,
            in2 => \N__18287\,
            in3 => \N__18278\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5_c\,
            carryout => \POWERLED.mult1_un68_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20195\,
            in1 => \N__18275\,
            in2 => \N__18269\,
            in3 => \N__18251\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6_c\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18248\,
            in3 => \N__18239\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => \POWERLED.mult1_un68_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18236\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18233\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18461\,
            in2 => \N__18361\,
            in3 => \N__18443\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18357\,
            in2 => \N__20252\,
            in3 => \N__18431\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20099\,
            in2 => \N__20231\,
            in3 => \N__18422\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20213\,
            in2 => \N__20107\,
            in3 => \N__18413\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18387\,
            in1 => \N__20168\,
            in2 => \N__18362\,
            in3 => \N__18401\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20135\,
            in3 => \N__18398\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20098\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_12_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18779\,
            lcout => \PCH_PWRGD.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32489\,
            ce => \N__18716\,
            sr => \N__18936\
        );

    \PCH_PWRGD.count_2_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__18841\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18882\,
            lcout => \PCH_PWRGD.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32686\,
            ce => \N__18714\,
            sr => \N__18935\
        );

    \PCH_PWRGD.count_RNIFV674_2_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__18677\,
            in1 => \N__18829\,
            in2 => \N__18845\,
            in3 => \N__18880\,
            lcout => \PCH_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__18881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18840\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIFV674_0_2_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__18679\,
            in1 => \N__18830\,
            in2 => \N__18821\,
            in3 => \N__18818\,
            lcout => \PCH_PWRGD.un12_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI37554_12_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18678\,
            in1 => \N__18785\,
            in2 => \_gnd_net_\,
            in3 => \N__18775\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => \PCH_PWRGD.countZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIORHA4_0_10_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__18756\,
            in1 => \N__18740\,
            in2 => \N__18722\,
            in3 => \N__18676\,
            lcout => \PCH_PWRGD.un12_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29549\,
            in1 => \N__18488\,
            in2 => \N__18509\,
            in3 => \N__18508\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_1_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29543\,
            in1 => \N__18476\,
            in2 => \_gnd_net_\,
            in3 => \N__18464\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_2_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29550\,
            in1 => \N__19085\,
            in2 => \_gnd_net_\,
            in3 => \N__19073\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_3_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29544\,
            in1 => \N__19069\,
            in2 => \_gnd_net_\,
            in3 => \N__19055\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_4_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29551\,
            in1 => \N__19052\,
            in2 => \_gnd_net_\,
            in3 => \N__19040\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_5_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29545\,
            in1 => \N__19037\,
            in2 => \_gnd_net_\,
            in3 => \N__19025\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_6_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29552\,
            in1 => \N__19022\,
            in2 => \_gnd_net_\,
            in3 => \N__19010\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_7_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29546\,
            in1 => \N__19007\,
            in2 => \_gnd_net_\,
            in3 => \N__18995\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__32634\,
            ce => 'H',
            sr => \N__19114\
        );

    \RSMRST_PWRGD.count_8_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29567\,
            in1 => \N__18991\,
            in2 => \_gnd_net_\,
            in3 => \N__18977\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__32887\,
            ce => 'H',
            sr => \N__19115\
        );

    \RSMRST_PWRGD.count_9_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29563\,
            in1 => \N__18974\,
            in2 => \_gnd_net_\,
            in3 => \N__18962\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__32887\,
            ce => 'H',
            sr => \N__19115\
        );

    \RSMRST_PWRGD.count_10_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29564\,
            in1 => \N__18959\,
            in2 => \_gnd_net_\,
            in3 => \N__18947\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__32887\,
            ce => 'H',
            sr => \N__19115\
        );

    \RSMRST_PWRGD.count_11_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29561\,
            in1 => \N__19208\,
            in2 => \_gnd_net_\,
            in3 => \N__19196\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__32887\,
            ce => 'H',
            sr => \N__19115\
        );

    \RSMRST_PWRGD.count_12_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29565\,
            in1 => \N__19192\,
            in2 => \_gnd_net_\,
            in3 => \N__19178\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__32887\,
            ce => 'H',
            sr => \N__19115\
        );

    \RSMRST_PWRGD.count_13_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29562\,
            in1 => \N__19174\,
            in2 => \_gnd_net_\,
            in3 => \N__19160\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__32887\,
            ce => 'H',
            sr => \N__19115\
        );

    \RSMRST_PWRGD.count_14_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29566\,
            in1 => \N__19157\,
            in2 => \_gnd_net_\,
            in3 => \N__19145\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__32887\,
            ce => 'H',
            sr => \N__19115\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27453\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19139\,
            in2 => \_gnd_net_\,
            in3 => \N__19142\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32899\,
            ce => \N__19127\,
            sr => \N__19104\
        );

    \POWERLED.count_RNI_2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19252\,
            in3 => \N__19326\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_3_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__20640\,
            in1 => \N__20730\,
            in2 => \N__19088\,
            in3 => \N__19287\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlt15_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_7_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19513\,
            in1 => \N__19548\,
            in2 => \N__19376\,
            in3 => \N__19591\,
            lcout => \POWERLED.un79_clk_100khzlto15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31998\,
            in1 => \N__25218\,
            in2 => \_gnd_net_\,
            in3 => \N__25183\,
            lcout => \POWERLED.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_10_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19410\,
            in1 => \N__20475\,
            in2 => \N__19464\,
            in3 => \N__21994\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_15_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20685\,
            in1 => \N__19358\,
            in2 => \N__19352\,
            in3 => \N__19650\,
            lcout => \POWERLED.count_RNIZ0Z_15\,
            ltout => \POWERLED.count_RNIZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIFPNR_0_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__25219\,
            in1 => \N__31799\,
            in2 => \N__19349\,
            in3 => \N__31999\,
            lcout => \POWERLED.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25140\,
            in2 => \N__25098\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \POWERLED.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_RNIB209_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25030\,
            in1 => \N__19327\,
            in2 => \_gnd_net_\,
            in3 => \N__19298\,
            lcout => \POWERLED.un1_count_cry_1_c_RNIBZ0Z209\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_1\,
            carryout => \POWERLED.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_2_c_RNIC419_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25036\,
            in1 => \N__19288\,
            in2 => \_gnd_net_\,
            in3 => \N__19259\,
            lcout => \POWERLED.un1_count_cry_2_c_RNICZ0Z419\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_2\,
            carryout => \POWERLED.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_3_c_RNID629_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25031\,
            in1 => \N__19248\,
            in2 => \_gnd_net_\,
            in3 => \N__19211\,
            lcout => \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_3\,
            carryout => \POWERLED.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNIE839_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25034\,
            in1 => \N__20731\,
            in2 => \_gnd_net_\,
            in3 => \N__19559\,
            lcout => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_4\,
            carryout => \POWERLED.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNIFA49_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25033\,
            in1 => \N__20641\,
            in2 => \_gnd_net_\,
            in3 => \N__19556\,
            lcout => \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_5\,
            carryout => \POWERLED.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_6_c_RNIGC59_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25035\,
            in1 => \N__19549\,
            in2 => \_gnd_net_\,
            in3 => \N__19517\,
            lcout => \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_6\,
            carryout => \POWERLED.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_7_c_RNIHE69_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25032\,
            in1 => \N__19506\,
            in2 => \_gnd_net_\,
            in3 => \N__19475\,
            lcout => \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_7\,
            carryout => \POWERLED.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_8_c_RNIIG79_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25041\,
            in1 => \N__19587\,
            in2 => \_gnd_net_\,
            in3 => \N__19472\,
            lcout => \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79\,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => \POWERLED.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_9_c_RNIJI89_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25038\,
            in1 => \_gnd_net_\,
            in2 => \N__19465\,
            in3 => \N__19421\,
            lcout => \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_9\,
            carryout => \POWERLED.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25043\,
            in1 => \N__19411\,
            in2 => \_gnd_net_\,
            in3 => \N__19382\,
            lcout => \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_10\,
            carryout => \POWERLED.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_11_c_RNISEH7_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25037\,
            in1 => \N__21990\,
            in2 => \_gnd_net_\,
            in3 => \N__19379\,
            lcout => \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_11\,
            carryout => \POWERLED.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_12_c_RNITGI7_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25042\,
            in1 => \N__20476\,
            in2 => \_gnd_net_\,
            in3 => \N__19661\,
            lcout => \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_12\,
            carryout => \POWERLED.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25039\,
            in1 => \N__20686\,
            in2 => \_gnd_net_\,
            in3 => \N__19658\,
            lcout => \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_13\,
            carryout => \POWERLED.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__19651\,
            in1 => \N__25040\,
            in2 => \_gnd_net_\,
            in3 => \N__19628\,
            lcout => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIA4NN_9_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19613\,
            in1 => \N__31988\,
            in2 => \_gnd_net_\,
            in3 => \N__19606\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI496F5_2_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__23884\,
            in1 => \N__20870\,
            in2 => \N__21786\,
            in3 => \N__20879\,
            lcout => \POWERLED.dutycycle_eena_1\,
            ltout => \POWERLED.dutycycle_eena_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN2MP8_2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__23778\,
            in1 => \N__19693\,
            in2 => \N__19568\,
            in3 => \N__20413\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNINQPO7_1_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__19711\,
            in1 => \N__23777\,
            in2 => \N__20510\,
            in3 => \N__19721\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIP27U5_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111111111"
        )
    port map (
            in0 => \N__30524\,
            in1 => \N__19565\,
            in2 => \N__26941\,
            in3 => \N__23883\,
            lcout => \POWERLED.dutycycle_eena\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIELPT3_1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__30522\,
            in2 => \N__28124\,
            in3 => \N__20878\,
            lcout => \POWERLED.N_108_f0_1\,
            ltout => \POWERLED.N_108_f0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIP27U5_1_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100110111"
        )
    port map (
            in0 => \N__30523\,
            in1 => \N__23882\,
            in2 => \N__19724\,
            in3 => \N__26475\,
            lcout => \POWERLED.dutycycle_eena_0\,
            ltout => \POWERLED.dutycycle_eena_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__19712\,
            in1 => \N__20503\,
            in2 => \N__19715\,
            in3 => \N__23780\,
            lcout => \POWERLED.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33077\,
            ce => 'H',
            sr => \N__22900\
        );

    \POWERLED.dutycycle_2_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0111000011111000"
        )
    port map (
            in0 => \N__23779\,
            in1 => \N__19703\,
            in2 => \N__19697\,
            in3 => \N__20414\,
            lcout => \POWERLED.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33077\,
            ce => 'H',
            sr => \N__22900\
        );

    \POWERLED.func_state_0_sqmuxa_0_o2_x1_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__22484\,
            in1 => \N__24906\,
            in2 => \N__28073\,
            in3 => \N__22068\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_0_sqmuxa_0_o2_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_sqmuxa_0_o2_ns_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27445\,
            in2 => \N__19682\,
            in3 => \N__24857\,
            lcout => \POWERLED.N_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBK1U_0_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20441\,
            in2 => \_gnd_net_\,
            in3 => \N__30550\,
            lcout => OPEN,
            ltout => \POWERLED.g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN3GO3_6_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__19814\,
            in1 => \N__19673\,
            in2 => \N__19679\,
            in3 => \N__26576\,
            lcout => \POWERLED.N_217_N_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIBVNS_0_4_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25758\,
            in2 => \_gnd_net_\,
            in3 => \N__28472\,
            lcout => OPEN,
            ltout => \POWERLED.N_300_N_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI6K332_4_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__28068\,
            in1 => \N__27885\,
            in2 => \N__19676\,
            in3 => \N__27097\,
            lcout => \POWERLED.N_4548_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOBU76_6_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__23893\,
            in1 => \N__19667\,
            in2 => \_gnd_net_\,
            in3 => \N__20396\,
            lcout => \POWERLED.dutycycle_eena_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6RAN_0_1_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__24907\,
            in1 => \N__28072\,
            in2 => \_gnd_net_\,
            in3 => \N__27795\,
            lcout => \POWERLED.N_353_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJ27K7_14_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19781\,
            in1 => \N__25756\,
            in2 => \N__21089\,
            in3 => \N__19790\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => \POWERLED.dutycycleZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19808\,
            in3 => \N__22940\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN3GO3_14_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111101111"
        )
    port map (
            in0 => \N__23298\,
            in1 => \N__24019\,
            in2 => \N__24107\,
            in3 => \N__21182\,
            lcout => OPEN,
            ltout => \POWERLED.N_86_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEB706_14_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23891\,
            in2 => \N__19793\,
            in3 => \N__23804\,
            lcout => \POWERLED.dutycycle_en_11\,
            ltout => \POWERLED.dutycycle_en_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__21088\,
            in1 => \N__19777\,
            in2 => \N__19784\,
            in3 => \N__25757\,
            lcout => \POWERLED.dutycycleZ1Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33090\,
            ce => 'H',
            sr => \N__22878\
        );

    \POWERLED.dutycycle_RNI_1_15_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23380\,
            in2 => \N__21199\,
            in3 => \N__22939\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIN3GO3_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111111"
        )
    port map (
            in0 => \N__23299\,
            in1 => \N__24020\,
            in2 => \N__19754\,
            in3 => \N__24104\,
            lcout => OPEN,
            ltout => \POWERLED.N_84_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIEB706_1_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23892\,
            in2 => \N__19727\,
            in3 => \N__23805\,
            lcout => \POWERLED.dutycycle_en_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__21019\,
            in1 => \N__24387\,
            in2 => \_gnd_net_\,
            in3 => \N__24248\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__21325\,
            in1 => \N__19850\,
            in2 => \N__25821\,
            in3 => \N__21122\,
            lcout => \POWERLED.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32949\,
            ce => 'H',
            sr => \N__22879\
        );

    \POWERLED.dutycycle_RNI_0_13_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24249\,
            in2 => \_gnd_net_\,
            in3 => \N__23021\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_10_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_9_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011010010"
        )
    port map (
            in0 => \N__23256\,
            in1 => \N__24394\,
            in2 => \N__19865\,
            in3 => \N__22969\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19862\,
            in3 => \N__23022\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI45I67_10_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__25797\,
            in1 => \N__19849\,
            in2 => \N__21326\,
            in3 => \N__21121\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => \POWERLED.dutycycleZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_9_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101000100"
        )
    port map (
            in0 => \N__21020\,
            in1 => \N__24388\,
            in2 => \N__19841\,
            in3 => \N__23255\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_4Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_11_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19838\,
            in2 => \N__19832\,
            in3 => \N__23468\,
            lcout => \POWERLED.un1_dutycycle_53_50_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19829\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19985\,
            in3 => \N__20030\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19937\,
            in3 => \N__20015\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27468\,
            in2 => \N__20012\,
            in3 => \N__19991\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19988\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19975\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19970\,
            in2 => \_gnd_net_\,
            in3 => \N__19950\,
            lcout => \POWERLED.mult1_un47_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIL58K7_15_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__19927\,
            in1 => \N__25801\,
            in2 => \N__19904\,
            in3 => \N__21061\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19880\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20057\,
            in2 => \N__20152\,
            in3 => \N__20243\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20148\,
            in2 => \N__20240\,
            in3 => \N__20222\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20219\,
            in2 => \N__20203\,
            in3 => \N__20207\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20199\,
            in2 => \N__20177\,
            in3 => \N__20162\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20103\,
            in1 => \N__20159\,
            in2 => \N__20153\,
            in3 => \N__20126\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20123\,
            in3 => \N__20114\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20078\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_7_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000100"
        )
    port map (
            in0 => \N__20285\,
            in1 => \N__24357\,
            in2 => \N__20276\,
            in3 => \N__23100\,
            lcout => \POWERLED.dutycycle_RNI_11Z0Z_7\,
            ltout => \POWERLED.dutycycle_RNI_11Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_12_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__23230\,
            in1 => \N__24179\,
            in2 => \N__20300\,
            in3 => \N__24344\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_9_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110101"
        )
    port map (
            in0 => \N__26599\,
            in1 => \N__26391\,
            in2 => \N__24386\,
            in3 => \N__23228\,
            lcout => \POWERLED.un1_dutycycle_53_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFO3M8_8_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21286\,
            in1 => \N__21304\,
            in2 => \N__25820\,
            in3 => \N__22672\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => \POWERLED.dutycycleZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__26600\,
            in1 => \_gnd_net_\,
            in2 => \N__20279\,
            in3 => \N__26392\,
            lcout => \POWERLED.un1_dutycycle_53_45_a0_1\,
            ltout => \POWERLED.un1_dutycycle_53_45_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_7_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__24267\,
            in1 => \N__23108\,
            in2 => \N__20267\,
            in3 => \N__24343\,
            lcout => \POWERLED.un1_dutycycle_53_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_7_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011011000"
        )
    port map (
            in0 => \N__26601\,
            in1 => \N__23099\,
            in2 => \N__26405\,
            in3 => \N__24356\,
            lcout => \POWERLED.un1_dutycycle_53_13_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110111111"
        )
    port map (
            in0 => \N__23229\,
            in1 => \N__24342\,
            in2 => \N__23128\,
            in3 => \N__26602\,
            lcout => \POWERLED.un1_dutycycle_53_13_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB5IA5_2_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21386\,
            in1 => \N__21380\,
            in2 => \N__21275\,
            in3 => \N__21392\,
            lcout => \HDA_STRAP.un4_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__21445\,
            in1 => \N__24623\,
            in2 => \N__21578\,
            in3 => \N__21506\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32685\,
            ce => \N__29397\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_1_2_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__21504\,
            in1 => \N__21564\,
            in2 => \_gnd_net_\,
            in3 => \N__21444\,
            lcout => OPEN,
            ltout => \HDA_STRAP.N_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000001100"
        )
    port map (
            in0 => \N__21565\,
            in1 => \N__20374\,
            in2 => \N__20378\,
            in3 => \N__20309\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32685\,
            ce => \N__29397\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__20375\,
            in1 => \N__21503\,
            in2 => \_gnd_net_\,
            in3 => \N__21570\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32685\,
            ce => \N__29397\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_1_0_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110101010"
        )
    port map (
            in0 => \N__20348\,
            in1 => \N__20333\,
            in2 => \N__30586\,
            in3 => \N__21505\,
            lcout => OPEN,
            ltout => \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21569\,
            in2 => \N__20336\,
            in3 => \N__20315\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32685\,
            ce => \N__29397\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_0_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101111"
        )
    port map (
            in0 => \N__21443\,
            in1 => \N__20332\,
            in2 => \N__21523\,
            in3 => \N__30576\,
            lcout => \HDA_STRAP.curr_state_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21499\,
            in2 => \_gnd_net_\,
            in3 => \N__30302\,
            lcout => \HDA_STRAP.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_1_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27778\,
            lcout => \POWERLED.N_341\,
            ltout => \POWERLED.N_341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__29249\,
            in1 => \_gnd_net_\,
            in2 => \N__20303\,
            in3 => \N__25595\,
            lcout => \POWERLED.un1_func_state25_6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__27103\,
            in1 => \N__27777\,
            in2 => \N__20816\,
            in3 => \N__22141\,
            lcout => \POWERLED.func_state_1_m2s2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_1_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25594\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_i_a3_1_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI2AJD2_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__28054\,
            in1 => \N__24778\,
            in2 => \N__20417\,
            in3 => \N__20384\,
            lcout => \POWERLED.N_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0RLE1_1_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__28053\,
            in1 => \N__27876\,
            in2 => \N__22049\,
            in3 => \N__27102\,
            lcout => \POWERLED.N_275_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31885\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26032\,
            lcout => suswarn_n,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJ9IE1_0_11_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__28031\,
            in1 => \N__24779\,
            in2 => \_gnd_net_\,
            in3 => \N__21630\,
            lcout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMJCH1_1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23949\,
            in2 => \_gnd_net_\,
            in3 => \N__28242\,
            lcout => \POWERLED.N_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_6_1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__22190\,
            in1 => \N__22140\,
            in2 => \_gnd_net_\,
            in3 => \N__27775\,
            lcout => OPEN,
            ltout => \POWERLED.g0_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBK1U_1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__21827\,
            in1 => \N__30555\,
            in2 => \N__20399\,
            in3 => \N__29242\,
            lcout => \POWERLED.g0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHL0V1_0_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101110111"
        )
    port map (
            in0 => \N__21914\,
            in1 => \N__20761\,
            in2 => \N__27889\,
            in3 => \N__22230\,
            lcout => \POWERLED.func_state_1_m0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010011"
        )
    port map (
            in0 => \N__27776\,
            in1 => \N__30554\,
            in2 => \N__29250\,
            in3 => \N__20999\,
            lcout => \POWERLED.dutycycle_1_0_iv_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__22474\,
            in1 => \N__24946\,
            in2 => \_gnd_net_\,
            in3 => \N__22384\,
            lcout => \POWERLED.N_326_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMQ0F_1_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__28471\,
            in1 => \N__27740\,
            in2 => \N__24955\,
            in3 => \N__24849\,
            lcout => \POWERLED.func_state_RNIMQ0FZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_0_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22221\,
            lcout => \POWERLED.N_2171_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9TUV2_0_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__21653\,
            in1 => \N__20429\,
            in2 => \N__21644\,
            in3 => \N__21811\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIG5G37_1_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__29231\,
            in1 => \N__21602\,
            in2 => \N__20423\,
            in3 => \N__21608\,
            lcout => \POWERLED.func_state_RNIG5G37Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_1_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__25136\,
            in1 => \N__25046\,
            in2 => \_gnd_net_\,
            in3 => \N__25078\,
            lcout => OPEN,
            ltout => \POWERLED.count_RNI_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGBFE_1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31890\,
            in1 => \_gnd_net_\,
            in2 => \N__20420\,
            in3 => \N__25109\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111010111"
        )
    port map (
            in0 => \N__22385\,
            in1 => \N__22475\,
            in2 => \N__24956\,
            in3 => \N__31889\,
            lcout => \POWERLED.N_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__20585\,
            in1 => \N__20591\,
            in2 => \N__23789\,
            in3 => \N__20570\,
            lcout => \POWERLED.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32776\,
            ce => 'H',
            sr => \N__22903\
        );

    \POWERLED.func_state_RNIBVNS_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__26884\,
            in1 => \N__25869\,
            in2 => \N__22247\,
            in3 => \N__27737\,
            lcout => \POWERLED.dutycycle_1_0_0\,
            ltout => \POWERLED.dutycycle_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJFRN7_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__23758\,
            in1 => \N__20584\,
            in2 => \N__20573\,
            in3 => \N__20569\,
            lcout => \POWERLED.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__22243\,
            in1 => \N__21640\,
            in2 => \_gnd_net_\,
            in3 => \N__27739\,
            lcout => \POWERLED.un1_func_state25_4_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI12UT8_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__23757\,
            in1 => \N__21763\,
            in2 => \N__20555\,
            in3 => \N__20524\,
            lcout => \POWERLED.func_state\,
            ltout => \POWERLED.func_state_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20513\,
            in3 => \N__25865\,
            lcout => \POWERLED.func_state_RNIBVNSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100011111"
        )
    port map (
            in0 => \N__27738\,
            in1 => \N__21011\,
            in2 => \N__25871\,
            in3 => \N__22242\,
            lcout => \POWERLED.dutycycle_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_1_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21639\,
            in2 => \_gnd_net_\,
            in3 => \N__27736\,
            lcout => \POWERLED.func_state_RNI_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI0M6O_13_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31987\,
            in1 => \N__20447\,
            in2 => \_gnd_net_\,
            in3 => \N__20455\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_13_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20459\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32798\,
            ce => \N__31763\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI2OIN_5_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31985\,
            in1 => \N__20702\,
            in2 => \_gnd_net_\,
            in3 => \N__20710\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_5_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20714\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32798\,
            ce => \N__31763\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI2P7O_14_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20657\,
            in1 => \N__32003\,
            in2 => \_gnd_net_\,
            in3 => \N__20665\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_14_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20669\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32798\,
            ce => \N__31763\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI4RJN_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31986\,
            in1 => \N__20612\,
            in2 => \_gnd_net_\,
            in3 => \N__20620\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_6_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20624\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32798\,
            ce => \N__31763\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHV5K7_13_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__20788\,
            in1 => \N__25717\,
            in2 => \N__20600\,
            in3 => \N__21103\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => \POWERLED.dutycycleZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN3GO3_13_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__25718\,
            in1 => \N__24099\,
            in2 => \N__20606\,
            in3 => \N__28449\,
            lcout => OPEN,
            ltout => \POWERLED.N_148_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEB706_13_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__23975\,
            in1 => \N__23948\,
            in2 => \N__20603\,
            in3 => \N__23742\,
            lcout => \POWERLED.dutycycle_en_10\,
            ltout => \POWERLED.dutycycle_en_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__21104\,
            in1 => \N__25722\,
            in2 => \N__20792\,
            in3 => \N__20789\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32794\,
            ce => 'H',
            sr => \N__22880\
        );

    \POWERLED.func_state_RNIOTGO_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__28055\,
            in1 => \N__20780\,
            in2 => \N__28250\,
            in3 => \N__30509\,
            lcout => OPEN,
            ltout => \POWERLED.N_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIES0I2_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__21775\,
            in1 => \N__25723\,
            in2 => \N__20771\,
            in3 => \N__23974\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQF354_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__28207\,
            in1 => \N__20768\,
            in2 => \N__20750\,
            in3 => \N__23741\,
            lcout => \POWERLED.count_clk_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_0_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23297\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.func_state_RNIBVNS_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIBVNS_1_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011101110111"
        )
    port map (
            in0 => \N__28456\,
            in1 => \N__25854\,
            in2 => \N__22172\,
            in3 => \N__22131\,
            lcout => \POWERLED.un1_count_off_1_sqmuxa_8_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25581\,
            in2 => \_gnd_net_\,
            in3 => \N__20803\,
            lcout => \POWERLED.dutycycle_RNI_8Z0Z_0\,
            ltout => \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20747\,
            in3 => \N__22132\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_1_0_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011110111111"
        )
    port map (
            in0 => \N__25900\,
            in1 => \N__25728\,
            in2 => \N__20744\,
            in3 => \N__25582\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_RNIBVNS_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMUFP1_1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__26769\,
            in1 => \N__25901\,
            in2 => \N__20891\,
            in3 => \N__20888\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIES0I2_1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28066\,
            in2 => \N__20882\,
            in3 => \N__30484\,
            lcout => \POWERLED.N_171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILP0F_2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__26240\,
            in1 => \N__27768\,
            in2 => \N__30521\,
            in3 => \N__27092\,
            lcout => \POWERLED.N_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_0_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25727\,
            in2 => \_gnd_net_\,
            in3 => \N__25583\,
            lcout => \POWERLED.func_state_RNIBVNS_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__23740\,
            in1 => \N__20839\,
            in2 => \N__20849\,
            in3 => \N__20828\,
            lcout => \POWERLED.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32948\,
            ce => 'H',
            sr => \N__22905\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI92UT3_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__23904\,
            in1 => \N__25759\,
            in2 => \N__20864\,
            in3 => \N__20978\,
            lcout => \POWERLED.dutycycle_set_0_0\,
            ltout => \POWERLED.dutycycle_set_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM1P2B_6_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__23739\,
            in1 => \N__20840\,
            in2 => \N__20831\,
            in3 => \N__20827\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => \POWERLED.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__26921\,
            in1 => \_gnd_net_\,
            in2 => \N__20819\,
            in3 => \N__26456\,
            lcout => \POWERLED.N_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__26922\,
            in2 => \N__26184\,
            in3 => \N__26554\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__26923\,
            in1 => \N__26577\,
            in2 => \N__26750\,
            in3 => \N__26458\,
            lcout => \POWERLED.N_392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_3_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__26455\,
            in1 => \N__26682\,
            in2 => \_gnd_net_\,
            in3 => \N__26555\,
            lcout => OPEN,
            ltout => \POWERLED.d_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_5_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__26165\,
            in1 => \N__22547\,
            in2 => \N__20966\,
            in3 => \N__26504\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26389\,
            in1 => \N__26932\,
            in2 => \_gnd_net_\,
            in3 => \N__26462\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001000"
        )
    port map (
            in0 => \N__23131\,
            in1 => \N__26388\,
            in2 => \N__24424\,
            in3 => \N__26677\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_3\,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_9_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__26565\,
            in1 => \_gnd_net_\,
            in2 => \N__20939\,
            in3 => \N__23258\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_7_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__23132\,
            in1 => \N__26568\,
            in2 => \N__20936\,
            in3 => \N__24264\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26567\,
            in1 => \N__20921\,
            in2 => \N__26190\,
            in3 => \N__23259\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_9_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001010"
        )
    port map (
            in0 => \N__23257\,
            in1 => \N__26566\,
            in2 => \N__20906\,
            in3 => \N__22505\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_13_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_11_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \N__23467\,
            in1 => \N__22511\,
            in2 => \N__21050\,
            in3 => \N__21047\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_7_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100010111"
        )
    port map (
            in0 => \N__23130\,
            in1 => \N__26387\,
            in2 => \N__24423\,
            in3 => \N__26564\,
            lcout => \POWERLED.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26938\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27019\,
            in2 => \N__26482\,
            in3 => \N__21002\,
            lcout => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26265\,
            in2 => \N__27053\,
            in3 => \N__20990\,
            lcout => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_1\,
            carryout => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27017\,
            in2 => \N__26696\,
            in3 => \N__20987\,
            lcout => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27042\,
            in2 => \N__26358\,
            in3 => \N__20984\,
            lcout => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27018\,
            in2 => \N__26191\,
            in3 => \N__20981\,
            lcout => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26578\,
            in2 => \N__27052\,
            in3 => \N__20969\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27013\,
            in2 => \N__23129\,
            in3 => \N__21131\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27020\,
            in2 => \N__24406\,
            in3 => \N__21128\,
            lcout => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_8_c_RNIMPUT_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25738\,
            in1 => \N__27024\,
            in2 => \N__23254\,
            in3 => \N__21125\,
            lcout => \POWERLED.dutycycle_rst_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_8_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27021\,
            in2 => \N__24265\,
            in3 => \N__21113\,
            lcout => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_9\,
            carryout => \POWERLED.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27025\,
            in2 => \N__23453\,
            in3 => \N__21110\,
            lcout => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_10\,
            carryout => \POWERLED.un1_dutycycle_94_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24152\,
            in2 => \N__27054\,
            in3 => \N__21107\,
            lcout => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_11\,
            carryout => \POWERLED.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27029\,
            in2 => \N__23020\,
            in3 => \N__21092\,
            lcout => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_12\,
            carryout => \POWERLED.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27022\,
            in2 => \N__21204\,
            in3 => \N__21074\,
            lcout => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_13\,
            carryout => \POWERLED.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27023\,
            in1 => \N__23371\,
            in2 => \_gnd_net_\,
            in3 => \N__21071\,
            lcout => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000001111"
        )
    port map (
            in0 => \N__23249\,
            in1 => \N__24268\,
            in2 => \N__23466\,
            in3 => \N__24158\,
            lcout => \POWERLED.g0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_9_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__23811\,
            in1 => \N__21245\,
            in2 => \N__23525\,
            in3 => \N__21232\,
            lcout => \POWERLED.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33050\,
            ce => 'H',
            sr => \N__22902\
        );

    \POWERLED.dutycycle_RNI_6_12_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__23250\,
            in1 => \N__24269\,
            in2 => \N__23162\,
            in3 => \N__24159\,
            lcout => OPEN,
            ltout => \POWERLED.g0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_13_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \N__23040\,
            in1 => \N__24185\,
            in2 => \N__21266\,
            in3 => \N__21263\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI67G18_9_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__21244\,
            in1 => \N__23521\,
            in2 => \N__21233\,
            in3 => \N__23810\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => \POWERLED.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_9_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__23168\,
            in1 => \_gnd_net_\,
            in2 => \N__21221\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.g0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_12_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__23449\,
            in1 => \N__24270\,
            in2 => \N__21218\,
            in3 => \N__24160\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_14_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__21205\,
            in1 => \_gnd_net_\,
            in2 => \N__21149\,
            in3 => \N__23035\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_7_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__21350\,
            in1 => \N__21362\,
            in2 => \N__21371\,
            in3 => \N__25805\,
            lcout => \POWERLED.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33139\,
            ce => 'H',
            sr => \N__22907\
        );

    \POWERLED.count_clk_RNI1J4E2_0_4_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__24009\,
            in1 => \N__23946\,
            in2 => \N__28475\,
            in3 => \N__25734\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_36_and_i_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEB706_7_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__24105\,
            in1 => \N__23809\,
            in2 => \N__21374\,
            in3 => \N__21335\,
            lcout => \POWERLED.dutycycle_RNIEB706Z0Z_7\,
            ltout => \POWERLED.dutycycle_RNIEB706Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN1M47_7_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__21361\,
            in1 => \N__25733\,
            in2 => \N__21353\,
            in3 => \N__21349\,
            lcout => \POWERLED.dutycycleZ1Z_6\,
            ltout => \POWERLED.dutycycleZ1Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_7_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21338\,
            in3 => \N__24008\,
            lcout => \POWERLED.un1_clk_100khz_36_and_i_0_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI1J4E2_4_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__28466\,
            in1 => \N__23945\,
            in2 => \_gnd_net_\,
            in3 => \N__25732\,
            lcout => \POWERLED.dutycycle_eena_3_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN3GO3_10_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__24106\,
            in1 => \N__28470\,
            in2 => \N__25793\,
            in3 => \N__24266\,
            lcout => OPEN,
            ltout => \POWERLED.N_143_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEB706_10_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001100"
        )
    port map (
            in0 => \N__24010\,
            in1 => \N__23812\,
            in2 => \N__21329\,
            in3 => \N__23947\,
            lcout => \POWERLED.dutycycle_en_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__21308\,
            in1 => \N__22673\,
            in2 => \N__21290\,
            in3 => \N__25822\,
            lcout => \POWERLED.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33052\,
            ce => 'H',
            sr => \N__22868\
        );

    \HDA_STRAP.count_RNI5DB61_6_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24484\,
            in1 => \N__24568\,
            in2 => \N__24524\,
            in3 => \N__24460\,
            lcout => \HDA_STRAP.un4_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIBJB61_7_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24439\,
            in1 => \N__24499\,
            in2 => \N__24545\,
            in3 => \N__24709\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI0NIR1_14_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24679\,
            in2 => \N__21395\,
            in3 => \N__24694\,
            lcout => \HDA_STRAP.un4_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI4CB61_17_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__23587\,
            in1 => \N__24664\,
            in2 => \N__23624\,
            in3 => \N__24637\,
            lcout => \HDA_STRAP.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI2L821_2_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23539\,
            in1 => \N__23554\,
            in2 => \N__23573\,
            in3 => \N__24583\,
            lcout => \HDA_STRAP.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIH91A_1_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21522\,
            in2 => \_gnd_net_\,
            in3 => \N__21563\,
            lcout => \HDA_STRAP.curr_state_RNIH91AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__21574\,
            in1 => \N__21508\,
            in2 => \N__24557\,
            in3 => \N__21452\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32748\,
            ce => \N__29396\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__21448\,
            in1 => \N__21577\,
            in2 => \N__21526\,
            in3 => \N__24509\,
            lcout => \HDA_STRAP.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32748\,
            ce => \N__29396\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__21572\,
            in1 => \N__21507\,
            in2 => \N__24473\,
            in3 => \N__21450\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32748\,
            ce => \N__29396\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__21447\,
            in1 => \N__21576\,
            in2 => \N__21525\,
            in3 => \N__24449\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32748\,
            ce => \N__29396\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__21571\,
            in1 => \N__21449\,
            in2 => \N__30310\,
            in3 => \N__21518\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32748\,
            ce => \N__29396\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_0_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__21446\,
            in1 => \N__21575\,
            in2 => \N__21524\,
            in3 => \N__23594\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32748\,
            ce => \N__29396\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011001100"
        )
    port map (
            in0 => \N__21573\,
            in1 => \N__24653\,
            in2 => \N__21527\,
            in3 => \N__21451\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32748\,
            ce => \N__29396\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__24952\,
            in1 => \N__22485\,
            in2 => \N__22040\,
            in3 => \N__22391\,
            lcout => \POWERLED.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_2_0_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22392\,
            in1 => \N__24954\,
            in2 => \N__22490\,
            in3 => \N__25584\,
            lcout => \POWERLED.func_state_RNIBVNS_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6RAN_1_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__24953\,
            in1 => \N__28027\,
            in2 => \_gnd_net_\,
            in3 => \N__27797\,
            lcout => \POWERLED.func_state_RNI6RANZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBK1U_1_1_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__21416\,
            in1 => \N__28249\,
            in2 => \N__25596\,
            in3 => \N__24809\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m2s2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHDGK3_1_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111111"
        )
    port map (
            in0 => \N__27798\,
            in1 => \N__24780\,
            in2 => \N__21410\,
            in3 => \N__23954\,
            lcout => \POWERLED.N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_rep1_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22029\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26033\,
            lcout => \SUSWARN_N_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI4VID3_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__21407\,
            in1 => \N__24746\,
            in2 => \N__21818\,
            in3 => \N__28160\,
            lcout => \POWERLED.func_state_1_m0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_en_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__21833\,
            in1 => \N__23695\,
            in2 => \N__24596\,
            in3 => \N__27902\,
            lcout => \POWERLED.count_off_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_154_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22030\,
            in2 => \_gnd_net_\,
            in3 => \N__26001\,
            lcout => \G_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_11_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28156\,
            lcout => \POWERLED.count_off_RNIZ0Z_11\,
            ltout => \POWERLED.count_off_RNIZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIJ9IE1_0_0_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25579\,
            in1 => \N__27979\,
            in2 => \N__21656\,
            in3 => \N__24788\,
            lcout => \POWERLED.N_310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIBK1U_11_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24808\,
            in1 => \N__25578\,
            in2 => \_gnd_net_\,
            in3 => \N__28157\,
            lcout => OPEN,
            ltout => \POWERLED.N_314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI18EF2_11_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__27106\,
            in1 => \N__23952\,
            in2 => \N__21647\,
            in3 => \N__21629\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHDGK3_0_1_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001011"
        )
    port map (
            in0 => \N__27796\,
            in1 => \N__24777\,
            in2 => \N__21611\,
            in3 => \N__21810\,
            lcout => \POWERLED.func_state_RNIHDGK3_0Z0Z_1\,
            ltout => \POWERLED.func_state_RNIHDGK3_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIB74H7_1_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000000000"
        )
    port map (
            in0 => \N__21598\,
            in1 => \N__21587\,
            in2 => \N__21581\,
            in3 => \N__29200\,
            lcout => \POWERLED.func_state_RNIB74H7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__32402\,
            in1 => \N__28799\,
            in2 => \N__31517\,
            in3 => \N__32150\,
            lcout => \VPP_VDDQ.un9_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22171\,
            in1 => \N__25870\,
            in2 => \N__22142\,
            in3 => \N__27105\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_287_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22222\,
            in1 => \N__22136\,
            in2 => \_gnd_net_\,
            in3 => \N__22170\,
            lcout => \POWERLED.func_state_RNI_1Z0Z_0\,
            ltout => \POWERLED.func_state_RNI_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBK1U_0_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__24807\,
            in1 => \_gnd_net_\,
            in2 => \N__21821\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.func_state_RNIBK1UZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIR2IB9_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__21751\,
            in1 => \N__21728\,
            in2 => \N__23699\,
            in3 => \N__21694\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => \POWERLED.func_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1GMT1_0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__28048\,
            in1 => \N__21683\,
            in2 => \N__21674\,
            in3 => \N__27835\,
            lcout => \POWERLED.un1_clk_100khz_48_and_i_o2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_m1_0_a2_0_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22473\,
            in1 => \N__24951\,
            in2 => \_gnd_net_\,
            in3 => \N__24845\,
            lcout => \POWERLED.un1_N_3_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_52_and_i_0_0_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__24950\,
            in1 => \N__22472\,
            in2 => \N__28067\,
            in3 => \N__22386\,
            lcout => \POWERLED.un1_clk_100khz_52_and_i_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0RLE1_0_1_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__28052\,
            in1 => \N__22048\,
            in2 => \N__27880\,
            in3 => \N__27104\,
            lcout => OPEN,
            ltout => \POWERLED.N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI80TT3_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__23953\,
            in1 => \N__21671\,
            in2 => \N__21659\,
            in3 => \N__25782\,
            lcout => \POWERLED.dutycycle_set_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_0_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27733\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22245\,
            lcout => \POWERLED.func_state_RNI_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_5_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25580\,
            in2 => \_gnd_net_\,
            in3 => \N__27732\,
            lcout => \POWERLED.func_state_RNI_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_1_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__27735\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28460\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_48_and_i_o2_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIC4OR2_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__30515\,
            in1 => \N__29201\,
            in2 => \N__21923\,
            in3 => \N__21920\,
            lcout => \POWERLED.func_state_RNIC4OR2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__27734\,
            in1 => \N__22246\,
            in2 => \_gnd_net_\,
            in3 => \N__28170\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNICAC53_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21913\,
            in1 => \N__28097\,
            in2 => \N__21902\,
            in3 => \N__27659\,
            lcout => \POWERLED.func_state_RNICAC53_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21899\,
            lcout => \POWERLED.un85_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_13_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25523\,
            lcout => \POWERLED.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32935\,
            ce => \N__31218\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_14_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25508\,
            lcout => \POWERLED.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32935\,
            ce => \N__31218\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25276\,
            lcout => \POWERLED.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32935\,
            ce => \N__31218\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_3_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25391\,
            lcout => \POWERLED.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32935\,
            ce => \N__31218\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_4_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25376\,
            lcout => \POWERLED.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32935\,
            ce => \N__31218\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUI5O_12_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21950\,
            in1 => \N__32002\,
            in2 => \_gnd_net_\,
            in3 => \N__21961\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_12_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21965\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32944\,
            ce => \N__31767\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIHTPD_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21944\,
            in2 => \N__25277\,
            in3 => \N__31143\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIL756_13_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31146\,
            in1 => \N__21938\,
            in2 => \_gnd_net_\,
            in3 => \N__25522\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINA66_14_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21932\,
            in1 => \N__31147\,
            in2 => \_gnd_net_\,
            in3 => \N__25507\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPD76_15_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31148\,
            in1 => \N__25478\,
            in2 => \_gnd_net_\,
            in3 => \N__25489\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIJ0RD_3_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22262\,
            in1 => \N__31144\,
            in2 => \_gnd_net_\,
            in3 => \N__25390\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIL3SD_4_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31145\,
            in1 => \N__22256\,
            in2 => \_gnd_net_\,
            in3 => \N__25375\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_5_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26153\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_5\,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__26788\,
            in1 => \_gnd_net_\,
            in2 => \N__22250\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_10Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_1_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25597\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27767\,
            lcout => \POWERLED.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__22244\,
            in1 => \N__22183\,
            in2 => \N__22169\,
            in3 => \N__22122\,
            lcout => \POWERLED.N_390\,
            ltout => \POWERLED.N_390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI39RS_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111111"
        )
    port map (
            in0 => \N__28065\,
            in1 => \N__22076\,
            in2 => \N__22052\,
            in3 => \N__22041\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_3_0_0_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIN7N72_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__24004\,
            in1 => \N__27859\,
            in2 => \N__22001\,
            in3 => \N__26016\,
            lcout => \POWERLED.dutycycle_eena_3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.slp_s3n_signal_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22464\,
            in2 => \_gnd_net_\,
            in3 => \N__24853\,
            lcout => slp_s3n_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_m1_e_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__22465\,
            in1 => \N__24922\,
            in2 => \_gnd_net_\,
            in3 => \N__22399\,
            lcout => \POWERLED.dutycycle_N_3_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILP0F_5_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__22334\,
            in1 => \N__22328\,
            in2 => \_gnd_net_\,
            in3 => \N__30483\,
            lcout => \POWERLED.un1_clk_100khz_52_and_i_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_5_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27794\,
            in1 => \_gnd_net_\,
            in2 => \N__26193\,
            in3 => \N__27093\,
            lcout => \POWERLED.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__25447\,
            in2 => \_gnd_net_\,
            in3 => \N__28473\,
            lcout => \POWERLED.un1_dutycycle_172_sm3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI1U7M2_5_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__26053\,
            in1 => \N__22555\,
            in2 => \N__26192\,
            in3 => \N__26039\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNICFHA6_5_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111000"
        )
    port map (
            in0 => \N__27113\,
            in1 => \N__22322\,
            in2 => \N__22316\,
            in3 => \N__30482\,
            lcout => OPEN,
            ltout => \POWERLED.N_225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIG6629_5_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22313\,
            in2 => \N__22304\,
            in3 => \N__23903\,
            lcout => \POWERLED.dutycycle_eena_14\,
            ltout => \POWERLED.dutycycle_eena_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNICPVSD_5_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__22286\,
            in1 => \N__22270\,
            in2 => \N__22301\,
            in3 => \N__23703\,
            lcout => \POWERLED.dutycycleZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__22271\,
            in1 => \N__22298\,
            in2 => \N__23738\,
            in3 => \N__22285\,
            lcout => \POWERLED.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33110\,
            ce => 'H',
            sr => \N__22906\
        );

    \POWERLED.dutycycle_3_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__25767\,
            in1 => \N__22499\,
            in2 => \N__22582\,
            in3 => \N__22595\,
            lcout => \POWERLED.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33123\,
            ce => 'H',
            sr => \N__22904\
        );

    \POWERLED.dutycycle_RNI59UL8_3_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__22498\,
            in1 => \N__22594\,
            in2 => \N__22583\,
            in3 => \N__25766\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => \POWERLED.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__26394\,
            in1 => \_gnd_net_\,
            in2 => \N__22562\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_3\,
            ltout => \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111111"
        )
    port map (
            in0 => \N__25891\,
            in1 => \N__26948\,
            in2 => \N__22559\,
            in3 => \N__26711\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_3_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26395\,
            in1 => \N__26681\,
            in2 => \_gnd_net_\,
            in3 => \N__23134\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_7_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__22520\,
            in1 => \_gnd_net_\,
            in2 => \N__23138\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_7_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111010"
        )
    port map (
            in0 => \N__26575\,
            in1 => \N__22519\,
            in2 => \N__24425\,
            in3 => \N__23133\,
            lcout => \POWERLED.un1_dutycycle_53_13_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111111"
        )
    port map (
            in0 => \N__26390\,
            in1 => \N__24416\,
            in2 => \N__26693\,
            in3 => \N__26574\,
            lcout => \POWERLED.un1_dutycycle_53_31_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4VJH7_3_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__24083\,
            in1 => \N__22687\,
            in2 => \N__26692\,
            in3 => \N__22708\,
            lcout => \POWERLED.dutycycle_en_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4VJH7_4_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__22688\,
            in1 => \N__24081\,
            in2 => \N__26401\,
            in3 => \N__22704\,
            lcout => \POWERLED.dutycycle_RNI4VJH7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4VJH7_8_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__24082\,
            in1 => \N__24414\,
            in2 => \N__22709\,
            in3 => \N__22686\,
            lcout => \POWERLED.dutycycle_en_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_7_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__24413\,
            in1 => \N__26357\,
            in2 => \_gnd_net_\,
            in3 => \N__23120\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_10_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_9_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__22741\,
            in1 => \N__23260\,
            in2 => \N__22652\,
            in3 => \N__24281\,
            lcout => \POWERLED.un1_dutycycle_53_10_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_7_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26613\,
            in2 => \_gnd_net_\,
            in3 => \N__23119\,
            lcout => \POWERLED.un1_dutycycle_53_31_a7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_9_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26770\,
            lcout => \POWERLED.N_2200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_12_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__26852\,
            in1 => \N__24415\,
            in2 => \_gnd_net_\,
            in3 => \N__24167\,
            lcout => \POWERLED.un2_count_clk_17_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI7CVL8_4_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__22631\,
            in1 => \N__25815\,
            in2 => \N__22619\,
            in3 => \N__22603\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__25813\,
            in1 => \N__22630\,
            in2 => \N__22607\,
            in3 => \N__22618\,
            lcout => \POWERLED.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33128\,
            ce => 'H',
            sr => \N__22901\
        );

    \POWERLED.dutycycle_RNIDP3K7_11_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22915\,
            in1 => \N__22720\,
            in2 => \N__25823\,
            in3 => \N__22924\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => \POWERLED.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_11_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23048\,
            in3 => \N__23244\,
            lcout => \POWERLED.un1_dutycycle_53_50_a0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_12_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__24168\,
            in1 => \N__24283\,
            in2 => \N__23465\,
            in3 => \N__23034\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__22970\,
            in1 => \N__22949\,
            in2 => \N__22943\,
            in3 => \N__24422\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__22916\,
            in1 => \N__25814\,
            in2 => \N__22727\,
            in3 => \N__22925\,
            lcout => \POWERLED.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33128\,
            ce => 'H',
            sr => \N__22901\
        );

    \POWERLED.dutycycle_RNI_11_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001010"
        )
    port map (
            in0 => \N__24282\,
            in1 => \N__23442\,
            in2 => \N__22745\,
            in3 => \N__23245\,
            lcout => \POWERLED.un1_dutycycle_53_50_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN3GO3_11_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__28446\,
            in1 => \N__25810\,
            in2 => \N__24100\,
            in3 => \N__23433\,
            lcout => OPEN,
            ltout => \POWERLED.N_144_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEB706_11_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011000100"
        )
    port map (
            in0 => \N__23944\,
            in1 => \N__23813\,
            in2 => \N__22730\,
            in3 => \N__24011\,
            lcout => \POWERLED.dutycycle_en_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIBVNS_4_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28448\,
            in2 => \_gnd_net_\,
            in3 => \N__25811\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNIBVNSZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOMK66_9_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111111"
        )
    port map (
            in0 => \N__24087\,
            in1 => \N__23174\,
            in2 => \N__23528\,
            in3 => \N__23951\,
            lcout => \POWERLED.dutycycle_eena_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFS4K7_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23513\,
            in1 => \N__25812\,
            in2 => \N__23488\,
            in3 => \N__23635\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => \POWERLED.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_12_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__23434\,
            in1 => \_gnd_net_\,
            in2 => \N__23393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_51_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_15_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__23390\,
            in1 => \N__23384\,
            in2 => \N__23333\,
            in3 => \N__23330\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBVNS_9_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111110"
        )
    port map (
            in0 => \N__28447\,
            in1 => \N__24012\,
            in2 => \N__23306\,
            in3 => \N__23231\,
            lcout => \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_7_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__23104\,
            in1 => \N__26622\,
            in2 => \N__24420\,
            in3 => \N__26380\,
            lcout => \POWERLED.dutycycle_RNI_8Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__26381\,
            in1 => \N__23106\,
            in2 => \N__26627\,
            in3 => \N__24398\,
            lcout => \POWERLED.N_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_3_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__23107\,
            in1 => \N__26694\,
            in2 => \N__24421\,
            in3 => \N__26383\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_7_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__26382\,
            in1 => \N__23105\,
            in2 => \_gnd_net_\,
            in3 => \N__26626\,
            lcout => OPEN,
            ltout => \POWERLED.g0_i_a6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_12_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__24402\,
            in1 => \N__24284\,
            in2 => \N__24188\,
            in3 => \N__24156\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIN3GO3_12_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__25809\,
            in1 => \N__24157\,
            in2 => \N__28474\,
            in3 => \N__24080\,
            lcout => OPEN,
            ltout => \POWERLED.N_145_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEB706_12_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__24013\,
            in1 => \N__23950\,
            in2 => \N__23816\,
            in3 => \N__23737\,
            lcout => \POWERLED.dutycycle_en_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_0_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23620\,
            in2 => \N__23609\,
            in3 => \N__23608\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23588\,
            in2 => \_gnd_net_\,
            in3 => \N__23576\,
            lcout => \HDA_STRAP.countZ0Z_1\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_0\,
            carryout => \HDA_STRAP.un1_count_1_cry_1\,
            clk => \N__32747\,
            ce => \N__29395\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23569\,
            in2 => \_gnd_net_\,
            in3 => \N__23558\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_1\,
            carryout => \HDA_STRAP.un1_count_1_cry_2\,
            clk => \N__32747\,
            ce => \N__29395\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23555\,
            in2 => \_gnd_net_\,
            in3 => \N__23543\,
            lcout => \HDA_STRAP.countZ0Z_3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_2\,
            carryout => \HDA_STRAP.un1_count_1_cry_3\,
            clk => \N__32747\,
            ce => \N__29395\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23540\,
            in2 => \_gnd_net_\,
            in3 => \N__24587\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_3\,
            carryout => \HDA_STRAP.un1_count_1_cry_4\,
            clk => \N__32747\,
            ce => \N__29395\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24584\,
            in2 => \_gnd_net_\,
            in3 => \N__24572\,
            lcout => \HDA_STRAP.countZ0Z_5\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_4\,
            carryout => \HDA_STRAP.un1_count_1_cry_5\,
            clk => \N__32747\,
            ce => \N__29395\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_6_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24569\,
            in2 => \_gnd_net_\,
            in3 => \N__24548\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_5\,
            carryout => \HDA_STRAP.un1_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24538\,
            in2 => \_gnd_net_\,
            in3 => \N__24527\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_6\,
            carryout => \HDA_STRAP.un1_count_1_cry_7\,
            clk => \N__32747\,
            ce => \N__29395\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_8_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24520\,
            in2 => \_gnd_net_\,
            in3 => \N__24503\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24500\,
            in2 => \_gnd_net_\,
            in3 => \N__24488\,
            lcout => \HDA_STRAP.countZ0Z_9\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_8\,
            carryout => \HDA_STRAP.un1_count_1_cry_9\,
            clk => \N__32911\,
            ce => \N__29401\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_10_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24485\,
            in2 => \_gnd_net_\,
            in3 => \N__24464\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_9\,
            carryout => \HDA_STRAP.un1_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_11_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24461\,
            in2 => \_gnd_net_\,
            in3 => \N__24443\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_10\,
            carryout => \HDA_STRAP.un1_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24440\,
            in2 => \_gnd_net_\,
            in3 => \N__24428\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_11\,
            carryout => \HDA_STRAP.un1_count_1_cry_12\,
            clk => \N__32911\,
            ce => \N__29401\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24710\,
            in2 => \_gnd_net_\,
            in3 => \N__24698\,
            lcout => \HDA_STRAP.countZ0Z_13\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_12\,
            carryout => \HDA_STRAP.un1_count_1_cry_13\,
            clk => \N__32911\,
            ce => \N__29401\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24695\,
            in2 => \_gnd_net_\,
            in3 => \N__24683\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_13\,
            carryout => \HDA_STRAP.un1_count_1_cry_14\,
            clk => \N__32911\,
            ce => \N__29401\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24680\,
            in2 => \_gnd_net_\,
            in3 => \N__24668\,
            lcout => \HDA_STRAP.countZ0Z_15\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_14\,
            carryout => \HDA_STRAP.un1_count_1_cry_15\,
            clk => \N__32911\,
            ce => \N__29401\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_16_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24665\,
            in2 => \_gnd_net_\,
            in3 => \N__24647\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_17_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24644\,
            in2 => \_gnd_net_\,
            in3 => \N__24626\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__27107\,
            in1 => \N__28030\,
            in2 => \N__27884\,
            in3 => \N__28159\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_o_N_305_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111100"
        )
    port map (
            in0 => \N__28029\,
            in1 => \N__24611\,
            in2 => \N__24602\,
            in3 => \N__30547\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__28200\,
            in1 => \N__28640\,
            in2 => \N__24599\,
            in3 => \N__27800\,
            lcout => \POWERLED.un1_func_state25_6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_ss0_i_0_x2_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29238\,
            in3 => \N__30546\,
            lcout => \POWERLED.N_150_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJ9IE1_11_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__24781\,
            in1 => \N__28028\,
            in2 => \_gnd_net_\,
            in3 => \N__28158\,
            lcout => \POWERLED.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIR1479_9_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24724\,
            in1 => \N__24733\,
            in2 => \_gnd_net_\,
            in3 => \N__30715\,
            lcout => \POWERLED.un3_count_off_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30925\,
            in2 => \_gnd_net_\,
            in3 => \N__29944\,
            lcout => \POWERLED.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32942\,
            ce => \N__30751\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__29980\,
            in1 => \_gnd_net_\,
            in2 => \N__30932\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32942\,
            ce => \N__30751\,
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNISUHQ2_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30923\,
            in2 => \_gnd_net_\,
            in3 => \N__29981\,
            lcout => \POWERLED.count_off_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI4C959_10_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__30924\,
            in1 => \N__24740\,
            in2 => \N__29948\,
            in3 => \N__30714\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => \POWERLED.count_offZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIR1479_0_9_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__24734\,
            in1 => \N__24725\,
            in2 => \N__24716\,
            in3 => \N__30753\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIG5N6N1_11_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25259\,
            in1 => \N__27548\,
            in2 => \N__24713\,
            in3 => \N__29831\,
            lcout => \POWERLED.count_off_RNIG5N6N1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDJM39_0_11_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000101"
        )
    port map (
            in0 => \N__29909\,
            in1 => \N__27599\,
            in2 => \N__27584\,
            in3 => \N__30752\,
            lcout => \POWERLED.un34_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25253\,
            in2 => \N__25223\,
            in3 => \N__25190\,
            lcout => \POWERLED.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32971\,
            ce => \N__31766\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIHTOU_8_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32401\,
            in1 => \N__32234\,
            in2 => \_gnd_net_\,
            in3 => \N__32207\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIM9AN_1_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28795\,
            in1 => \N__32400\,
            in2 => \_gnd_net_\,
            in3 => \N__31510\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_1\,
            ltout => \VPP_VDDQ.un1_count_2_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25151\,
            in3 => \N__32149\,
            lcout => \VPP_VDDQ.count_2_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25141\,
            in2 => \N__25099\,
            in3 => \N__25044\,
            lcout => \POWERLED.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32971\,
            ce => \N__31766\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25091\,
            in2 => \_gnd_net_\,
            in3 => \N__25045\,
            lcout => \POWERLED.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32971\,
            ce => \N__31766\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.VCCST_EN_0_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24844\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIN6TD_5_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31202\,
            in1 => \N__25301\,
            in2 => \_gnd_net_\,
            in3 => \N__25360\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_5_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33099\,
            ce => \N__31223\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIP9UD_6_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31203\,
            in1 => \N__25295\,
            in2 => \_gnd_net_\,
            in3 => \N__25348\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_6_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33099\,
            ce => \N__31223\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNITF0E_8_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31204\,
            in1 => \N__25289\,
            in2 => \_gnd_net_\,
            in3 => \N__25333\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_8_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33099\,
            ce => \N__31223\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIVI1E_9_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31205\,
            in1 => \N__25283\,
            in2 => \_gnd_net_\,
            in3 => \N__25321\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_9_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33099\,
            ce => \N__31223\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31352\,
            in2 => \N__31085\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31315\,
            in1 => \_gnd_net_\,
            in2 => \N__28609\,
            in3 => \N__25262\,
            lcout => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_1\,
            carryout => \POWERLED.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31251\,
            in1 => \_gnd_net_\,
            in2 => \N__28585\,
            in3 => \N__25379\,
            lcout => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_2\,
            carryout => \POWERLED.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31316\,
            in1 => \_gnd_net_\,
            in2 => \N__28503\,
            in3 => \N__25364\,
            lcout => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_3\,
            carryout => \POWERLED.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31252\,
            in1 => \_gnd_net_\,
            in2 => \N__31032\,
            in3 => \N__25352\,
            lcout => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_4\,
            carryout => \POWERLED.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31317\,
            in1 => \_gnd_net_\,
            in2 => \N__28560\,
            in3 => \N__25340\,
            lcout => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_5\,
            carryout => \POWERLED.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31253\,
            in1 => \_gnd_net_\,
            in2 => \N__28313\,
            in3 => \N__25337\,
            lcout => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_6\,
            carryout => \POWERLED.un1_count_clk_2_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31318\,
            in1 => \_gnd_net_\,
            in2 => \N__28528\,
            in3 => \N__25325\,
            lcout => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_7_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31319\,
            in1 => \_gnd_net_\,
            in2 => \N__31002\,
            in3 => \N__25310\,
            lcout => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28724\,
            in3 => \N__25307\,
            lcout => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_9_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31424\,
            in2 => \_gnd_net_\,
            in3 => \N__25304\,
            lcout => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_10_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31366\,
            in2 => \_gnd_net_\,
            in3 => \N__25526\,
            lcout => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_11\,
            carryout => \POWERLED.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31320\,
            in1 => \_gnd_net_\,
            in2 => \N__28693\,
            in3 => \N__25511\,
            lcout => \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_12\,
            carryout => \POWERLED.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__31321\,
            in1 => \_gnd_net_\,
            in2 => \N__28672\,
            in3 => \N__25496\,
            lcout => \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_13\,
            carryout => \POWERLED.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__28708\,
            in1 => \N__31322\,
            in2 => \_gnd_net_\,
            in3 => \N__25493\,
            lcout => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_15_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25490\,
            lcout => \POWERLED.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32943\,
            ce => \N__31217\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31206\,
            in1 => \N__25460\,
            in2 => \_gnd_net_\,
            in3 => \N__25471\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_7_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25472\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32972\,
            ce => \N__31207\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__25454\,
            in1 => \N__26831\,
            in2 => \_gnd_net_\,
            in3 => \N__28424\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25436\,
            in3 => \N__25412\,
            lcout => \POWERLED.mult1_un47_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__26097\,
            in1 => \N__26098\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBVNS_5_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__26170\,
            in1 => \N__25889\,
            in2 => \N__26063\,
            in3 => \N__26832\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m4_bm_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMUFP1_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25846\,
            in2 => \N__26042\,
            in3 => \N__25907\,
            lcout => \POWERLED.dutycycle_RNIMUFP1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_9_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32008\,
            in2 => \_gnd_net_\,
            in3 => \N__26031\,
            lcout => \G_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_2_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__25890\,
            in1 => \N__26171\,
            in2 => \N__26288\,
            in3 => \N__26707\,
            lcout => \POWERLED.un1_dutycycle_172_m4_bm_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_4_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28428\,
            in2 => \_gnd_net_\,
            in3 => \N__27077\,
            lcout => \POWERLED.N_20_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBVNS_2_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25818\,
            in1 => \N__25603\,
            in2 => \_gnd_net_\,
            in3 => \N__26282\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMUFP1_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000011101"
        )
    port map (
            in0 => \N__25847\,
            in1 => \N__26840\,
            in2 => \N__25826\,
            in3 => \N__26833\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m3_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1U7M2_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__25819\,
            in1 => \N__25604\,
            in2 => \N__25529\,
            in3 => \N__27119\,
            lcout => \POWERLED.un1_dutycycle_172_m3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__26487\,
            in1 => \N__26939\,
            in2 => \N__27098\,
            in3 => \N__28429\,
            lcout => \POWERLED.un1_dutycycle_96_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__26940\,
            in1 => \N__26851\,
            in2 => \N__28461\,
            in3 => \N__26488\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__26675\,
            in1 => \N__26273\,
            in2 => \_gnd_net_\,
            in3 => \N__26607\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101001011"
        )
    port map (
            in0 => \N__26834\,
            in1 => \N__26483\,
            in2 => \N__26810\,
            in3 => \N__26396\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_2_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26807\,
            in3 => \N__26274\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__26795\,
            in1 => \N__26777\,
            in2 => \N__28462\,
            in3 => \N__26749\,
            lcout => \POWERLED.dutycycle_RNI_9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_3_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__26676\,
            in1 => \N__26393\,
            in2 => \N__26492\,
            in3 => \N__26606\,
            lcout => \POWERLED.un1_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__26489\,
            in1 => \N__26397\,
            in2 => \N__26286\,
            in3 => \N__26166\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27272\,
            in1 => \N__27254\,
            in2 => \N__27215\,
            in3 => \N__27160\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27488\,
            in1 => \N__27506\,
            in2 => \N__27377\,
            in3 => \N__27524\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27173\,
            in1 => \N__27182\,
            in2 => \N__27176\,
            in3 => \N__27167\,
            lcout => \VPP_VDDQ.un6_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27319\,
            in1 => \N__27334\,
            in2 => \N__27290\,
            in3 => \N__27349\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27304\,
            in1 => \N__27148\,
            in2 => \N__27236\,
            in3 => \N__27133\,
            lcout => \VPP_VDDQ.un6_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29588\,
            in1 => \N__27161\,
            in2 => \N__29162\,
            in3 => \N__29161\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29584\,
            in1 => \N__27149\,
            in2 => \_gnd_net_\,
            in3 => \N__27137\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29589\,
            in1 => \N__27134\,
            in2 => \_gnd_net_\,
            in3 => \N__27122\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29585\,
            in1 => \N__27350\,
            in2 => \_gnd_net_\,
            in3 => \N__27338\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29590\,
            in1 => \N__27335\,
            in2 => \_gnd_net_\,
            in3 => \N__27323\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29586\,
            in1 => \N__27320\,
            in2 => \_gnd_net_\,
            in3 => \N__27308\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_6_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29591\,
            in1 => \N__27305\,
            in2 => \_gnd_net_\,
            in3 => \N__27293\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29587\,
            in1 => \N__27289\,
            in2 => \_gnd_net_\,
            in3 => \N__27275\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__33142\,
            ce => 'H',
            sr => \N__29129\
        );

    \VPP_VDDQ.count_8_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29583\,
            in1 => \N__27271\,
            in2 => \_gnd_net_\,
            in3 => \N__27257\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__33138\,
            ce => 'H',
            sr => \N__29128\
        );

    \VPP_VDDQ.count_9_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29579\,
            in1 => \N__27253\,
            in2 => \_gnd_net_\,
            in3 => \N__27239\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__33138\,
            ce => 'H',
            sr => \N__29128\
        );

    \VPP_VDDQ.count_10_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29580\,
            in1 => \N__27232\,
            in2 => \_gnd_net_\,
            in3 => \N__27218\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__33138\,
            ce => 'H',
            sr => \N__29128\
        );

    \VPP_VDDQ.count_11_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29577\,
            in1 => \N__27211\,
            in2 => \_gnd_net_\,
            in3 => \N__27197\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__33138\,
            ce => 'H',
            sr => \N__29128\
        );

    \VPP_VDDQ.count_12_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29581\,
            in1 => \N__27523\,
            in2 => \_gnd_net_\,
            in3 => \N__27509\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__33138\,
            ce => 'H',
            sr => \N__29128\
        );

    \VPP_VDDQ.count_13_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29578\,
            in1 => \N__27505\,
            in2 => \_gnd_net_\,
            in3 => \N__27491\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__33138\,
            ce => 'H',
            sr => \N__29128\
        );

    \VPP_VDDQ.count_14_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29582\,
            in1 => \N__27487\,
            in2 => \_gnd_net_\,
            in3 => \N__27473\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__33138\,
            ce => 'H',
            sr => \N__29128\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27449\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27373\,
            in2 => \_gnd_net_\,
            in3 => \N__27380\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33140\,
            ce => \N__29093\,
            sr => \N__29121\
        );

    \POWERLED.count_off_RNIJLV69_5_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__30921\,
            in1 => \N__29761\,
            in2 => \N__27359\,
            in3 => \N__30761\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29762\,
            in3 => \N__30922\,
            lcout => \POWERLED.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32906\,
            ce => \N__30782\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30160\,
            in2 => \_gnd_net_\,
            in3 => \N__30917\,
            lcout => \POWERLED.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32906\,
            ce => \N__30782\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30918\,
            lcout => \POWERLED.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32906\,
            ce => \N__30782\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNILVQ39_15_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__30920\,
            in1 => \N__27563\,
            in2 => \N__30784\,
            in3 => \N__30184\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30919\,
            lcout => \POWERLED.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32906\,
            ce => \N__30782\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIPU279_8_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__30916\,
            in1 => \N__27557\,
            in2 => \N__30785\,
            in3 => \N__30005\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29794\,
            in2 => \_gnd_net_\,
            in3 => \N__30931\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33029\,
            ce => \N__30765\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDCS69_0_2_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__29776\,
            in1 => \N__27641\,
            in2 => \N__30777\,
            in3 => \N__27632\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI8GSR41_2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27614\,
            in1 => \N__30116\,
            in2 => \N__27551\,
            in3 => \N__27539\,
            lcout => \POWERLED.un34_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNILO079_0_6_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__29819\,
            in1 => \N__27533\,
            in2 => \N__30778\,
            in3 => \N__28271\,
            lcout => \POWERLED.un34_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNIPOEQ2_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29741\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30929\,
            lcout => \POWERLED.count_off_1_6\,
            ltout => \POWERLED.count_off_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNILO079_6_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__30734\,
            in1 => \N__28270\,
            in2 => \N__27527\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un3_count_off_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNILGAQ2_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29795\,
            in2 => \_gnd_net_\,
            in3 => \N__30930\,
            lcout => \POWERLED.count_off_1_2\,
            ltout => \POWERLED.count_off_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDCS69_2_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30735\,
            in1 => \_gnd_net_\,
            in2 => \N__27635\,
            in3 => \N__27631\,
            lcout => \POWERLED.un3_count_off_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNINR179_7_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30766\,
            in1 => \N__27607\,
            in2 => \_gnd_net_\,
            in3 => \N__27623\,
            lcout => \POWERLED.un3_count_off_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNIQQFQ2_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30032\,
            in2 => \_gnd_net_\,
            in3 => \N__30853\,
            lcout => \POWERLED.count_off_1_7\,
            ltout => \POWERLED.count_off_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNINR179_0_7_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__30787\,
            in1 => \N__27608\,
            in2 => \N__27617\,
            in3 => \N__30020\,
            lcout => \POWERLED.un34_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30031\,
            in2 => \_gnd_net_\,
            in3 => \N__30857\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32907\,
            ce => \N__30786\,
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNI570P2_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30854\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29921\,
            lcout => \POWERLED.count_off_1_11\,
            ltout => \POWERLED.count_off_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDJM39_11_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27574\,
            in2 => \N__27587\,
            in3 => \N__30767\,
            lcout => \POWERLED.un3_count_off_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30855\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29920\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32907\,
            ce => \N__30786\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29740\,
            in2 => \_gnd_net_\,
            in3 => \N__30856\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32907\,
            ce => \N__30786\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIJ9IE1_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28282\,
            in1 => \N__28262\,
            in2 => \_gnd_net_\,
            in3 => \N__28087\,
            lcout => OPEN,
            ltout => \POWERLED.N_289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIU8AB2_7_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__28632\,
            in1 => \N__28241\,
            in2 => \N__28211\,
            in3 => \N__28208\,
            lcout => \POWERLED.N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_8_1_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__28178\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28120\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_2_tz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIRKB61_1_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__28283\,
            in1 => \N__28001\,
            in2 => \N__28100\,
            in3 => \N__27883\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27882\,
            in1 => \N__28088\,
            in2 => \N__28041\,
            in3 => \N__28281\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_304_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100011"
        )
    port map (
            in0 => \N__28633\,
            in1 => \N__27881\,
            in2 => \N__27799\,
            in3 => \N__28340\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_4_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28561\,
            in2 => \_gnd_net_\,
            in3 => \N__28510\,
            lcout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_2_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__28615\,
            in1 => \N__28534\,
            in2 => \N__27650\,
            in3 => \N__28591\,
            lcout => \POWERLED.N_352\,
            ltout => \POWERLED.N_352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_7_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28315\,
            in2 => \N__28643\,
            in3 => \N__30968\,
            lcout => \POWERLED.N_394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__31607\,
            in1 => \N__33660\,
            in2 => \_gnd_net_\,
            in3 => \N__32001\,
            lcout => \VPP_VDDQ.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33431\,
            lcout => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__28616\,
            in1 => \N__28592\,
            in2 => \N__28568\,
            in3 => \N__28535\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_4_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__28511\,
            in1 => \N__28316\,
            in2 => \N__28478\,
            in3 => \N__30967\,
            lcout => \POWERLED.N_2182_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__31039\,
            in1 => \N__31076\,
            in2 => \_gnd_net_\,
            in3 => \N__31051\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_9_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__28322\,
            in1 => \N__28314\,
            in2 => \N__28286\,
            in3 => \N__31003\,
            lcout => \POWERLED.count_clk_RNIZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_10_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__28736\,
            in1 => \_gnd_net_\,
            in2 => \N__31314\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33048\,
            ce => \N__31201\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8SH6_10_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__31162\,
            in1 => \N__31285\,
            in2 => \N__28745\,
            in3 => \N__28735\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => \POWERLED.count_clkZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_15_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31367\,
            in1 => \N__31423\,
            in2 => \N__28712\,
            in3 => \N__28709\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_13_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31345\,
            in1 => \N__28694\,
            in2 => \N__28676\,
            in3 => \N__28673\,
            lcout => \POWERLED.N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31286\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31346\,
            lcout => \POWERLED.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33048\,
            ce => \N__31201\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31347\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31283\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIQF8B_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28655\,
            in2 => \N__28649\,
            in3 => \N__31161\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => \POWERLED.count_clkZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__31078\,
            in1 => \_gnd_net_\,
            in2 => \N__28646\,
            in3 => \N__31284\,
            lcout => \POWERLED.count_clk_RNIZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33397\,
            in1 => \N__33557\,
            in2 => \N__33297\,
            in3 => \N__28822\,
            lcout => \VPP_VDDQ.count_2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33558\,
            in1 => \N__33277\,
            in2 => \N__28826\,
            in3 => \N__33402\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33100\,
            ce => \N__32429\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__28948\,
            in1 => \N__33567\,
            in2 => \N__33451\,
            in3 => \N__33282\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJ0QU_9_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28805\,
            in1 => \_gnd_net_\,
            in2 => \N__28808\,
            in3 => \N__32363\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33399\,
            in1 => \N__33560\,
            in2 => \N__28949\,
            in3 => \N__33281\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33100\,
            ce => \N__32429\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33278\,
            in1 => \N__31541\,
            in2 => \N__33620\,
            in3 => \N__33401\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33100\,
            ce => \N__32429\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33398\,
            in1 => \N__33559\,
            in2 => \N__31484\,
            in3 => \N__33280\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33100\,
            ce => \N__32429\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33279\,
            in1 => \N__33400\,
            in2 => \N__33621\,
            in3 => \N__29006\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33100\,
            ce => \N__32429\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI5BIU_0_2_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__32359\,
            in1 => \N__31460\,
            in2 => \N__28874\,
            in3 => \N__31447\,
            lcout => \VPP_VDDQ.un9_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIBKLU_0_5_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__28981\,
            in1 => \N__32361\,
            in2 => \N__28889\,
            in3 => \N__28898\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFQ6J3_1_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28775\,
            in1 => \N__28760\,
            in2 => \N__28754\,
            in3 => \N__28751\,
            lcout => \VPP_VDDQ.un9_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI9HKU_0_4_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000111"
        )
    port map (
            in0 => \N__28907\,
            in1 => \N__32360\,
            in2 => \N__31703\,
            in3 => \N__28918\,
            lcout => \VPP_VDDQ.un9_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI9HKU_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32357\,
            in1 => \_gnd_net_\,
            in2 => \N__28919\,
            in3 => \N__28906\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33428\,
            in1 => \N__33268\,
            in2 => \N__33657\,
            in3 => \N__29002\,
            lcout => \VPP_VDDQ.count_2_1_5\,
            ltout => \VPP_VDDQ.count_2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIBKLU_5_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32358\,
            in1 => \_gnd_net_\,
            in2 => \N__28892\,
            in3 => \N__28885\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI5BIU_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31459\,
            in1 => \N__28870\,
            in2 => \_gnd_net_\,
            in3 => \N__32356\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32135\,
            in2 => \N__28862\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28844\,
            in2 => \_gnd_net_\,
            in3 => \N__28838\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31448\,
            in2 => \_gnd_net_\,
            in3 => \N__28835\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28832\,
            in2 => \_gnd_net_\,
            in3 => \N__28811\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29012\,
            in2 => \_gnd_net_\,
            in3 => \N__28991\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31696\,
            in2 => \_gnd_net_\,
            in3 => \N__28988\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32075\,
            in2 => \_gnd_net_\,
            in3 => \N__28985\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28982\,
            in2 => \_gnd_net_\,
            in3 => \N__28952\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31574\,
            in2 => \_gnd_net_\,
            in3 => \N__28934\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33671\,
            in2 => \_gnd_net_\,
            in3 => \N__28931\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32192\,
            in2 => \_gnd_net_\,
            in3 => \N__28928\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32065\,
            in2 => \_gnd_net_\,
            in3 => \N__28925\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29054\,
            in3 => \N__28922\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32029\,
            in2 => \_gnd_net_\,
            in3 => \N__29078\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29038\,
            in2 => \_gnd_net_\,
            in3 => \N__29075\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_15_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32030\,
            in1 => \N__32066\,
            in2 => \N__29039\,
            in3 => \N__29053\,
            lcout => \VPP_VDDQ.un9_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33290\,
            in1 => \N__33465\,
            in2 => \N__33664\,
            in3 => \N__29071\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33136\,
            ce => \N__32418\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__29072\,
            in1 => \N__33654\,
            in2 => \N__33473\,
            in3 => \N__33293\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI98N41_13_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32381\,
            in1 => \_gnd_net_\,
            in2 => \N__29063\,
            in3 => \N__29060\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33655\,
            in1 => \N__33470\,
            in2 => \N__33299\,
            in3 => \N__29026\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIDEP41_15_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29018\,
            in2 => \N__29042\,
            in3 => \N__32382\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__33466\,
            in2 => \N__33665\,
            in3 => \N__29027\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33136\,
            ce => \N__32418\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33464\,
            in1 => \N__33647\,
            in2 => \N__32056\,
            in3 => \N__33292\,
            lcout => \VPP_VDDQ.count_2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33136\,
            ce => \N__32418\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__29268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29138\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29267\,
            lcout => \VPP_VDDQ.N_360\,
            ltout => \VPP_VDDQ.N_360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29620\,
            in2 => \N__29165\,
            in3 => \N__29681\,
            lcout => \VPP_VDDQ.N_264_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110010101010"
        )
    port map (
            in0 => \N__29137\,
            in1 => \N__29726\,
            in2 => \N__29624\,
            in3 => \N__29575\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__29576\,
            in1 => \N__29084\,
            in2 => \N__29141\,
            in3 => \N__29646\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNITROD7_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__29725\,
            in1 => \N__29617\,
            in2 => \N__29714\,
            in3 => \N__29547\,
            lcout => \VPP_VDDQ.curr_state_RNITROD7Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_RNITROD7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29548\,
            in1 => \_gnd_net_\,
            in2 => \N__29096\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.N_27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__29675\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29618\,
            lcout => \VPP_VDDQ.N_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29673\,
            in2 => \_gnd_net_\,
            in3 => \N__29640\,
            lcout => \VPP_VDDQ.N_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI8I855_0_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29674\,
            in1 => \N__29616\,
            in2 => \_gnd_net_\,
            in3 => \N__29704\,
            lcout => \VPP_VDDQ.N_214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010101110"
        )
    port map (
            in0 => \N__29680\,
            in1 => \N__29619\,
            in2 => \N__29651\,
            in3 => \N__29705\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33112\,
            ce => \N__29416\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29679\,
            in2 => \_gnd_net_\,
            in3 => \N__29650\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33112\,
            ce => \N__29416\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIFMN39_12_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29306\,
            in1 => \N__30911\,
            in2 => \N__29888\,
            in3 => \N__30775\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_1_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29817\,
            in2 => \_gnd_net_\,
            in3 => \N__30066\,
            lcout => \POWERLED.count_off_RNIZ0Z_1\,
            ltout => \POWERLED.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIL3SN8_1_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29294\,
            in1 => \N__30912\,
            in2 => \N__29309\,
            in3 => \N__30776\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30913\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29884\,
            lcout => \POWERLED.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33068\,
            ce => \N__30783\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29300\,
            in2 => \_gnd_net_\,
            in3 => \N__30915\,
            lcout => \POWERLED.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33068\,
            ce => \N__30783\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30914\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29857\,
            lcout => \POWERLED.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33068\,
            ce => \N__30783\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHPO39_13_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29840\,
            in1 => \N__30910\,
            in2 => \N__29861\,
            in3 => \N__30774\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => \POWERLED.count_offZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_15_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30143\,
            in1 => \N__30065\,
            in2 => \N__29834\,
            in3 => \N__30199\,
            lcout => \POWERLED.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29818\,
            in2 => \N__30068\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNIN70F_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29801\,
            in2 => \_gnd_net_\,
            in3 => \N__29786\,
            lcout => \POWERLED.un3_count_off_1_cry_1_c_RNIN70FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_1\,
            carryout => \POWERLED.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30077\,
            in2 => \_gnd_net_\,
            in3 => \N__29783\,
            lcout => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_2\,
            carryout => \POWERLED.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30128\,
            in2 => \_gnd_net_\,
            in3 => \N__29780\,
            lcout => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_3\,
            carryout => \POWERLED.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_4_c_RNIQD3F_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29777\,
            in3 => \N__29750\,
            lcout => \POWERLED.un3_count_off_1_cry_4_c_RNIQD3FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_4\,
            carryout => \POWERLED.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNIRF4F_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29747\,
            in2 => \_gnd_net_\,
            in3 => \N__29729\,
            lcout => \POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_5\,
            carryout => \POWERLED.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNISH5F_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30038\,
            in2 => \_gnd_net_\,
            in3 => \N__30023\,
            lcout => \POWERLED.un3_count_off_1_cry_6_c_RNISH5FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_6\,
            carryout => \POWERLED.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_7_c_RNITJ6F_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30016\,
            in2 => \_gnd_net_\,
            in3 => \N__29996\,
            lcout => \POWERLED.un3_count_off_1_cry_7_c_RNITJ6FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_7\,
            carryout => \POWERLED.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNIUL7F_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29993\,
            in2 => \_gnd_net_\,
            in3 => \N__29966\,
            lcout => \POWERLED.un3_count_off_1_cry_8_c_RNIUL7FZ0\,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_9_c_RNIVN8F_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29963\,
            in2 => \_gnd_net_\,
            in3 => \N__29930\,
            lcout => \POWERLED.un3_count_off_1_cry_9_c_RNIVN8FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_9\,
            carryout => \POWERLED.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNI7ULD_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29927\,
            in2 => \_gnd_net_\,
            in3 => \N__29912\,
            lcout => \POWERLED.un3_count_off_1_cry_10_c_RNI7ULDZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_10\,
            carryout => \POWERLED.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_11_c_RNI80ND_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29905\,
            in2 => \_gnd_net_\,
            in3 => \N__29873\,
            lcout => \POWERLED.un3_count_off_1_cry_11_c_RNI80NDZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_11\,
            carryout => \POWERLED.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_12_c_RNI92OD_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29870\,
            in2 => \_gnd_net_\,
            in3 => \N__29846\,
            lcout => \POWERLED.un3_count_off_1_cry_12_c_RNI92ODZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_12\,
            carryout => \POWERLED.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_13_c_RNIA4PD_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30139\,
            in2 => \_gnd_net_\,
            in3 => \N__29843\,
            lcout => \POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_13\,
            carryout => \POWERLED.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_14_c_RNIB6QD_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30203\,
            in2 => \_gnd_net_\,
            in3 => \N__30188\,
            lcout => \POWERLED.un3_count_off_1_cry_14_c_RNIB6QDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJSP39_14_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__30173\,
            in1 => \N__30888\,
            in2 => \N__30161\,
            in3 => \N__30773\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30106\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33028\,
            ce => \N__30788\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHIU69_4_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__30794\,
            in1 => \N__30859\,
            in2 => \N__30950\,
            in3 => \N__30756\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => \POWERLED.count_offZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIFFT69_0_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__30757\,
            in1 => \N__30095\,
            in2 => \N__30119\,
            in3 => \N__30086\,
            lcout => \POWERLED.un34_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNIMIBQ2_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30107\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30858\,
            lcout => \POWERLED.count_off_1_3\,
            ltout => \POWERLED.count_off_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIFFT69_3_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30755\,
            in1 => \_gnd_net_\,
            in2 => \N__30089\,
            in3 => \N__30085\,
            lcout => \POWERLED.un3_count_off_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIK2SN8_0_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__30956\,
            in1 => \N__30860\,
            in2 => \N__30067\,
            in3 => \N__30754\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => \POWERLED.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__30861\,
            in1 => \_gnd_net_\,
            in2 => \N__30959\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33028\,
            ce => \N__30788\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30946\,
            in2 => \_gnd_net_\,
            in3 => \N__30863\,
            lcout => \POWERLED.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33028\,
            ce => \N__30788\,
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_3_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30611\,
            in1 => \N__30599\,
            in2 => \N__30587\,
            in3 => \N__30428\,
            lcout => OPEN,
            ltout => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30398\,
            in2 => \N__30392\,
            in3 => \N__30389\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__30254\,
            in1 => \N__31659\,
            in2 => \N__30245\,
            in3 => \N__30230\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_okZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNI9SRO4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30338\,
            in3 => \N__30328\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNINI731_0_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__30227\,
            in1 => \N__33661\,
            in2 => \N__31661\,
            in3 => \N__31801\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_en\,
            ltout => \VPP_VDDQ.delayed_vddq_ok_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__30241\,
            in1 => \N__31658\,
            in2 => \N__30248\,
            in3 => \N__30229\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33049\,
            ce => 'H',
            sr => \N__30215\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30228\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.N_53_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIH136_11_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__31394\,
            in1 => \N__31160\,
            in2 => \N__31409\,
            in3 => \N__31309\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_11_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31405\,
            lcout => \POWERLED.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33051\,
            ce => \N__31219\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_12_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31378\,
            in2 => \_gnd_net_\,
            in3 => \N__31313\,
            lcout => \POWERLED.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33051\,
            ce => \N__31219\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIJ446_12_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__31310\,
            in1 => \N__31388\,
            in2 => \N__31382\,
            in3 => \N__31192\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__31348\,
            in1 => \N__31312\,
            in2 => \_gnd_net_\,
            in3 => \N__31077\,
            lcout => \POWERLED.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33051\,
            ce => \N__31219\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIRG8B_1_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31229\,
            in2 => \N__31191\,
            in3 => \N__31091\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => \POWERLED.count_clkZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__31052\,
            in1 => \N__31040\,
            in2 => \N__31007\,
            in3 => \N__31004\,
            lcout => \POWERLED.N_176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__31599\,
            in1 => \N__33545\,
            in2 => \N__33450\,
            in3 => \N__33269\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31490\,
            in2 => \N__31544\,
            in3 => \N__32000\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33555\,
            in1 => \N__31540\,
            in2 => \N__31520\,
            in3 => \N__33270\,
            lcout => \VPP_VDDQ.count_2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__33393\,
            in1 => \N__33547\,
            in2 => \N__31603\,
            in3 => \N__33273\,
            lcout => \VPP_VDDQ.curr_state_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33127\,
            ce => \N__31772\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33271\,
            in1 => \N__33556\,
            in2 => \N__31483\,
            in3 => \N__33391\,
            lcout => \VPP_VDDQ.count_2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33392\,
            in1 => \N__33546\,
            in2 => \N__32285\,
            in3 => \N__33272\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI7EJU_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32362\,
            in1 => \_gnd_net_\,
            in2 => \N__31451\,
            in3 => \N__32267\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__31433\,
            in1 => \N__33615\,
            in2 => \N__31660\,
            in3 => \N__31677\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33135\,
            ce => \N__31771\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33429\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33207\,
            lcout => \VPP_VDDQ.N_385\,
            ltout => \VPP_VDDQ.N_385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__31653\,
            in1 => \N__33616\,
            in2 => \N__31427\,
            in3 => \N__31678\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.m4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32018\,
            in2 => \N__32012\,
            in3 => \N__32009\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__31595\,
            in1 => \N__31676\,
            in2 => \N__31805\,
            in3 => \N__31794\,
            lcout => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIDNMU_6_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31685\,
            in2 => \N__31706\,
            in3 => \N__32243\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33208\,
            in1 => \N__33430\,
            in2 => \N__32258\,
            in3 => \N__33617\,
            lcout => \VPP_VDDQ.count_2_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_a2_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31679\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31654\,
            lcout => \N_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__33432\,
            in1 => \N__32137\,
            in2 => \N__33618\,
            in3 => \N__33236\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIL8AN_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32114\,
            in2 => \N__31577\,
            in3 => \N__32331\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__32333\,
            in1 => \N__31573\,
            in2 => \N__32090\,
            in3 => \N__32096\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIQODG5_10_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32183\,
            in1 => \N__31559\,
            in2 => \N__31553\,
            in3 => \N__31550\,
            lcout => \VPP_VDDQ.N_1_i\,
            ltout => \VPP_VDDQ.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_0_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__33434\,
            in1 => \N__33656\,
            in2 => \N__32153\,
            in3 => \N__32136\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33141\,
            ce => \N__32403\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33238\,
            in1 => \N__33554\,
            in2 => \N__32108\,
            in3 => \N__33435\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33141\,
            ce => \N__32403\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33433\,
            in1 => \N__32104\,
            in2 => \N__33619\,
            in3 => \N__33237\,
            lcout => \VPP_VDDQ.count_2_1_7\,
            ltout => \VPP_VDDQ.count_2_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFQNU_7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32086\,
            in2 => \N__32078\,
            in3 => \N__32332\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33241\,
            in1 => \N__33313\,
            in2 => \N__33662\,
            in3 => \N__33454\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI75M41_12_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32380\,
            in2 => \N__32069\,
            in3 => \N__33152\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33240\,
            in1 => \N__33625\,
            in2 => \N__32057\,
            in3 => \N__33453\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIBBO41_14_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__32039\,
            in1 => \N__32379\,
            in2 => \N__32033\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33242\,
            in1 => \N__32281\,
            in2 => \N__33663\,
            in3 => \N__33456\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33111\,
            ce => \N__32425\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33455\,
            in1 => \N__33244\,
            in2 => \N__33659\,
            in3 => \N__32254\,
            lcout => \VPP_VDDQ.count_2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33111\,
            ce => \N__32425\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33243\,
            in1 => \N__33626\,
            in2 => \N__32219\,
            in3 => \N__33457\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33111\,
            ce => \N__32425\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33452\,
            in1 => \N__33239\,
            in2 => \N__33658\,
            in3 => \N__32218\,
            lcout => \VPP_VDDQ.count_2_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33284\,
            in1 => \N__33703\,
            in2 => \N__33472\,
            in3 => \N__33634\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33146\,
            ce => \N__32409\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33631\,
            in1 => \N__33459\,
            in2 => \N__33298\,
            in3 => \N__32173\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI52L41_11_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32159\,
            in2 => \N__32195\,
            in3 => \N__32377\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => \VPP_VDDQ.count_2Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIS3FU_0_10_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__32378\,
            in1 => \N__33686\,
            in2 => \N__32186\,
            in3 => \N__33692\,
            lcout => \VPP_VDDQ.un9_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33285\,
            in1 => \N__33633\,
            in2 => \N__32174\,
            in3 => \N__33471\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33146\,
            ce => \N__32409\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33630\,
            in1 => \N__33458\,
            in2 => \N__33704\,
            in3 => \N__33283\,
            lcout => \VPP_VDDQ.count_2_1_10\,
            ltout => \VPP_VDDQ.count_2_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIS3FU_10_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33685\,
            in2 => \N__33674\,
            in3 => \N__32376\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33632\,
            in1 => \N__33460\,
            in2 => \N__33314\,
            in3 => \N__33286\,
            lcout => \VPP_VDDQ.count_2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33146\,
            ce => \N__32409\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
