// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 7 2022 11:04:43

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    output SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__34245;
    wire N__34244;
    wire N__34243;
    wire N__34236;
    wire N__34235;
    wire N__34234;
    wire N__34227;
    wire N__34226;
    wire N__34225;
    wire N__34218;
    wire N__34217;
    wire N__34216;
    wire N__34209;
    wire N__34208;
    wire N__34207;
    wire N__34200;
    wire N__34199;
    wire N__34198;
    wire N__34191;
    wire N__34190;
    wire N__34189;
    wire N__34182;
    wire N__34181;
    wire N__34180;
    wire N__34173;
    wire N__34172;
    wire N__34171;
    wire N__34164;
    wire N__34163;
    wire N__34162;
    wire N__34155;
    wire N__34154;
    wire N__34153;
    wire N__34146;
    wire N__34145;
    wire N__34144;
    wire N__34137;
    wire N__34136;
    wire N__34135;
    wire N__34128;
    wire N__34127;
    wire N__34126;
    wire N__34119;
    wire N__34118;
    wire N__34117;
    wire N__34110;
    wire N__34109;
    wire N__34108;
    wire N__34101;
    wire N__34100;
    wire N__34099;
    wire N__34092;
    wire N__34091;
    wire N__34090;
    wire N__34083;
    wire N__34082;
    wire N__34081;
    wire N__34074;
    wire N__34073;
    wire N__34072;
    wire N__34065;
    wire N__34064;
    wire N__34063;
    wire N__34056;
    wire N__34055;
    wire N__34054;
    wire N__34047;
    wire N__34046;
    wire N__34045;
    wire N__34038;
    wire N__34037;
    wire N__34036;
    wire N__34029;
    wire N__34028;
    wire N__34027;
    wire N__34020;
    wire N__34019;
    wire N__34018;
    wire N__34011;
    wire N__34010;
    wire N__34009;
    wire N__34002;
    wire N__34001;
    wire N__34000;
    wire N__33993;
    wire N__33992;
    wire N__33991;
    wire N__33984;
    wire N__33983;
    wire N__33982;
    wire N__33975;
    wire N__33974;
    wire N__33973;
    wire N__33966;
    wire N__33965;
    wire N__33964;
    wire N__33957;
    wire N__33956;
    wire N__33955;
    wire N__33948;
    wire N__33947;
    wire N__33946;
    wire N__33939;
    wire N__33938;
    wire N__33937;
    wire N__33930;
    wire N__33929;
    wire N__33928;
    wire N__33921;
    wire N__33920;
    wire N__33919;
    wire N__33912;
    wire N__33911;
    wire N__33910;
    wire N__33903;
    wire N__33902;
    wire N__33901;
    wire N__33894;
    wire N__33893;
    wire N__33892;
    wire N__33885;
    wire N__33884;
    wire N__33883;
    wire N__33876;
    wire N__33875;
    wire N__33874;
    wire N__33867;
    wire N__33866;
    wire N__33865;
    wire N__33858;
    wire N__33857;
    wire N__33856;
    wire N__33849;
    wire N__33848;
    wire N__33847;
    wire N__33840;
    wire N__33839;
    wire N__33838;
    wire N__33831;
    wire N__33830;
    wire N__33829;
    wire N__33822;
    wire N__33821;
    wire N__33820;
    wire N__33813;
    wire N__33812;
    wire N__33811;
    wire N__33804;
    wire N__33803;
    wire N__33802;
    wire N__33795;
    wire N__33794;
    wire N__33793;
    wire N__33786;
    wire N__33785;
    wire N__33784;
    wire N__33777;
    wire N__33776;
    wire N__33775;
    wire N__33768;
    wire N__33767;
    wire N__33766;
    wire N__33759;
    wire N__33758;
    wire N__33757;
    wire N__33750;
    wire N__33749;
    wire N__33748;
    wire N__33741;
    wire N__33740;
    wire N__33739;
    wire N__33732;
    wire N__33731;
    wire N__33730;
    wire N__33723;
    wire N__33722;
    wire N__33721;
    wire N__33704;
    wire N__33703;
    wire N__33700;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33664;
    wire N__33663;
    wire N__33662;
    wire N__33661;
    wire N__33660;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33655;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33634;
    wire N__33633;
    wire N__33632;
    wire N__33631;
    wire N__33630;
    wire N__33627;
    wire N__33626;
    wire N__33625;
    wire N__33622;
    wire N__33621;
    wire N__33620;
    wire N__33619;
    wire N__33618;
    wire N__33617;
    wire N__33616;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33598;
    wire N__33593;
    wire N__33588;
    wire N__33577;
    wire N__33568;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33560;
    wire N__33559;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33555;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33547;
    wire N__33546;
    wire N__33545;
    wire N__33538;
    wire N__33535;
    wire N__33522;
    wire N__33507;
    wire N__33502;
    wire N__33495;
    wire N__33488;
    wire N__33473;
    wire N__33472;
    wire N__33471;
    wire N__33470;
    wire N__33467;
    wire N__33466;
    wire N__33465;
    wire N__33464;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33455;
    wire N__33454;
    wire N__33453;
    wire N__33452;
    wire N__33451;
    wire N__33450;
    wire N__33447;
    wire N__33436;
    wire N__33435;
    wire N__33434;
    wire N__33433;
    wire N__33432;
    wire N__33431;
    wire N__33430;
    wire N__33429;
    wire N__33428;
    wire N__33419;
    wire N__33406;
    wire N__33403;
    wire N__33402;
    wire N__33401;
    wire N__33400;
    wire N__33399;
    wire N__33398;
    wire N__33397;
    wire N__33394;
    wire N__33393;
    wire N__33392;
    wire N__33391;
    wire N__33386;
    wire N__33377;
    wire N__33374;
    wire N__33369;
    wire N__33366;
    wire N__33361;
    wire N__33346;
    wire N__33337;
    wire N__33332;
    wire N__33329;
    wire N__33314;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33299;
    wire N__33298;
    wire N__33297;
    wire N__33294;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33287;
    wire N__33286;
    wire N__33285;
    wire N__33284;
    wire N__33283;
    wire N__33282;
    wire N__33281;
    wire N__33280;
    wire N__33279;
    wire N__33278;
    wire N__33277;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33257;
    wire N__33254;
    wire N__33245;
    wire N__33244;
    wire N__33243;
    wire N__33242;
    wire N__33241;
    wire N__33240;
    wire N__33239;
    wire N__33238;
    wire N__33237;
    wire N__33236;
    wire N__33225;
    wire N__33220;
    wire N__33209;
    wire N__33208;
    wire N__33207;
    wire N__33204;
    wire N__33197;
    wire N__33184;
    wire N__33177;
    wire N__33170;
    wire N__33165;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33142;
    wire N__33141;
    wire N__33140;
    wire N__33139;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33132;
    wire N__33129;
    wire N__33128;
    wire N__33127;
    wire N__33124;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33113;
    wire N__33112;
    wire N__33111;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33100;
    wire N__33099;
    wire N__33094;
    wire N__33091;
    wire N__33090;
    wire N__33087;
    wire N__33086;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33078;
    wire N__33077;
    wire N__33072;
    wire N__33071;
    wire N__33070;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33066;
    wire N__33063;
    wire N__33060;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33052;
    wire N__33051;
    wire N__33050;
    wire N__33049;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33029;
    wire N__33028;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32989;
    wire N__32986;
    wire N__32985;
    wire N__32982;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32974;
    wire N__32973;
    wire N__32972;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32964;
    wire N__32963;
    wire N__32960;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32949;
    wire N__32948;
    wire N__32945;
    wire N__32944;
    wire N__32943;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32928;
    wire N__32927;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32911;
    wire N__32908;
    wire N__32907;
    wire N__32906;
    wire N__32901;
    wire N__32900;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32888;
    wire N__32887;
    wire N__32884;
    wire N__32879;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32851;
    wire N__32848;
    wire N__32845;
    wire N__32844;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32819;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32798;
    wire N__32795;
    wire N__32794;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32777;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32769;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32748;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32731;
    wire N__32728;
    wire N__32719;
    wire N__32714;
    wire N__32709;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32686;
    wire N__32685;
    wire N__32680;
    wire N__32677;
    wire N__32672;
    wire N__32669;
    wire N__32660;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32640;
    wire N__32635;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32612;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32592;
    wire N__32587;
    wire N__32580;
    wire N__32573;
    wire N__32570;
    wire N__32569;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32548;
    wire N__32541;
    wire N__32534;
    wire N__32529;
    wire N__32526;
    wire N__32521;
    wire N__32512;
    wire N__32507;
    wire N__32504;
    wire N__32493;
    wire N__32490;
    wire N__32489;
    wire N__32482;
    wire N__32479;
    wire N__32472;
    wire N__32467;
    wire N__32460;
    wire N__32455;
    wire N__32452;
    wire N__32449;
    wire N__32446;
    wire N__32429;
    wire N__32426;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32418;
    wire N__32413;
    wire N__32410;
    wire N__32409;
    wire N__32404;
    wire N__32403;
    wire N__32402;
    wire N__32401;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32383;
    wire N__32382;
    wire N__32381;
    wire N__32380;
    wire N__32379;
    wire N__32378;
    wire N__32377;
    wire N__32376;
    wire N__32369;
    wire N__32364;
    wire N__32363;
    wire N__32362;
    wire N__32361;
    wire N__32360;
    wire N__32359;
    wire N__32358;
    wire N__32357;
    wire N__32356;
    wire N__32351;
    wire N__32346;
    wire N__32339;
    wire N__32334;
    wire N__32333;
    wire N__32332;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32312;
    wire N__32303;
    wire N__32296;
    wire N__32285;
    wire N__32282;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32218;
    wire N__32215;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32173;
    wire N__32170;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32138;
    wire N__32137;
    wire N__32136;
    wire N__32135;
    wire N__32132;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32104;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32087;
    wire N__32086;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32065;
    wire N__32060;
    wire N__32057;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32009;
    wire N__32008;
    wire N__32005;
    wire N__32004;
    wire N__32003;
    wire N__32002;
    wire N__32001;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31995;
    wire N__31994;
    wire N__31993;
    wire N__31992;
    wire N__31991;
    wire N__31990;
    wire N__31989;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31943;
    wire N__31938;
    wire N__31931;
    wire N__31928;
    wire N__31921;
    wire N__31916;
    wire N__31913;
    wire N__31908;
    wire N__31901;
    wire N__31896;
    wire N__31891;
    wire N__31890;
    wire N__31889;
    wire N__31886;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31872;
    wire N__31865;
    wire N__31862;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31835;
    wire N__31832;
    wire N__31827;
    wire N__31818;
    wire N__31805;
    wire N__31802;
    wire N__31801;
    wire N__31800;
    wire N__31799;
    wire N__31796;
    wire N__31795;
    wire N__31794;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31772;
    wire N__31771;
    wire N__31770;
    wire N__31769;
    wire N__31768;
    wire N__31767;
    wire N__31766;
    wire N__31765;
    wire N__31764;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31745;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31678;
    wire N__31677;
    wire N__31676;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31660;
    wire N__31659;
    wire N__31658;
    wire N__31655;
    wire N__31654;
    wire N__31653;
    wire N__31650;
    wire N__31643;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31612;
    wire N__31607;
    wire N__31604;
    wire N__31603;
    wire N__31600;
    wire N__31599;
    wire N__31596;
    wire N__31595;
    wire N__31592;
    wire N__31587;
    wire N__31584;
    wire N__31577;
    wire N__31574;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31484;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31460;
    wire N__31459;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31423;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31409;
    wire N__31406;
    wire N__31405;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31348;
    wire N__31347;
    wire N__31346;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31332;
    wire N__31329;
    wire N__31322;
    wire N__31321;
    wire N__31320;
    wire N__31319;
    wire N__31318;
    wire N__31317;
    wire N__31316;
    wire N__31315;
    wire N__31314;
    wire N__31313;
    wire N__31312;
    wire N__31311;
    wire N__31310;
    wire N__31309;
    wire N__31304;
    wire N__31299;
    wire N__31290;
    wire N__31287;
    wire N__31286;
    wire N__31285;
    wire N__31284;
    wire N__31283;
    wire N__31272;
    wire N__31265;
    wire N__31254;
    wire N__31253;
    wire N__31252;
    wire N__31251;
    wire N__31244;
    wire N__31237;
    wire N__31234;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31219;
    wire N__31218;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31207;
    wire N__31206;
    wire N__31205;
    wire N__31204;
    wire N__31203;
    wire N__31202;
    wire N__31201;
    wire N__31198;
    wire N__31193;
    wire N__31192;
    wire N__31191;
    wire N__31188;
    wire N__31183;
    wire N__31174;
    wire N__31171;
    wire N__31166;
    wire N__31163;
    wire N__31162;
    wire N__31161;
    wire N__31160;
    wire N__31157;
    wire N__31152;
    wire N__31149;
    wire N__31148;
    wire N__31147;
    wire N__31146;
    wire N__31145;
    wire N__31144;
    wire N__31143;
    wire N__31136;
    wire N__31131;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31107;
    wire N__31100;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31078;
    wire N__31077;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31052;
    wire N__31051;
    wire N__31048;
    wire N__31045;
    wire N__31040;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31007;
    wire N__31004;
    wire N__31003;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30968;
    wire N__30967;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30935;
    wire N__30932;
    wire N__30931;
    wire N__30930;
    wire N__30929;
    wire N__30926;
    wire N__30925;
    wire N__30924;
    wire N__30923;
    wire N__30922;
    wire N__30921;
    wire N__30920;
    wire N__30919;
    wire N__30918;
    wire N__30917;
    wire N__30916;
    wire N__30915;
    wire N__30914;
    wire N__30913;
    wire N__30912;
    wire N__30911;
    wire N__30910;
    wire N__30903;
    wire N__30894;
    wire N__30889;
    wire N__30888;
    wire N__30877;
    wire N__30864;
    wire N__30863;
    wire N__30862;
    wire N__30861;
    wire N__30860;
    wire N__30859;
    wire N__30858;
    wire N__30857;
    wire N__30856;
    wire N__30855;
    wire N__30854;
    wire N__30853;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30823;
    wire N__30812;
    wire N__30809;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30787;
    wire N__30786;
    wire N__30785;
    wire N__30784;
    wire N__30783;
    wire N__30782;
    wire N__30779;
    wire N__30778;
    wire N__30777;
    wire N__30776;
    wire N__30775;
    wire N__30774;
    wire N__30773;
    wire N__30768;
    wire N__30767;
    wire N__30766;
    wire N__30765;
    wire N__30762;
    wire N__30761;
    wire N__30758;
    wire N__30757;
    wire N__30756;
    wire N__30755;
    wire N__30754;
    wire N__30753;
    wire N__30752;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30735;
    wire N__30734;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30716;
    wire N__30715;
    wire N__30714;
    wire N__30711;
    wire N__30704;
    wire N__30695;
    wire N__30688;
    wire N__30683;
    wire N__30680;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30654;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30632;
    wire N__30623;
    wire N__30620;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30586;
    wire N__30585;
    wire N__30584;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30576;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30555;
    wire N__30554;
    wire N__30551;
    wire N__30550;
    wire N__30549;
    wire N__30548;
    wire N__30547;
    wire N__30546;
    wire N__30543;
    wire N__30536;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30524;
    wire N__30523;
    wire N__30522;
    wire N__30521;
    wire N__30516;
    wire N__30515;
    wire N__30510;
    wire N__30509;
    wire N__30506;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30488;
    wire N__30485;
    wire N__30484;
    wire N__30483;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30465;
    wire N__30458;
    wire N__30453;
    wire N__30448;
    wire N__30441;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30418;
    wire N__30417;
    wire N__30416;
    wire N__30415;
    wire N__30412;
    wire N__30403;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30311;
    wire N__30310;
    wire N__30307;
    wire N__30306;
    wire N__30303;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30280;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30241;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30229;
    wire N__30228;
    wire N__30227;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30188;
    wire N__30185;
    wire N__30184;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30143;
    wire N__30140;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30106;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30085;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30067;
    wire N__30066;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30043;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30031;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30005;
    wire N__30004;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29980;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29944;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29920;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29888;
    wire N__29885;
    wire N__29884;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29857;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29818;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29794;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29762;
    wire N__29761;
    wire N__29758;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29729;
    wire N__29726;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29673;
    wire N__29668;
    wire N__29665;
    wire N__29658;
    wire N__29651;
    wire N__29650;
    wire N__29647;
    wire N__29646;
    wire N__29641;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29624;
    wire N__29621;
    wire N__29620;
    wire N__29619;
    wire N__29618;
    wire N__29617;
    wire N__29616;
    wire N__29611;
    wire N__29608;
    wire N__29601;
    wire N__29598;
    wire N__29591;
    wire N__29590;
    wire N__29589;
    wire N__29588;
    wire N__29587;
    wire N__29586;
    wire N__29585;
    wire N__29584;
    wire N__29583;
    wire N__29582;
    wire N__29581;
    wire N__29580;
    wire N__29579;
    wire N__29578;
    wire N__29577;
    wire N__29576;
    wire N__29575;
    wire N__29574;
    wire N__29573;
    wire N__29572;
    wire N__29571;
    wire N__29570;
    wire N__29569;
    wire N__29568;
    wire N__29567;
    wire N__29566;
    wire N__29565;
    wire N__29564;
    wire N__29563;
    wire N__29562;
    wire N__29561;
    wire N__29560;
    wire N__29559;
    wire N__29558;
    wire N__29557;
    wire N__29556;
    wire N__29555;
    wire N__29554;
    wire N__29553;
    wire N__29552;
    wire N__29551;
    wire N__29550;
    wire N__29549;
    wire N__29548;
    wire N__29547;
    wire N__29546;
    wire N__29545;
    wire N__29544;
    wire N__29543;
    wire N__29542;
    wire N__29541;
    wire N__29540;
    wire N__29539;
    wire N__29530;
    wire N__29521;
    wire N__29512;
    wire N__29505;
    wire N__29500;
    wire N__29491;
    wire N__29484;
    wire N__29475;
    wire N__29468;
    wire N__29459;
    wire N__29450;
    wire N__29441;
    wire N__29436;
    wire N__29427;
    wire N__29422;
    wire N__29417;
    wire N__29416;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29401;
    wire N__29398;
    wire N__29397;
    wire N__29396;
    wire N__29395;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29269;
    wire N__29268;
    wire N__29267;
    wire N__29264;
    wire N__29261;
    wire N__29256;
    wire N__29251;
    wire N__29250;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29242;
    wire N__29239;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29202;
    wire N__29201;
    wire N__29200;
    wire N__29197;
    wire N__29190;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29165;
    wire N__29162;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29152;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29137;
    wire N__29132;
    wire N__29129;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29071;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29053;
    wire N__29050;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29038;
    wire N__29035;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28952;
    wire N__28949;
    wire N__28948;
    wire N__28945;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28918;
    wire N__28915;
    wire N__28910;
    wire N__28907;
    wire N__28906;
    wire N__28901;
    wire N__28898;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28870;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28822;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28735;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28694;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28676;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28633;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28616;
    wire N__28615;
    wire N__28610;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28592;
    wire N__28591;
    wire N__28586;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28561;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28535;
    wire N__28534;
    wire N__28529;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28511;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28478;
    wire N__28475;
    wire N__28474;
    wire N__28473;
    wire N__28472;
    wire N__28471;
    wire N__28470;
    wire N__28467;
    wire N__28466;
    wire N__28463;
    wire N__28462;
    wire N__28461;
    wire N__28460;
    wire N__28457;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28449;
    wire N__28448;
    wire N__28447;
    wire N__28446;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28429;
    wire N__28428;
    wire N__28425;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28368;
    wire N__28365;
    wire N__28360;
    wire N__28349;
    wire N__28346;
    wire N__28341;
    wire N__28340;
    wire N__28337;
    wire N__28332;
    wire N__28329;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28315;
    wire N__28314;
    wire N__28313;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28286;
    wire N__28283;
    wire N__28282;
    wire N__28281;
    wire N__28274;
    wire N__28271;
    wire N__28270;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28242;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28221;
    wire N__28218;
    wire N__28211;
    wire N__28208;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28178;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28160;
    wire N__28159;
    wire N__28158;
    wire N__28157;
    wire N__28156;
    wire N__28153;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28135;
    wire N__28124;
    wire N__28121;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28076;
    wire N__28073;
    wire N__28072;
    wire N__28069;
    wire N__28068;
    wire N__28067;
    wire N__28066;
    wire N__28065;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28055;
    wire N__28054;
    wire N__28053;
    wire N__28052;
    wire N__28049;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28031;
    wire N__28030;
    wire N__28029;
    wire N__28028;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28010;
    wire N__28005;
    wire N__28002;
    wire N__28001;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27983;
    wire N__27980;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27965;
    wire N__27962;
    wire N__27957;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27931;
    wire N__27926;
    wire N__27919;
    wire N__27914;
    wire N__27909;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27889;
    wire N__27886;
    wire N__27885;
    wire N__27884;
    wire N__27883;
    wire N__27882;
    wire N__27881;
    wire N__27880;
    wire N__27877;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27860;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27845;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27832;
    wire N__27827;
    wire N__27824;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27800;
    wire N__27799;
    wire N__27798;
    wire N__27797;
    wire N__27796;
    wire N__27795;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27783;
    wire N__27780;
    wire N__27779;
    wire N__27778;
    wire N__27777;
    wire N__27776;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27768;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27756;
    wire N__27749;
    wire N__27744;
    wire N__27741;
    wire N__27740;
    wire N__27739;
    wire N__27738;
    wire N__27737;
    wire N__27736;
    wire N__27735;
    wire N__27734;
    wire N__27733;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27694;
    wire N__27685;
    wire N__27678;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27631;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27607;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27509;
    wire N__27506;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27491;
    wire N__27488;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27473;
    wire N__27470;
    wire N__27469;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27461;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27453;
    wire N__27450;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27410;
    wire N__27405;
    wire N__27400;
    wire N__27397;
    wire N__27392;
    wire N__27387;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27338;
    wire N__27335;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27323;
    wire N__27320;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27308;
    wire N__27305;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27293;
    wire N__27290;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27275;
    wire N__27272;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27257;
    wire N__27254;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27149;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27137;
    wire N__27134;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27106;
    wire N__27105;
    wire N__27104;
    wire N__27103;
    wire N__27102;
    wire N__27099;
    wire N__27098;
    wire N__27097;
    wire N__27094;
    wire N__27093;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27081;
    wire N__27078;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27055;
    wire N__27054;
    wire N__27053;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27042;
    wire N__27039;
    wire N__27030;
    wire N__27029;
    wire N__27026;
    wire N__27025;
    wire N__27024;
    wire N__27023;
    wire N__27022;
    wire N__27021;
    wire N__27020;
    wire N__27019;
    wire N__27018;
    wire N__27017;
    wire N__27014;
    wire N__27013;
    wire N__27010;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26994;
    wire N__26985;
    wire N__26976;
    wire N__26963;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26941;
    wire N__26940;
    wire N__26939;
    wire N__26938;
    wire N__26937;
    wire N__26934;
    wire N__26933;
    wire N__26932;
    wire N__26929;
    wire N__26924;
    wire N__26923;
    wire N__26922;
    wire N__26921;
    wire N__26918;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26884;
    wire N__26879;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26859;
    wire N__26852;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26828;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26770;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26755;
    wire N__26750;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26711;
    wire N__26708;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26696;
    wire N__26695;
    wire N__26694;
    wire N__26693;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26682;
    wire N__26681;
    wire N__26678;
    wire N__26677;
    wire N__26676;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26655;
    wire N__26652;
    wire N__26647;
    wire N__26644;
    wire N__26627;
    wire N__26626;
    wire N__26623;
    wire N__26622;
    wire N__26619;
    wire N__26614;
    wire N__26613;
    wire N__26608;
    wire N__26607;
    wire N__26606;
    wire N__26603;
    wire N__26602;
    wire N__26601;
    wire N__26600;
    wire N__26599;
    wire N__26596;
    wire N__26591;
    wire N__26588;
    wire N__26579;
    wire N__26578;
    wire N__26577;
    wire N__26576;
    wire N__26575;
    wire N__26574;
    wire N__26569;
    wire N__26568;
    wire N__26567;
    wire N__26566;
    wire N__26565;
    wire N__26564;
    wire N__26559;
    wire N__26556;
    wire N__26555;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26543;
    wire N__26540;
    wire N__26529;
    wire N__26524;
    wire N__26519;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26491;
    wire N__26490;
    wire N__26489;
    wire N__26488;
    wire N__26487;
    wire N__26484;
    wire N__26483;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26475;
    wire N__26472;
    wire N__26463;
    wire N__26462;
    wire N__26459;
    wire N__26458;
    wire N__26457;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26426;
    wire N__26417;
    wire N__26412;
    wire N__26405;
    wire N__26402;
    wire N__26401;
    wire N__26398;
    wire N__26397;
    wire N__26396;
    wire N__26395;
    wire N__26394;
    wire N__26393;
    wire N__26392;
    wire N__26391;
    wire N__26390;
    wire N__26389;
    wire N__26388;
    wire N__26387;
    wire N__26384;
    wire N__26383;
    wire N__26382;
    wire N__26381;
    wire N__26380;
    wire N__26377;
    wire N__26372;
    wire N__26367;
    wire N__26364;
    wire N__26359;
    wire N__26358;
    wire N__26357;
    wire N__26354;
    wire N__26347;
    wire N__26344;
    wire N__26335;
    wire N__26332;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26311;
    wire N__26300;
    wire N__26297;
    wire N__26288;
    wire N__26287;
    wire N__26286;
    wire N__26283;
    wire N__26282;
    wire N__26279;
    wire N__26278;
    wire N__26275;
    wire N__26274;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26266;
    wire N__26265;
    wire N__26260;
    wire N__26253;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26241;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26215;
    wire N__26210;
    wire N__26207;
    wire N__26198;
    wire N__26195;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26191;
    wire N__26190;
    wire N__26185;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26171;
    wire N__26170;
    wire N__26167;
    wire N__26166;
    wire N__26165;
    wire N__26162;
    wire N__26157;
    wire N__26154;
    wire N__26153;
    wire N__26150;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26128;
    wire N__26125;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26098;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26053;
    wire N__26050;
    wire N__26047;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26032;
    wire N__26031;
    wire N__26030;
    wire N__26029;
    wire N__26028;
    wire N__26027;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26003;
    wire N__26002;
    wire N__26001;
    wire N__26000;
    wire N__25997;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25933;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25900;
    wire N__25895;
    wire N__25892;
    wire N__25891;
    wire N__25890;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25878;
    wire N__25871;
    wire N__25870;
    wire N__25869;
    wire N__25866;
    wire N__25865;
    wire N__25862;
    wire N__25855;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25847;
    wire N__25846;
    wire N__25843;
    wire N__25838;
    wire N__25833;
    wire N__25826;
    wire N__25823;
    wire N__25822;
    wire N__25821;
    wire N__25820;
    wire N__25819;
    wire N__25818;
    wire N__25817;
    wire N__25816;
    wire N__25815;
    wire N__25814;
    wire N__25813;
    wire N__25812;
    wire N__25811;
    wire N__25810;
    wire N__25809;
    wire N__25806;
    wire N__25805;
    wire N__25802;
    wire N__25801;
    wire N__25798;
    wire N__25797;
    wire N__25794;
    wire N__25793;
    wire N__25788;
    wire N__25783;
    wire N__25782;
    wire N__25775;
    wire N__25768;
    wire N__25767;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25759;
    wire N__25758;
    wire N__25757;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25742;
    wire N__25739;
    wire N__25738;
    wire N__25735;
    wire N__25734;
    wire N__25733;
    wire N__25732;
    wire N__25729;
    wire N__25728;
    wire N__25727;
    wire N__25724;
    wire N__25723;
    wire N__25722;
    wire N__25719;
    wire N__25718;
    wire N__25717;
    wire N__25712;
    wire N__25707;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25691;
    wire N__25680;
    wire N__25677;
    wire N__25668;
    wire N__25665;
    wire N__25660;
    wire N__25657;
    wire N__25652;
    wire N__25649;
    wire N__25644;
    wire N__25637;
    wire N__25628;
    wire N__25623;
    wire N__25604;
    wire N__25603;
    wire N__25598;
    wire N__25597;
    wire N__25596;
    wire N__25595;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25580;
    wire N__25579;
    wire N__25578;
    wire N__25573;
    wire N__25568;
    wire N__25563;
    wire N__25556;
    wire N__25553;
    wire N__25548;
    wire N__25541;
    wire N__25538;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25511;
    wire N__25508;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25471;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25436;
    wire N__25433;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25412;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25391;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25379;
    wire N__25376;
    wire N__25375;
    wire N__25372;
    wire N__25369;
    wire N__25364;
    wire N__25361;
    wire N__25360;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25348;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25333;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25321;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25249;
    wire N__25248;
    wire N__25247;
    wire N__25244;
    wire N__25237;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25219;
    wire N__25218;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25208;
    wire N__25205;
    wire N__25200;
    wire N__25197;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25183;
    wire N__25182;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25170;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25141;
    wire N__25140;
    wire N__25137;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25099;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25084;
    wire N__25079;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25051;
    wire N__25046;
    wire N__25045;
    wire N__25044;
    wire N__25043;
    wire N__25042;
    wire N__25041;
    wire N__25040;
    wire N__25039;
    wire N__25038;
    wire N__25037;
    wire N__25036;
    wire N__25035;
    wire N__25034;
    wire N__25033;
    wire N__25032;
    wire N__25031;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25014;
    wire N__25005;
    wire N__24998;
    wire N__24989;
    wire N__24986;
    wire N__24981;
    wire N__24972;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24955;
    wire N__24954;
    wire N__24953;
    wire N__24952;
    wire N__24951;
    wire N__24950;
    wire N__24947;
    wire N__24946;
    wire N__24943;
    wire N__24942;
    wire N__24935;
    wire N__24930;
    wire N__24923;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24911;
    wire N__24908;
    wire N__24907;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24895;
    wire N__24890;
    wire N__24887;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24862;
    wire N__24857;
    wire N__24854;
    wire N__24853;
    wire N__24850;
    wire N__24849;
    wire N__24846;
    wire N__24845;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24821;
    wire N__24816;
    wire N__24809;
    wire N__24808;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24781;
    wire N__24780;
    wire N__24779;
    wire N__24778;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24733;
    wire N__24728;
    wire N__24725;
    wire N__24724;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24698;
    wire N__24695;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24683;
    wire N__24680;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24668;
    wire N__24665;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24572;
    wire N__24569;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24488;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24428;
    wire N__24425;
    wire N__24424;
    wire N__24423;
    wire N__24422;
    wire N__24421;
    wire N__24420;
    wire N__24417;
    wire N__24416;
    wire N__24415;
    wire N__24414;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24406;
    wire N__24403;
    wire N__24402;
    wire N__24399;
    wire N__24398;
    wire N__24395;
    wire N__24394;
    wire N__24389;
    wire N__24388;
    wire N__24387;
    wire N__24386;
    wire N__24383;
    wire N__24378;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24358;
    wire N__24357;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24345;
    wire N__24344;
    wire N__24343;
    wire N__24342;
    wire N__24339;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24323;
    wire N__24318;
    wire N__24311;
    wire N__24302;
    wire N__24295;
    wire N__24284;
    wire N__24283;
    wire N__24282;
    wire N__24281;
    wire N__24280;
    wire N__24279;
    wire N__24276;
    wire N__24271;
    wire N__24270;
    wire N__24269;
    wire N__24268;
    wire N__24267;
    wire N__24266;
    wire N__24265;
    wire N__24264;
    wire N__24263;
    wire N__24260;
    wire N__24255;
    wire N__24250;
    wire N__24249;
    wire N__24248;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24218;
    wire N__24213;
    wire N__24206;
    wire N__24203;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24168;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24160;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24156;
    wire N__24153;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24136;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24107;
    wire N__24106;
    wire N__24105;
    wire N__24104;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24087;
    wire N__24084;
    wire N__24083;
    wire N__24082;
    wire N__24081;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24020;
    wire N__24019;
    wire N__24014;
    wire N__24013;
    wire N__24012;
    wire N__24011;
    wire N__24010;
    wire N__24009;
    wire N__24008;
    wire N__24005;
    wire N__24004;
    wire N__24001;
    wire N__23996;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23976;
    wire N__23975;
    wire N__23974;
    wire N__23971;
    wire N__23966;
    wire N__23961;
    wire N__23954;
    wire N__23953;
    wire N__23952;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23947;
    wire N__23946;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23905;
    wire N__23904;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23893;
    wire N__23892;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23884;
    wire N__23883;
    wire N__23882;
    wire N__23879;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23852;
    wire N__23847;
    wire N__23840;
    wire N__23829;
    wire N__23816;
    wire N__23813;
    wire N__23812;
    wire N__23811;
    wire N__23810;
    wire N__23809;
    wire N__23808;
    wire N__23807;
    wire N__23806;
    wire N__23805;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23793;
    wire N__23790;
    wire N__23789;
    wire N__23784;
    wire N__23781;
    wire N__23780;
    wire N__23779;
    wire N__23778;
    wire N__23777;
    wire N__23772;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23758;
    wire N__23757;
    wire N__23752;
    wire N__23743;
    wire N__23742;
    wire N__23741;
    wire N__23740;
    wire N__23739;
    wire N__23738;
    wire N__23737;
    wire N__23734;
    wire N__23729;
    wire N__23722;
    wire N__23717;
    wire N__23712;
    wire N__23707;
    wire N__23704;
    wire N__23703;
    wire N__23700;
    wire N__23699;
    wire N__23696;
    wire N__23695;
    wire N__23688;
    wire N__23683;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23656;
    wire N__23653;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23624;
    wire N__23621;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23609;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23543;
    wire N__23540;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23516;
    wire N__23513;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23492;
    wire N__23489;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23471;
    wire N__23470;
    wire N__23469;
    wire N__23468;
    wire N__23467;
    wire N__23466;
    wire N__23465;
    wire N__23462;
    wire N__23457;
    wire N__23454;
    wire N__23453;
    wire N__23450;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23442;
    wire N__23435;
    wire N__23434;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23422;
    wire N__23417;
    wire N__23414;
    wire N__23409;
    wire N__23406;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23380;
    wire N__23379;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23371;
    wire N__23368;
    wire N__23367;
    wire N__23366;
    wire N__23363;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23344;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23299;
    wire N__23298;
    wire N__23297;
    wire N__23294;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23269;
    wire N__23264;
    wire N__23261;
    wire N__23260;
    wire N__23259;
    wire N__23258;
    wire N__23257;
    wire N__23256;
    wire N__23255;
    wire N__23254;
    wire N__23251;
    wire N__23250;
    wire N__23249;
    wire N__23246;
    wire N__23245;
    wire N__23244;
    wire N__23237;
    wire N__23232;
    wire N__23231;
    wire N__23230;
    wire N__23229;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23217;
    wire N__23214;
    wire N__23209;
    wire N__23204;
    wire N__23201;
    wire N__23194;
    wire N__23191;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23134;
    wire N__23133;
    wire N__23132;
    wire N__23131;
    wire N__23130;
    wire N__23129;
    wire N__23128;
    wire N__23121;
    wire N__23120;
    wire N__23119;
    wire N__23112;
    wire N__23109;
    wire N__23108;
    wire N__23107;
    wire N__23106;
    wire N__23105;
    wire N__23104;
    wire N__23101;
    wire N__23100;
    wire N__23099;
    wire N__23096;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23073;
    wire N__23066;
    wire N__23057;
    wire N__23048;
    wire N__23045;
    wire N__23044;
    wire N__23041;
    wire N__23040;
    wire N__23037;
    wire N__23036;
    wire N__23035;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23023;
    wire N__23022;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23009;
    wire N__23006;
    wire N__23001;
    wire N__22998;
    wire N__22993;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22975;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22939;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22924;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22910;
    wire N__22907;
    wire N__22906;
    wire N__22905;
    wire N__22904;
    wire N__22903;
    wire N__22902;
    wire N__22901;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22884;
    wire N__22881;
    wire N__22880;
    wire N__22879;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22793;
    wire N__22790;
    wire N__22783;
    wire N__22778;
    wire N__22775;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22745;
    wire N__22742;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22709;
    wire N__22708;
    wire N__22705;
    wire N__22704;
    wire N__22701;
    wire N__22696;
    wire N__22691;
    wire N__22688;
    wire N__22687;
    wire N__22686;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22630;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22618;
    wire N__22615;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22603;
    wire N__22598;
    wire N__22595;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22583;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22555;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22520;
    wire N__22519;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22498;
    wire N__22493;
    wire N__22490;
    wire N__22489;
    wire N__22486;
    wire N__22485;
    wire N__22484;
    wire N__22481;
    wire N__22476;
    wire N__22475;
    wire N__22474;
    wire N__22473;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22465;
    wire N__22464;
    wire N__22461;
    wire N__22456;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22440;
    wire N__22437;
    wire N__22432;
    wire N__22429;
    wire N__22424;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22392;
    wire N__22391;
    wire N__22388;
    wire N__22387;
    wire N__22386;
    wire N__22385;
    wire N__22384;
    wire N__22381;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22351;
    wire N__22346;
    wire N__22341;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22285;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22246;
    wire N__22245;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22239;
    wire N__22234;
    wire N__22231;
    wire N__22230;
    wire N__22223;
    wire N__22222;
    wire N__22221;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22172;
    wire N__22171;
    wire N__22170;
    wire N__22169;
    wire N__22166;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22142;
    wire N__22141;
    wire N__22140;
    wire N__22137;
    wire N__22136;
    wire N__22133;
    wire N__22132;
    wire N__22131;
    wire N__22128;
    wire N__22123;
    wire N__22122;
    wire N__22119;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22100;
    wire N__22097;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22076;
    wire N__22073;
    wire N__22072;
    wire N__22069;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22052;
    wire N__22049;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22041;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22030;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22018;
    wire N__22015;
    wire N__22010;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21994;
    wire N__21991;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21973;
    wire N__21970;
    wire N__21965;
    wire N__21962;
    wire N__21961;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21881;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21811;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21794;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21764;
    wire N__21763;
    wire N__21760;
    wire N__21755;
    wire N__21752;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21740;
    wire N__21737;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21640;
    wire N__21639;
    wire N__21636;
    wire N__21631;
    wire N__21630;
    wire N__21629;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21575;
    wire N__21574;
    wire N__21573;
    wire N__21572;
    wire N__21571;
    wire N__21570;
    wire N__21569;
    wire N__21566;
    wire N__21565;
    wire N__21564;
    wire N__21563;
    wire N__21548;
    wire N__21537;
    wire N__21534;
    wire N__21527;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21519;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21508;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21504;
    wire N__21503;
    wire N__21500;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21480;
    wire N__21473;
    wire N__21466;
    wire N__21463;
    wire N__21452;
    wire N__21451;
    wire N__21450;
    wire N__21449;
    wire N__21448;
    wire N__21447;
    wire N__21446;
    wire N__21445;
    wire N__21444;
    wire N__21443;
    wire N__21428;
    wire N__21421;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21361;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21349;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21325;
    wire N__21322;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21244;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21232;
    wire N__21229;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21211;
    wire N__21206;
    wire N__21205;
    wire N__21204;
    wire N__21201;
    wire N__21200;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21168;
    wire N__21163;
    wire N__21158;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21121;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21103;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21088;
    wire N__21085;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21019;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20878;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20839;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20827;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20792;
    wire N__20789;
    wire N__20788;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20731;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20714;
    wire N__20711;
    wire N__20710;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20669;
    wire N__20666;
    wire N__20665;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20641;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20624;
    wire N__20621;
    wire N__20620;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20573;
    wire N__20570;
    wire N__20569;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20476;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20459;
    wire N__20456;
    wire N__20455;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20413;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20374;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20332;
    wire N__20327;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20203;
    wire N__20200;
    wire N__20199;
    wire N__20196;
    wire N__20195;
    wire N__20192;
    wire N__20187;
    wire N__20184;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20152;
    wire N__20149;
    wire N__20148;
    wire N__20145;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20107;
    wire N__20104;
    wire N__20103;
    wire N__20100;
    wire N__20099;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20085;
    wire N__20078;
    wire N__20075;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20047;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19975;
    wire N__19974;
    wire N__19971;
    wire N__19970;
    wire N__19967;
    wire N__19962;
    wire N__19957;
    wire N__19952;
    wire N__19951;
    wire N__19950;
    wire N__19945;
    wire N__19942;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19904;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19880;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19849;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19711;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19651;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19633;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19621;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19595;
    wire N__19592;
    wire N__19591;
    wire N__19588;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19549;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19492;
    wire N__19487;
    wire N__19484;
    wire N__19483;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19465;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19411;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19394;
    wire N__19393;
    wire N__19390;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19342;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19310;
    wire N__19307;
    wire N__19306;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19288;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19271;
    wire N__19268;
    wire N__19267;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19252;
    wire N__19249;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19211;
    wire N__19208;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19196;
    wire N__19193;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19160;
    wire N__19157;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19088;
    wire N__19085;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19073;
    wire N__19070;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19055;
    wire N__19052;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19025;
    wire N__19022;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19010;
    wire N__19007;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18995;
    wire N__18992;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18977;
    wire N__18974;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18962;
    wire N__18959;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18936;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18928;
    wire N__18927;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18893;
    wire N__18890;
    wire N__18883;
    wire N__18882;
    wire N__18881;
    wire N__18880;
    wire N__18879;
    wire N__18876;
    wire N__18867;
    wire N__18860;
    wire N__18857;
    wire N__18850;
    wire N__18845;
    wire N__18842;
    wire N__18841;
    wire N__18840;
    wire N__18833;
    wire N__18830;
    wire N__18829;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18757;
    wire N__18756;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18740;
    wire N__18737;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18722;
    wire N__18719;
    wire N__18718;
    wire N__18717;
    wire N__18716;
    wire N__18715;
    wire N__18714;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18703;
    wire N__18702;
    wire N__18701;
    wire N__18698;
    wire N__18697;
    wire N__18694;
    wire N__18693;
    wire N__18692;
    wire N__18691;
    wire N__18690;
    wire N__18689;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18681;
    wire N__18680;
    wire N__18679;
    wire N__18678;
    wire N__18677;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18666;
    wire N__18665;
    wire N__18664;
    wire N__18663;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18647;
    wire N__18642;
    wire N__18637;
    wire N__18636;
    wire N__18635;
    wire N__18634;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18618;
    wire N__18609;
    wire N__18606;
    wire N__18601;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18577;
    wire N__18570;
    wire N__18567;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18547;
    wire N__18542;
    wire N__18539;
    wire N__18532;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18476;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18391;
    wire N__18388;
    wire N__18387;
    wire N__18384;
    wire N__18383;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18369;
    wire N__18362;
    wire N__18361;
    wire N__18358;
    wire N__18357;
    wire N__18354;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18313;
    wire N__18310;
    wire N__18309;
    wire N__18306;
    wire N__18305;
    wire N__18302;
    wire N__18297;
    wire N__18294;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18268;
    wire N__18265;
    wire N__18264;
    wire N__18261;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18187;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18173;
    wire N__18170;
    wire N__18169;
    wire N__18164;
    wire N__18161;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18136;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18028;
    wire N__18027;
    wire N__18024;
    wire N__18023;
    wire N__18022;
    wire N__18017;
    wire N__18012;
    wire N__18009;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17981;
    wire N__17978;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17785;
    wire N__17780;
    wire N__17779;
    wire N__17778;
    wire N__17777;
    wire N__17774;
    wire N__17769;
    wire N__17766;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17731;
    wire N__17728;
    wire N__17727;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17643;
    wire N__17642;
    wire N__17641;
    wire N__17640;
    wire N__17637;
    wire N__17626;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17596;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17551;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17528;
    wire N__17527;
    wire N__17524;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17500;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17488;
    wire N__17487;
    wire N__17486;
    wire N__17485;
    wire N__17484;
    wire N__17483;
    wire N__17482;
    wire N__17481;
    wire N__17480;
    wire N__17479;
    wire N__17478;
    wire N__17467;
    wire N__17460;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17449;
    wire N__17448;
    wire N__17447;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17414;
    wire N__17409;
    wire N__17396;
    wire N__17395;
    wire N__17394;
    wire N__17393;
    wire N__17392;
    wire N__17391;
    wire N__17390;
    wire N__17389;
    wire N__17388;
    wire N__17387;
    wire N__17386;
    wire N__17385;
    wire N__17384;
    wire N__17383;
    wire N__17382;
    wire N__17381;
    wire N__17380;
    wire N__17379;
    wire N__17378;
    wire N__17377;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17359;
    wire N__17356;
    wire N__17347;
    wire N__17336;
    wire N__17335;
    wire N__17334;
    wire N__17333;
    wire N__17332;
    wire N__17331;
    wire N__17330;
    wire N__17323;
    wire N__17320;
    wire N__17307;
    wire N__17306;
    wire N__17295;
    wire N__17292;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17270;
    wire N__17267;
    wire N__17266;
    wire N__17265;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17249;
    wire N__17246;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17191;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17176;
    wire N__17175;
    wire N__17170;
    wire N__17167;
    wire N__17162;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17147;
    wire N__17144;
    wire N__17143;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17125;
    wire N__17122;
    wire N__17117;
    wire N__17116;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17081;
    wire N__17080;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17054;
    wire N__17053;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__17001;
    wire N__16998;
    wire N__16991;
    wire N__16990;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16946;
    wire N__16943;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16931;
    wire N__16928;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16909;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16892;
    wire N__16891;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16815;
    wire N__16814;
    wire N__16813;
    wire N__16810;
    wire N__16803;
    wire N__16800;
    wire N__16795;
    wire N__16790;
    wire N__16789;
    wire N__16786;
    wire N__16785;
    wire N__16782;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16768;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16747;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16729;
    wire N__16726;
    wire N__16725;
    wire N__16720;
    wire N__16717;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16693;
    wire N__16690;
    wire N__16689;
    wire N__16686;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16515;
    wire N__16514;
    wire N__16513;
    wire N__16510;
    wire N__16503;
    wire N__16500;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16483;
    wire N__16480;
    wire N__16479;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16450;
    wire N__16447;
    wire N__16446;
    wire N__16443;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16310;
    wire N__16307;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16223;
    wire N__16220;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16190;
    wire N__16187;
    wire N__16186;
    wire N__16185;
    wire N__16184;
    wire N__16183;
    wire N__16182;
    wire N__16177;
    wire N__16168;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16120;
    wire N__16119;
    wire N__16118;
    wire N__16117;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16099;
    wire N__16092;
    wire N__16089;
    wire N__16084;
    wire N__16079;
    wire N__16076;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16068;
    wire N__16067;
    wire N__16062;
    wire N__16057;
    wire N__16054;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15982;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15952;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15910;
    wire N__15907;
    wire N__15902;
    wire N__15899;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15868;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15840;
    wire N__15837;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15820;
    wire N__15817;
    wire N__15816;
    wire N__15813;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15670;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15595;
    wire N__15594;
    wire N__15591;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15557;
    wire N__15556;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15538;
    wire N__15533;
    wire N__15530;
    wire N__15529;
    wire N__15528;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15439;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15431;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15404;
    wire N__15403;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15385;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15179;
    wire N__15176;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15161;
    wire N__15158;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15146;
    wire N__15143;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15128;
    wire N__15125;
    wire N__15124;
    wire N__15121;
    wire N__15118;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15095;
    wire N__15092;
    wire N__15091;
    wire N__15088;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15071;
    wire N__15068;
    wire N__15067;
    wire N__15064;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15047;
    wire N__15044;
    wire N__15043;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15020;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14984;
    wire N__14981;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14969;
    wire N__14966;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14954;
    wire N__14951;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14939;
    wire N__14936;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14924;
    wire N__14921;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14909;
    wire N__14906;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14891;
    wire N__14888;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14876;
    wire N__14873;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14861;
    wire N__14858;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14843;
    wire N__14840;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14828;
    wire N__14825;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14813;
    wire N__14810;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14795;
    wire N__14792;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14780;
    wire N__14777;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14765;
    wire N__14762;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14750;
    wire N__14747;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14725;
    wire N__14724;
    wire N__14723;
    wire N__14720;
    wire N__14713;
    wire N__14708;
    wire N__14705;
    wire N__14704;
    wire N__14703;
    wire N__14700;
    wire N__14695;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14674;
    wire N__14671;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14659;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14638;
    wire N__14635;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14558;
    wire N__14555;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14543;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14531;
    wire N__14528;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14513;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14494;
    wire N__14489;
    wire N__14486;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14474;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14462;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14447;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14413;
    wire N__14412;
    wire N__14409;
    wire N__14406;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14375;
    wire N__14372;
    wire N__14371;
    wire N__14370;
    wire N__14369;
    wire N__14366;
    wire N__14361;
    wire N__14358;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14330;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14318;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14306;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14291;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14279;
    wire N__14278;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14252;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14240;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14225;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14197;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14187;
    wire N__14184;
    wire N__14179;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14068;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14050;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13975;
    wire N__13974;
    wire N__13973;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13961;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13949;
    wire N__13946;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13849;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13773;
    wire N__13772;
    wire N__13769;
    wire N__13764;
    wire N__13761;
    wire N__13754;
    wire N__13751;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13723;
    wire N__13720;
    wire N__13719;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13691;
    wire N__13688;
    wire N__13687;
    wire N__13686;
    wire N__13685;
    wire N__13684;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13660;
    wire N__13659;
    wire N__13658;
    wire N__13657;
    wire N__13646;
    wire N__13643;
    wire N__13642;
    wire N__13641;
    wire N__13638;
    wire N__13637;
    wire N__13636;
    wire N__13627;
    wire N__13624;
    wire N__13619;
    wire N__13616;
    wire N__13615;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13591;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire VCCG0;
    wire bfn_1_2_0_;
    wire \DSW_PWRGD.un1_count_1_cry_0 ;
    wire \DSW_PWRGD.un1_count_1_cry_1 ;
    wire \DSW_PWRGD.un1_count_1_cry_2 ;
    wire \DSW_PWRGD.un1_count_1_cry_3 ;
    wire \DSW_PWRGD.un1_count_1_cry_4 ;
    wire \DSW_PWRGD.un1_count_1_cry_5 ;
    wire \DSW_PWRGD.un1_count_1_cry_6 ;
    wire \DSW_PWRGD.un1_count_1_cry_7 ;
    wire bfn_1_3_0_;
    wire \DSW_PWRGD.un1_count_1_cry_8 ;
    wire \DSW_PWRGD.un1_count_1_cry_9 ;
    wire \DSW_PWRGD.un1_count_1_cry_10 ;
    wire \DSW_PWRGD.un1_count_1_cry_11 ;
    wire \DSW_PWRGD.un1_count_1_cry_12 ;
    wire \DSW_PWRGD.un1_count_1_cry_13 ;
    wire \DSW_PWRGD.un1_count_1_cry_14 ;
    wire \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_1_4_0_;
    wire \DSW_PWRGD.un1_curr_state10_0 ;
    wire v33dsw_ok;
    wire \DSW_PWRGD.curr_stateZ0Z_1 ;
    wire \DSW_PWRGD.curr_stateZ0Z_0 ;
    wire DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_;
    wire G_27;
    wire G_27_cascade_;
    wire \DSW_PWRGD.N_27_1 ;
    wire bfn_1_10_0_;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire bfn_1_11_0_;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_s_8_cascade_ ;
    wire bfn_1_12_0_;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_7_l_fx ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_axb_4_l_fx ;
    wire bfn_1_13_0_;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un124_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire bfn_1_14_0_;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire bfn_1_15_0_;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire bfn_1_16_0_;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire \PCH_PWRGD.count_rst_6_cascade_ ;
    wire \PCH_PWRGD.count_rst_14_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.count_RNIZ0Z_1 ;
    wire \PCH_PWRGD.count_RNIZ0Z_1_cascade_ ;
    wire \PCH_PWRGD.count_0_1 ;
    wire \DSW_PWRGD.countZ0Z_3 ;
    wire \DSW_PWRGD.countZ0Z_4 ;
    wire \DSW_PWRGD.countZ0Z_0 ;
    wire \DSW_PWRGD.countZ0Z_1 ;
    wire \PCH_PWRGD.delayed_vccin_ok_0 ;
    wire \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0_cascade_ ;
    wire \DSW_PWRGD.countZ0Z_11 ;
    wire \DSW_PWRGD.countZ0Z_10 ;
    wire \DSW_PWRGD.countZ0Z_6 ;
    wire \DSW_PWRGD.countZ0Z_5 ;
    wire \DSW_PWRGD.countZ0Z_9 ;
    wire \DSW_PWRGD.countZ0Z_7 ;
    wire \DSW_PWRGD.countZ0Z_8 ;
    wire \DSW_PWRGD.countZ0Z_2 ;
    wire \PCH_PWRGD.N_2126_i_cascade_ ;
    wire \PCH_PWRGD.N_381_cascade_ ;
    wire \PCH_PWRGD.N_254_0 ;
    wire \DSW_PWRGD.countZ0Z_12 ;
    wire \DSW_PWRGD.countZ0Z_13 ;
    wire \DSW_PWRGD.countZ0Z_14 ;
    wire \DSW_PWRGD.countZ0Z_15 ;
    wire \DSW_PWRGD.un4_count_11 ;
    wire \DSW_PWRGD.un4_count_10 ;
    wire \DSW_PWRGD.un4_count_8_cascade_ ;
    wire \DSW_PWRGD.un4_count_9 ;
    wire \DSW_PWRGD.N_1_i ;
    wire \PCH_PWRGD.N_381 ;
    wire \PCH_PWRGD.N_2126_i ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.N_255_0_cascade_ ;
    wire \COUNTER.counterZ0Z_0 ;
    wire bfn_2_5_0_;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire bfn_2_6_0_;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire bfn_2_7_0_;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire bfn_2_8_0_;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \POWERLED.un1_count_cry_0_i ;
    wire bfn_2_9_0_;
    wire \POWERLED.N_4527_i ;
    wire \POWERLED.un85_clk_100khz_cry_0 ;
    wire \POWERLED.N_4528_i ;
    wire \POWERLED.un85_clk_100khz_cry_1 ;
    wire \POWERLED.un85_clk_100khz_3 ;
    wire \POWERLED.N_4529_i ;
    wire \POWERLED.un85_clk_100khz_cry_2 ;
    wire \POWERLED.un85_clk_100khz_4 ;
    wire \POWERLED.N_4530_i ;
    wire \POWERLED.un85_clk_100khz_cry_3 ;
    wire \POWERLED.N_4531_i ;
    wire \POWERLED.un85_clk_100khz_cry_4 ;
    wire \POWERLED.un85_clk_100khz_6 ;
    wire \POWERLED.N_4532_i ;
    wire \POWERLED.un85_clk_100khz_cry_5 ;
    wire \POWERLED.N_4533_i ;
    wire \POWERLED.un85_clk_100khz_cry_6 ;
    wire \POWERLED.un85_clk_100khz_cry_7 ;
    wire \POWERLED.N_4534_i ;
    wire bfn_2_10_0_;
    wire \POWERLED.N_4535_i ;
    wire \POWERLED.un85_clk_100khz_cry_8 ;
    wire \POWERLED.N_4536_i ;
    wire \POWERLED.un85_clk_100khz_cry_9 ;
    wire \POWERLED.N_4537_i ;
    wire \POWERLED.un85_clk_100khz_cry_10 ;
    wire \POWERLED.N_4538_i ;
    wire \POWERLED.un85_clk_100khz_cry_11 ;
    wire \POWERLED.N_4539_i ;
    wire \POWERLED.un85_clk_100khz_cry_12 ;
    wire \POWERLED.N_4540_i ;
    wire \POWERLED.un85_clk_100khz_cry_13 ;
    wire \POWERLED.N_4541_i ;
    wire \POWERLED.un85_clk_100khz_cry_14 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_2_11_0_;
    wire \POWERLED.un85_clk_100khz_1 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.un85_clk_100khz_9 ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.un85_clk_100khz_5 ;
    wire \POWERLED.un85_clk_100khz_11 ;
    wire v33a_enn;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.un85_clk_100khz_13 ;
    wire \POWERLED.un85_clk_100khz_8 ;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.un85_clk_100khz_7 ;
    wire \POWERLED.un85_clk_100khz_12 ;
    wire \POWERLED.mult1_un61_sum_i_8 ;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire \POWERLED.un85_clk_100khz_14 ;
    wire vpp_ok;
    wire vddq_en;
    wire bfn_2_15_0_;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \PCH_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire \PCH_PWRGD.m4_0_0_cascade_ ;
    wire \PCH_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.curr_state_0_1 ;
    wire \PCH_PWRGD.count_0_8 ;
    wire \PCH_PWRGD.countZ0Z_9_cascade_ ;
    wire \PCH_PWRGD.count_rst_6 ;
    wire \PCH_PWRGD.curr_state_RNI3DJUZ0Z_0 ;
    wire \PCH_PWRGD.curr_state_0_0 ;
    wire \PCH_PWRGD.count_rst_11 ;
    wire \PCH_PWRGD.count_rst_11_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_3_cascade_ ;
    wire \PCH_PWRGD.count_0_3 ;
    wire \PCH_PWRGD.count_rst_10_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_4_cascade_ ;
    wire \PCH_PWRGD.count_0_4 ;
    wire \PCH_PWRGD.count_0_0 ;
    wire \PCH_PWRGD.count_rst_3_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_11_cascade_ ;
    wire \PCH_PWRGD.count_rst_3 ;
    wire \PCH_PWRGD.count_0_11 ;
    wire \PCH_PWRGD.un12_clk_100khz_7 ;
    wire \PCH_PWRGD.un12_clk_100khz_4_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_5 ;
    wire \PCH_PWRGD.un12_clk_100khz_13_cascade_ ;
    wire \PCH_PWRGD.N_1_i ;
    wire \PCH_PWRGD.N_1_i_cascade_ ;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2_cascade_ ;
    wire \PCH_PWRGD.curr_state_7_1 ;
    wire \PCH_PWRGD.countZ0Z_15_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_8 ;
    wire \PCH_PWRGD.count_0_14 ;
    wire \PCH_PWRGD.count_0_13 ;
    wire \PCH_PWRGD.count_0_15 ;
    wire N_187_cascade_;
    wire v33a_ok;
    wire v5a_ok;
    wire slp_susn;
    wire v1p8a_ok;
    wire rsmrst_pwrgd_signal_cascade_;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_4_7_0_;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire COUNTER_un4_counter_7;
    wire bfn_4_8_0_;
    wire v5s_enn;
    wire bfn_4_9_0_;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire G_2121;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.un85_clk_100khz_0 ;
    wire \POWERLED.mult1_un159_sum_i ;
    wire bfn_4_10_0_;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.un85_clk_100khz_2 ;
    wire \POWERLED.un2_count_clk_17_0_a2_5_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_46_0_cascade_ ;
    wire bfn_4_13_0_;
    wire \POWERLED.mult1_un47_sum_i ;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un54_sum_s_8_cascade_ ;
    wire bfn_4_14_0_;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8_cascade_ ;
    wire bfn_4_15_0_;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \PCH_PWRGD.un2_count_1_axb_5_cascade_ ;
    wire \PCH_PWRGD.count_0_5 ;
    wire \PCH_PWRGD.un12_clk_100khz_6 ;
    wire \PCH_PWRGD.count_rst_9 ;
    wire \PCH_PWRGD.count_rst_7_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_7_cascade_ ;
    wire \PCH_PWRGD.count_0_7 ;
    wire \PCH_PWRGD.count_0_9 ;
    wire \PCH_PWRGD.countZ0Z_1 ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire bfn_5_2_0_;
    wire \PCH_PWRGD.un2_count_1_cry_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_2 ;
    wire \PCH_PWRGD.countZ0Z_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_3 ;
    wire \PCH_PWRGD.un2_count_1_axb_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_5 ;
    wire \PCH_PWRGD.countZ0Z_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_6 ;
    wire \PCH_PWRGD.un2_count_1_axb_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_8 ;
    wire bfn_5_3_0_;
    wire \PCH_PWRGD.un2_count_1_cry_9 ;
    wire \PCH_PWRGD.un2_count_1_axb_11 ;
    wire \PCH_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_10 ;
    wire \PCH_PWRGD.un2_count_1_cry_11 ;
    wire \PCH_PWRGD.countZ0Z_13 ;
    wire \PCH_PWRGD.count_rst_1 ;
    wire \PCH_PWRGD.un2_count_1_cry_12 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.count_rst_0 ;
    wire \PCH_PWRGD.un2_count_1_cry_13 ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.un2_count_1_cry_14 ;
    wire \PCH_PWRGD.count_rst ;
    wire \PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ;
    wire \PCH_PWRGD.N_386 ;
    wire \PCH_PWRGD.countZ0Z_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire \PCH_PWRGD.count_rst_5 ;
    wire \RSMRST_PWRGD.un4_count_9_cascade_ ;
    wire \RSMRST_PWRGD.N_1_i ;
    wire \RSMRST_PWRGD.un4_count_8 ;
    wire \RSMRST_PWRGD.un4_count_10 ;
    wire \RSMRST_PWRGD.un4_count_11 ;
    wire \POWERLED.g0_i_o3_0_cascade_ ;
    wire \POWERLED.pwm_outZ0 ;
    wire \POWERLED.g0_i_o3_0 ;
    wire pwrbtn_led;
    wire \POWERLED.curr_state_3_0_cascade_ ;
    wire \POWERLED.curr_stateZ0Z_0_cascade_ ;
    wire \POWERLED.count_0_sqmuxa_i_cascade_ ;
    wire \POWERLED.count_RNIZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.count_rst_8 ;
    wire \PCH_PWRGD.count_0_6 ;
    wire \PCH_PWRGD.un2_count_1_axb_10 ;
    wire RSMRST_PWRGD_curr_state_0;
    wire N_187;
    wire G_11_cascade_;
    wire \POWERLED.count_0_4 ;
    wire \POWERLED.count_0_2 ;
    wire \POWERLED.count_0_11 ;
    wire \POWERLED.count_0_3 ;
    wire \POWERLED.count_0_15 ;
    wire \POWERLED.count_0_7 ;
    wire \POWERLED.count_0_8 ;
    wire \POWERLED.count_0_10 ;
    wire bfn_5_10_0_;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum ;
    wire bfn_5_11_0_;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_0_cZ0 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_1_cZ0 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_2_cZ0 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_3_cZ0 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_4_cZ0 ;
    wire \POWERLED.mult1_un103_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_5_cZ0 ;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_7_cZ0 ;
    wire \POWERLED.mult1_un89_sum ;
    wire bfn_5_12_0_;
    wire \POWERLED.un1_dutycycle_53_cry_8_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_9_cZ0 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_10 ;
    wire \POWERLED.un1_dutycycle_53_cry_11 ;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_12 ;
    wire \POWERLED.un1_dutycycle_53_cry_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_15 ;
    wire bfn_5_13_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.CO2_THRU_CO ;
    wire bfn_5_14_0_;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un68_sum_cry_2_c ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_3_c ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_4_c ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_5_c ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6_c ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un82_sum ;
    wire bfn_5_15_0_;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire \PCH_PWRGD.un2_count_1_axb_2 ;
    wire \PCH_PWRGD.count_0_sqmuxa ;
    wire \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSCZ0 ;
    wire \PCH_PWRGD.count_0_2 ;
    wire \PCH_PWRGD.count_rst_12_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.un12_clk_100khz_3 ;
    wire \PCH_PWRGD.count_0_12 ;
    wire \PCH_PWRGD.count_rst_2 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.count_rst_4 ;
    wire \PCH_PWRGD.count_0_10 ;
    wire \PCH_PWRGD.countZ0Z_12_cascade_ ;
    wire \PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0 ;
    wire \PCH_PWRGD.un12_clk_100khz_2 ;
    wire \RSMRST_PWRGD.N_256_i ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire bfn_6_3_0_;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire bfn_6_4_0_;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_6_5_0_;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.N_27_2 ;
    wire G_11;
    wire \POWERLED.un79_clk_100khzlto4_0_cascade_ ;
    wire \POWERLED.un79_clk_100khzlt15_0_cascade_ ;
    wire \POWERLED.pwm_out_1_sqmuxa ;
    wire \POWERLED.un79_clk_100khzlto15_5 ;
    wire \POWERLED.un79_clk_100khzlto15_6_cascade_ ;
    wire \POWERLED.count_RNIZ0Z_15_cascade_ ;
    wire \POWERLED.N_8 ;
    wire bfn_6_7_0_;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.un1_count_cry_1_c_RNIBZ0Z209 ;
    wire \POWERLED.un1_count_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.un1_count_cry_2_c_RNICZ0Z419 ;
    wire \POWERLED.un1_count_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ;
    wire \POWERLED.un1_count_cry_3 ;
    wire \POWERLED.un1_count_cry_4 ;
    wire \POWERLED.un1_count_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59 ;
    wire \POWERLED.un1_count_cry_6 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69 ;
    wire \POWERLED.un1_count_cry_7 ;
    wire \POWERLED.un1_count_cry_8 ;
    wire bfn_6_8_0_;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ;
    wire \POWERLED.un1_count_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7 ;
    wire \POWERLED.un1_count_cry_10 ;
    wire \POWERLED.un1_count_cry_11 ;
    wire \POWERLED.un1_count_cry_12 ;
    wire \POWERLED.un1_count_cry_13 ;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.un1_count_cry_14 ;
    wire \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ;
    wire \POWERLED.count_0_9 ;
    wire \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79 ;
    wire \POWERLED.countZ0Z_9 ;
    wire \POWERLED.dutycycle_eena_1_cascade_ ;
    wire \POWERLED.N_108_f0_1 ;
    wire \POWERLED.N_108_f0_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_0 ;
    wire \POWERLED.dutycycle_eena_0_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_1 ;
    wire \POWERLED.dutycycle_eena_1 ;
    wire \POWERLED.dutycycleZ1Z_2 ;
    wire \POWERLED.func_state_0_sqmuxa_0_o2_xZ0Z1_cascade_ ;
    wire \POWERLED.g1_1_cascade_ ;
    wire \POWERLED.N_300_N_0_cascade_ ;
    wire \POWERLED.N_4548_0 ;
    wire \POWERLED.N_217_N_0 ;
    wire \POWERLED.N_353_0 ;
    wire \POWERLED.dutycycleZ0Z_10_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_14 ;
    wire \POWERLED.N_86_f0_cascade_ ;
    wire \POWERLED.dutycycle_en_11 ;
    wire \POWERLED.dutycycle_en_11_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_14 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_15 ;
    wire \POWERLED.N_2215_i ;
    wire \POWERLED.N_84_f0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_10_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_13 ;
    wire \POWERLED.dutycycleZ1Z_10 ;
    wire \POWERLED.dutycycleZ0Z_2_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_10 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_9_cascade_ ;
    wire \POWERLED.mult1_un47_sum ;
    wire bfn_6_13_0_;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.un1_dutycycle_53_i_29 ;
    wire \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ;
    wire \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ;
    wire \POWERLED.mult1_un47_sum_s_4_sf ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.dutycycle_en_12 ;
    wire \POWERLED.mult1_un75_sum ;
    wire bfn_6_14_0_;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.dutycycle_RNI_11Z0Z_7_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_12 ;
    wire \POWERLED.un1_dutycycle_53_4_1 ;
    wire \POWERLED.dutycycleZ0Z_3_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_45_a0_1 ;
    wire \POWERLED.un1_dutycycle_53_45_a0_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_10_1 ;
    wire \HDA_STRAP.N_14_cascade_ ;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire hda_sdo_atp;
    wire gpio_fpga_soc_1;
    wire \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_ ;
    wire PCH_PWRGD_delayed_vccin_ok;
    wire \HDA_STRAP.curr_state_RNO_0Z0Z_0 ;
    wire \HDA_STRAP.N_5_0 ;
    wire \POWERLED.N_341_cascade_ ;
    wire \POWERLED.dutycycle_1_0_iv_i_a3_1_0_2_cascade_ ;
    wire \POWERLED.N_64 ;
    wire \POWERLED.g0_0_a3_1_cascade_ ;
    wire \POWERLED.g0_3_1 ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_2 ;
    wire \POWERLED.func_state_RNIMQ0FZ0Z_1 ;
    wire \POWERLED.N_309 ;
    wire \POWERLED.func_state_1_m0_1_cascade_ ;
    wire \POWERLED.count_RNI_0_1_cascade_ ;
    wire \POWERLED.dutycycle_1_0_0 ;
    wire \POWERLED.dutycycleZ1Z_0 ;
    wire \POWERLED.dutycycle_1_0_0_cascade_ ;
    wire \POWERLED.dutycycle_eena ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.func_state_RNIG5G37Z0Z_1 ;
    wire \POWERLED.func_state_cascade_ ;
    wire \POWERLED.dutycycle_1_0_1 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7 ;
    wire \POWERLED.count_0_13 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ;
    wire \POWERLED.count_0_5 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ;
    wire \POWERLED.count_0_14 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49 ;
    wire \POWERLED.count_0_6 ;
    wire \POWERLED.dutycycleZ0Z_11_cascade_ ;
    wire \POWERLED.N_148_N_cascade_ ;
    wire \POWERLED.dutycycle_en_10 ;
    wire \POWERLED.dutycycle_en_10_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.un1_func_state25_4_i_a2_1 ;
    wire \POWERLED.N_301_cascade_ ;
    wire \POWERLED.N_341 ;
    wire \POWERLED.count_clk_en_1_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_ ;
    wire \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_cascade_ ;
    wire \POWERLED.func_state_RNIBVNS_1Z0Z_0_cascade_ ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_ns_1 ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ;
    wire \POWERLED.N_171 ;
    wire \POWERLED.N_283 ;
    wire \POWERLED.N_275_0 ;
    wire \POWERLED.dutycycle_set_0_0 ;
    wire \POWERLED.dutycycle_eena_13_0 ;
    wire \POWERLED.dutycycle_set_0_0_cascade_ ;
    wire \POWERLED.dutycycle_0_6 ;
    wire \POWERLED.dutycycleZ0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_0 ;
    wire \POWERLED.d_i3_mux_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_5 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_7 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_3 ;
    wire \POWERLED.dutycycle_RNIZ0Z_5 ;
    wire \POWERLED.un1_dutycycle_53_13_4_1 ;
    wire \POWERLED.un1_dutycycle_53_13_4_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_13_3 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_11 ;
    wire \POWERLED.g0_0_1 ;
    wire bfn_7_12_0_;
    wire \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_0_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_cZ0 ;
    wire bfn_7_13_0_;
    wire \POWERLED.un1_dutycycle_94_cry_8_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ;
    wire \POWERLED.un1_dutycycle_94_cry_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_12 ;
    wire \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_13 ;
    wire \POWERLED.un1_dutycycle_94_cry_14 ;
    wire \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ;
    wire \POWERLED.g0_i_1_cascade_ ;
    wire \POWERLED.g0_i_0 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_13 ;
    wire \POWERLED.dutycycleZ1Z_9 ;
    wire \POWERLED.dutycycle_rst_1 ;
    wire \POWERLED.dutycycleZ0Z_4_cascade_ ;
    wire \POWERLED.g0_1_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_14 ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_0_0_cascade_ ;
    wire \POWERLED.dutycycle_RNIEB706Z0Z_7 ;
    wire \POWERLED.dutycycleZ1Z_7 ;
    wire \POWERLED.dutycycle_RNIEB706Z0Z_7_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ;
    wire \POWERLED.dutycycleZ1Z_6_cascade_ ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_d_0 ;
    wire \POWERLED.N_143_N_cascade_ ;
    wire \POWERLED.dutycycle_en_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ;
    wire \POWERLED.dutycycleZ1Z_8 ;
    wire \HDA_STRAP.un4_count_12 ;
    wire \HDA_STRAP.un4_count_9_cascade_ ;
    wire \HDA_STRAP.un4_count_13 ;
    wire \HDA_STRAP.un4_count_11 ;
    wire \HDA_STRAP.un4_count_10 ;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire \HDA_STRAP.un4_count ;
    wire \POWERLED.func_state_1_m2s2_i_0 ;
    wire \POWERLED.func_state_1_m2s2_i_1_cascade_ ;
    wire \POWERLED.func_state_1_m0_0_1_0 ;
    wire \POWERLED.count_off_RNIZ0Z_11_cascade_ ;
    wire \POWERLED.N_310 ;
    wire \POWERLED.N_314_cascade_ ;
    wire \POWERLED.count_off_RNIZ0Z_11 ;
    wire \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_ ;
    wire \POWERLED.func_state_RNIHDGK3_0Z0Z_1 ;
    wire \POWERLED.N_67 ;
    wire \POWERLED.func_state_1_m0_0 ;
    wire \POWERLED.func_state_RNIHDGK3_0Z0Z_1_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_o_N_287_N ;
    wire \POWERLED.func_state_RNI_1Z0Z_0 ;
    wire \POWERLED.func_state_RNI_1Z0Z_0_cascade_ ;
    wire \POWERLED.func_state_RNIBK1UZ0Z_0 ;
    wire \POWERLED.N_326_0 ;
    wire \POWERLED.func_stateZ1Z_0 ;
    wire \POWERLED.func_state_RNIB74H7Z0Z_1 ;
    wire \POWERLED.func_state_RNI6RANZ0Z_1 ;
    wire \POWERLED.func_stateZ0Z_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ;
    wire \POWERLED.N_275_cascade_ ;
    wire \POWERLED.un1_clk_100khz_48_and_i_o2_2_0_cascade_ ;
    wire \POWERLED.un1_clk_100khz_48_and_i_o2_3_0 ;
    wire \POWERLED.N_197 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.un85_clk_100khz_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7 ;
    wire \POWERLED.count_0_12 ;
    wire \POWERLED.count_clk_0_2 ;
    wire \POWERLED.count_clk_0_13 ;
    wire \POWERLED.count_clk_0_14 ;
    wire \POWERLED.count_clk_0_3 ;
    wire \POWERLED.count_clk_0_4 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_ ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI_10Z0Z_0 ;
    wire \POWERLED.N_337 ;
    wire SUSWARN_N_fast;
    wire \POWERLED.N_390_cascade_ ;
    wire SUSWARN_N_rep1;
    wire \POWERLED.dutycycle_eena_3_0_0_sx_cascade_ ;
    wire slp_s3n;
    wire rsmrstn;
    wire \POWERLED.N_222 ;
    wire \POWERLED.un1_dutycycle_172_sm3 ;
    wire \POWERLED.un1_clk_100khz_52_and_i_m2_1 ;
    wire \POWERLED.un1_dutycycle_172_m4_cascade_ ;
    wire \POWERLED.un1_clk_100khz_52_and_i_0Z0Z_0 ;
    wire \POWERLED.N_225_cascade_ ;
    wire \POWERLED.dutycycle_eena_14_cascade_ ;
    wire \POWERLED.dutycycle_eena_14 ;
    wire \POWERLED.dutycycle_set_1 ;
    wire \POWERLED.dutycycle_0_5 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ;
    wire \POWERLED.dutycycleZ1Z_3 ;
    wire \POWERLED.dutycycleZ0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_3 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_3 ;
    wire \POWERLED.un1_dutycycle_53_13_2 ;
    wire \POWERLED.un1_dutycycle_53_31_4_1 ;
    wire \POWERLED.dutycycle_en_8 ;
    wire \POWERLED.dutycycle_eena_3_0_1 ;
    wire \POWERLED.dutycycle_eena_3_d_0 ;
    wire \POWERLED.dutycycle_en_3 ;
    wire \POWERLED.un1_dutycycle_53_10_1_0_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_10_1_0 ;
    wire \POWERLED.un2_count_clk_17_0_a2_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ;
    wire \POWERLED.dutycycle_RNI4VJH7Z0Z_4 ;
    wire \POWERLED.dutycycleZ1Z_4 ;
    wire \POWERLED.dutycycleZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.dutycycle_RNI_11Z0Z_7 ;
    wire \POWERLED.un1_dutycycle_53_50_a0_1 ;
    wire \POWERLED.un1_dutycycle_53_2_1_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ;
    wire \POWERLED.dutycycleZ1Z_11 ;
    wire \POWERLED.N_209_iZ0 ;
    wire \POWERLED.un1_dutycycle_53_31_a7_0 ;
    wire \POWERLED.N_144_N_cascade_ ;
    wire \POWERLED.dutycycle_en_7 ;
    wire \POWERLED.count_clk_RNIBVNSZ0Z_4_cascade_ ;
    wire \POWERLED.dutycycle_eena_2 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_7_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_50_3 ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.un1_dutycycle_53_51_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_50_4 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_15 ;
    wire \POWERLED.func_state_RNIBVNSZ0Z_1 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_1 ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_7 ;
    wire \POWERLED.N_8_1 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_3 ;
    wire \POWERLED.dutycycleZ1Z_6 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.g0_i_a6_0_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_12 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.func_state_RNIC4OR2Z0Z_0 ;
    wire \POWERLED.N_390 ;
    wire \POWERLED.N_209 ;
    wire \POWERLED.N_145_N_cascade_ ;
    wire G_154;
    wire \POWERLED.dutycycle_en_9 ;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire \HDA_STRAP.curr_state_RNIH91AZ0Z_1 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_0 ;
    wire bfn_9_1_0_;
    wire \HDA_STRAP.countZ0Z_1 ;
    wire \HDA_STRAP.un1_count_1_cry_0 ;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.un1_count_1_cry_1 ;
    wire \HDA_STRAP.countZ0Z_3 ;
    wire \HDA_STRAP.un1_count_1_cry_2 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.un1_count_1_cry_3 ;
    wire \HDA_STRAP.countZ0Z_5 ;
    wire \HDA_STRAP.un1_count_1_cry_4 ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_6 ;
    wire \HDA_STRAP.un1_count_1_cry_5 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.un1_count_1_cry_6 ;
    wire \HDA_STRAP.un1_count_1_cry_7 ;
    wire \HDA_STRAP.countZ0Z_8 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_8 ;
    wire bfn_9_2_0_;
    wire \HDA_STRAP.countZ0Z_9 ;
    wire \HDA_STRAP.un1_count_1_cry_8 ;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_10 ;
    wire \HDA_STRAP.un1_count_1_cry_9 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_11 ;
    wire \HDA_STRAP.un1_count_1_cry_10 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.un1_count_1_cry_11 ;
    wire \HDA_STRAP.countZ0Z_13 ;
    wire \HDA_STRAP.un1_count_1_cry_12 ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.un1_count_1_cry_13 ;
    wire \HDA_STRAP.countZ0Z_15 ;
    wire \HDA_STRAP.un1_count_1_cry_14 ;
    wire \HDA_STRAP.un1_count_1_cry_15 ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_16 ;
    wire bfn_9_3_0_;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \HDA_STRAP.un1_count_1_cry_16 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_17 ;
    wire \POWERLED.un1_func_state25_6_0_a2_1 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_305_N_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_0_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_1 ;
    wire \POWERLED.N_150_i ;
    wire \POWERLED.N_154 ;
    wire \POWERLED.N_389 ;
    wire \POWERLED.count_off_0_10 ;
    wire \POWERLED.count_off_1_9 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_offZ0Z_10_cascade_ ;
    wire \POWERLED.un34_clk_100khz_4_cascade_ ;
    wire \POWERLED.un34_clk_100khz_5 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire \POWERLED.count_RNIZ0Z_15 ;
    wire \POWERLED.curr_state_1_0 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_1_cascade_ ;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.count_0_1 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.count_0_sqmuxa_i ;
    wire \POWERLED.count_0_0 ;
    wire slp_s4n;
    wire RSMRST_PWRGD_RSMRSTn_2_fast;
    wire \POWERLED.count_clk_0_5 ;
    wire \POWERLED.count_clk_0_6 ;
    wire \POWERLED.count_clk_0_8 ;
    wire \POWERLED.count_clk_0_9 ;
    wire bfn_9_7_0_;
    wire \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_1 ;
    wire \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_2 ;
    wire \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_3 ;
    wire \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_4 ;
    wire \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_5 ;
    wire \POWERLED.un1_count_clk_2_cry_6 ;
    wire \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_7_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_8_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ;
    wire bfn_9_8_0_;
    wire \POWERLED.un1_count_clk_2_cry_9_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_10_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_11 ;
    wire \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_12 ;
    wire \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_13 ;
    wire \POWERLED.un1_count_clk_2_cry_14 ;
    wire \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ;
    wire \POWERLED.count_clk_0_15 ;
    wire \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ;
    wire \POWERLED.count_clk_0_7 ;
    wire \POWERLED.N_392 ;
    wire \POWERLED.mult1_un40_sum_i_5 ;
    wire \POWERLED.mult1_un47_sum_cry_5_THRU_CO ;
    wire \POWERLED.mult1_un47_sum_s_6 ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire \POWERLED.func_state_RNIBVNS_0Z0Z_0 ;
    wire \POWERLED.un1_dutycycle_172_m4_bm_rn_0_cascade_ ;
    wire \POWERLED.dutycycle_RNIMUFP1Z0Z_2 ;
    wire COUNTER_un4_counter_7_THRU_CO;
    wire G_9;
    wire \POWERLED.un1_dutycycle_172_m4_bm_sn ;
    wire \POWERLED.N_20_i ;
    wire \POWERLED.dutycycle_N_3_mux_0 ;
    wire \POWERLED.un1_count_off_1_sqmuxa_2_0_cascade_ ;
    wire \POWERLED.func_state_RNIBVNS_0Z0Z_1 ;
    wire \POWERLED.N_2171_i ;
    wire \POWERLED.un1_dutycycle_172_m3_ns_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_0 ;
    wire \POWERLED.un1_dutycycle_172_m3 ;
    wire \POWERLED.N_2200_i ;
    wire \POWERLED.un1_dutycycle_96_0_a3_1 ;
    wire \POWERLED.dutycycle ;
    wire \POWERLED.N_327 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_5 ;
    wire \POWERLED.un1_dutycycle_53_axb_3_1_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_2 ;
    wire \POWERLED.N_342 ;
    wire \POWERLED.N_155 ;
    wire \POWERLED.N_336 ;
    wire \POWERLED.dutycycle_RNI_9Z0Z_0 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.un1_i3_mux ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.dutycycleZ1Z_5 ;
    wire \POWERLED.dutycycle_RNIZ0Z_1 ;
    wire \VPP_VDDQ.un6_count_10 ;
    wire \VPP_VDDQ.un6_count_8_cascade_ ;
    wire \VPP_VDDQ.un6_count_11 ;
    wire \VPP_VDDQ.un6_count_9 ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire bfn_9_13_0_;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire bfn_9_14_0_;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_9_15_0_;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \POWERLED.count_off_0_5 ;
    wire \POWERLED.count_off_0_15 ;
    wire \POWERLED.count_off_0_8 ;
    wire \POWERLED.un34_clk_100khz_0_cascade_ ;
    wire \POWERLED.un34_clk_100khz_12 ;
    wire \POWERLED.un34_clk_100khz_1 ;
    wire \POWERLED.count_off_1_6 ;
    wire \POWERLED.count_off_1_6_cascade_ ;
    wire \POWERLED.count_off_1_2 ;
    wire \POWERLED.count_off_1_2_cascade_ ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.count_off_1_7 ;
    wire \POWERLED.count_off_1_7_cascade_ ;
    wire \POWERLED.un34_clk_100khz_3 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_off_1_11 ;
    wire \POWERLED.count_off_1_11_cascade_ ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_0 ;
    wire \POWERLED.func_state_RNI_2Z0Z_1 ;
    wire \POWERLED.N_289_cascade_ ;
    wire \POWERLED.func_state_RNIBVNS_2Z0Z_0 ;
    wire \POWERLED.count_off_RNIG5N6N1Z0Z_11 ;
    wire \POWERLED.func_state_RNI_5Z0Z_1 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_2_tz_0_cascade_ ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_2 ;
    wire \POWERLED.func_state_RNI_2Z0Z_0 ;
    wire gpio_fpga_soc_4;
    wire \POWERLED.un1_func_state25_6_0_o_N_304_N ;
    wire \POWERLED.un1_N_3_mux_0 ;
    wire \POWERLED.func_state ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_2_0 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_3_0 ;
    wire \POWERLED.N_352_cascade_ ;
    wire \POWERLED.N_394 ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ;
    wire \POWERLED.N_2182_i ;
    wire \POWERLED.N_352 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_2_2_cascade_ ;
    wire \POWERLED.count_clk_RNIZ0Z_9 ;
    wire \POWERLED.count_clk_0_10 ;
    wire \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.count_clkZ0Z_10_cascade_ ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_4_cascade_ ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.count_clk_0_0 ;
    wire \POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_1_9_cascade_ ;
    wire \VPP_VDDQ.count_2_0_9 ;
    wire \VPP_VDDQ.count_2Z0Z_1 ;
    wire \VPP_VDDQ.un9_clk_100khz_2 ;
    wire \VPP_VDDQ.un9_clk_100khz_0 ;
    wire \VPP_VDDQ.un9_clk_100khz_1_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_3 ;
    wire \VPP_VDDQ.count_2Z0Z_4 ;
    wire \VPP_VDDQ.count_2_1_4 ;
    wire \VPP_VDDQ.count_2_1_5 ;
    wire \VPP_VDDQ.count_2_1_5_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_5 ;
    wire \VPP_VDDQ.count_2Z0Z_2 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_1 ;
    wire bfn_11_11_0_;
    wire \VPP_VDDQ.un1_count_2_1_axb_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6 ;
    wire \VPP_VDDQ.count_2Z0Z_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ;
    wire bfn_11_12_0_;
    wire \VPP_VDDQ.un1_count_2_1_cry_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ;
    wire \VPP_VDDQ.count_2_1_13_cascade_ ;
    wire \VPP_VDDQ.count_2_0_13 ;
    wire \VPP_VDDQ.count_2Z0Z_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_15 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ;
    wire \VPP_VDDQ.count_2_0_15 ;
    wire vpp_en;
    wire vccst_en;
    wire \VPP_VDDQ.N_360_cascade_ ;
    wire \VPP_VDDQ.N_264_i ;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire \VPP_VDDQ.curr_state_RNITROD7Z0Z_0 ;
    wire \VPP_VDDQ.curr_state_RNITROD7Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.N_27_0 ;
    wire \VPP_VDDQ.N_382 ;
    wire \VPP_VDDQ.N_186 ;
    wire \VPP_VDDQ.N_214 ;
    wire \VPP_VDDQ.un6_count ;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire \VPP_VDDQ.N_360 ;
    wire \VPP_VDDQ.curr_stateZ0Z_0 ;
    wire N_27_g;
    wire \POWERLED.count_off_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.count_off_0_12 ;
    wire \POWERLED.count_off_RNIZ0Z_1 ;
    wire \POWERLED.count_off_0_1 ;
    wire \POWERLED.count_off_0_13 ;
    wire \POWERLED.count_offZ0Z_13_cascade_ ;
    wire \POWERLED.un34_clk_100khz_11 ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire bfn_12_4_0_;
    wire \POWERLED.un3_count_off_1_axb_2 ;
    wire \POWERLED.un3_count_off_1_cry_1_c_RNIN70FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_1 ;
    wire \POWERLED.un3_count_off_1_cry_2 ;
    wire \POWERLED.un3_count_off_1_cry_3 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.un3_count_off_1_cry_4_c_RNIQD3FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_4 ;
    wire \POWERLED.un3_count_off_1_axb_6 ;
    wire \POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_5 ;
    wire \POWERLED.un3_count_off_1_axb_7 ;
    wire \POWERLED.un3_count_off_1_cry_6_c_RNISH5FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_6 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.un3_count_off_1_cry_7_c_RNITJ6FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_7 ;
    wire \POWERLED.un3_count_off_1_cry_8 ;
    wire \POWERLED.un3_count_off_1_axb_9 ;
    wire \POWERLED.un3_count_off_1_cry_8_c_RNIUL7FZ0 ;
    wire bfn_12_5_0_;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.un3_count_off_1_cry_9_c_RNIVN8FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_9 ;
    wire \POWERLED.un3_count_off_1_axb_11 ;
    wire \POWERLED.un3_count_off_1_cry_10_c_RNI7ULDZ0 ;
    wire \POWERLED.un3_count_off_1_cry_10 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.un3_count_off_1_cry_11_c_RNI80NDZ0 ;
    wire \POWERLED.un3_count_off_1_cry_11 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.un3_count_off_1_cry_12_c_RNI92ODZ0 ;
    wire \POWERLED.un3_count_off_1_cry_12 ;
    wire \POWERLED.un3_count_off_1_cry_13 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.un3_count_off_1_cry_14 ;
    wire \POWERLED.un3_count_off_1_cry_14_c_RNIB6QDZ0 ;
    wire \POWERLED.count_off_0_14 ;
    wire \POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.count_offZ0Z_4_cascade_ ;
    wire \POWERLED.un34_clk_100khz_2 ;
    wire \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ;
    wire \POWERLED.count_off_1_3 ;
    wire \POWERLED.count_off_1_3_cascade_ ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.un3_count_off_1_axb_3 ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.count_offZ0Z_0_cascade_ ;
    wire \POWERLED.count_off_0_0 ;
    wire \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ;
    wire \POWERLED.N_116 ;
    wire \POWERLED.count_off_0_4 ;
    wire \POWERLED.count_off_enZ0 ;
    wire v33s_ok;
    wire vccst_cpu_ok;
    wire slp_s3n_signal;
    wire rsmrst_pwrgd_signal;
    wire v5s_ok;
    wire \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ;
    wire dsw_pwrok;
    wire vccin_en;
    wire \VPP_VDDQ.delayed_vddq_okZ0_cascade_ ;
    wire pch_pwrok;
    wire vccst_pwrgd;
    wire \VPP_VDDQ.delayed_vddq_ok_en ;
    wire \VPP_VDDQ.delayed_vddq_ok_en_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_ok_0 ;
    wire \VPP_VDDQ.N_53 ;
    wire \VPP_VDDQ.N_53_i ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ;
    wire \POWERLED.count_clk_0_11 ;
    wire \POWERLED.count_clk_0_12 ;
    wire \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.func_state_RNICAC53_0_0 ;
    wire \POWERLED.count_clk_0_1 ;
    wire \POWERLED.count_clk_en ;
    wire \POWERLED.count_clk_RNIZ0Z_0 ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.N_163 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.count_clkZ0Z_1_cascade_ ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.N_176 ;
    wire \VPP_VDDQ.N_47_cascade_ ;
    wire \VPP_VDDQ.count_2_RNIZ0Z_1 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_2_1_1 ;
    wire \VPP_VDDQ.curr_state_2_0_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ;
    wire \VPP_VDDQ.count_2_1_2 ;
    wire \VPP_VDDQ.count_2_1_3_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_3 ;
    wire \VPP_VDDQ.N_385 ;
    wire \VPP_VDDQ.N_385_cascade_ ;
    wire \VPP_VDDQ.curr_state_2_0_0 ;
    wire \VPP_VDDQ.m4_0_cascade_ ;
    wire suswarn_n;
    wire \VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ;
    wire N_579_g;
    wire \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_6 ;
    wire \VPP_VDDQ.count_2_1_6 ;
    wire \VPP_VDDQ.curr_state_2_RNIZ0Z_1 ;
    wire vddq_ok;
    wire N_362;
    wire \VPP_VDDQ.count_2_1_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_9 ;
    wire \VPP_VDDQ.un9_clk_100khz_12 ;
    wire \VPP_VDDQ.un9_clk_100khz_4_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_11 ;
    wire \VPP_VDDQ.N_1_i_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0 ;
    wire \VPP_VDDQ.count_2_0_0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ;
    wire \VPP_VDDQ.count_2_1_7 ;
    wire \VPP_VDDQ.count_2Z0Z_7 ;
    wire \VPP_VDDQ.count_2_1_7_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_7 ;
    wire \VPP_VDDQ.count_2_1_12_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ;
    wire \VPP_VDDQ.count_2_0_14 ;
    wire \VPP_VDDQ.count_2_1_14_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ;
    wire \VPP_VDDQ.count_2_0_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7 ;
    wire \VPP_VDDQ.count_2_0_6 ;
    wire \VPP_VDDQ.count_2_0_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ;
    wire \VPP_VDDQ.count_2_1_8 ;
    wire \VPP_VDDQ.count_2_1_11_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_11 ;
    wire \VPP_VDDQ.count_2Z0Z_11_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ;
    wire \VPP_VDDQ.count_2_0_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ;
    wire \VPP_VDDQ.count_2_1_10 ;
    wire \VPP_VDDQ.count_2Z0Z_10 ;
    wire \VPP_VDDQ.count_2_1_10_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_10 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ;
    wire \VPP_VDDQ.N_1_i ;
    wire \VPP_VDDQ.count_2_0_12 ;
    wire fpga_osc;
    wire \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ;
    wire _gnd_net_;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__34245),
            .DIN(N__34244),
            .DOUT(N__34243),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__34245),
            .PADOUT(N__34244),
            .PADIN(N__34243),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__34236),
            .DIN(N__34235),
            .DOUT(N__34234),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__34236),
            .PADOUT(N__34235),
            .PADIN(N__34234),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15452),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__34227),
            .DIN(N__34226),
            .DOUT(N__34225),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__34227),
            .PADOUT(N__34226),
            .PADIN(N__34225),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16306),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__34218),
            .DIN(N__34217),
            .DOUT(N__34216),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__34218),
            .PADOUT(N__34217),
            .PADIN(N__34216),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15761),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__34209),
            .DIN(N__34208),
            .DOUT(N__34207),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__34209),
            .PADOUT(N__34208),
            .PADIN(N__34207),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__34200),
            .DIN(N__34199),
            .DOUT(N__34198),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__34200),
            .PADOUT(N__34199),
            .PADIN(N__34198),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__34191),
            .DIN(N__34190),
            .DOUT(N__34189),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__34191),
            .PADOUT(N__34190),
            .PADIN(N__34189),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__34182),
            .DIN(N__34181),
            .DOUT(N__34180),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__34182),
            .PADOUT(N__34181),
            .PADIN(N__34180),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__34173),
            .DIN(N__34172),
            .DOUT(N__34171),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__34173),
            .PADOUT(N__34172),
            .PADIN(N__34171),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16333),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__34164),
            .DIN(N__34163),
            .DOUT(N__34162),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__34164),
            .PADOUT(N__34163),
            .PADIN(N__34162),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__34155),
            .DIN(N__34154),
            .DOUT(N__34153),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__34155),
            .PADOUT(N__34154),
            .PADIN(N__34153),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__34146),
            .DIN(N__34145),
            .DOUT(N__34144),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__34146),
            .PADOUT(N__34145),
            .PADIN(N__34144),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17582),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__34137),
            .DIN(N__34136),
            .DOUT(N__34135),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__34137),
            .PADOUT(N__34136),
            .PADIN(N__34135),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__34128),
            .DIN(N__34127),
            .DOUT(N__34126),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__34128),
            .PADOUT(N__34127),
            .PADIN(N__34126),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__34119),
            .DIN(N__34118),
            .DOUT(N__34117),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__34119),
            .PADOUT(N__34118),
            .PADIN(N__34117),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__34110),
            .DIN(N__34109),
            .DOUT(N__34108),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__34110),
            .PADOUT(N__34109),
            .PADIN(N__34108),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__34101),
            .DIN(N__34100),
            .DOUT(N__34099),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__34101),
            .PADOUT(N__34100),
            .PADIN(N__34099),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29269),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__34092),
            .DIN(N__34091),
            .DOUT(N__34090),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__34092),
            .PADOUT(N__34091),
            .PADIN(N__34090),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33dsw_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__34083),
            .DIN(N__34082),
            .DOUT(N__34081),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__34083),
            .PADOUT(N__34082),
            .PADIN(N__34081),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__34074),
            .DIN(N__34073),
            .DOUT(N__34072),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__34074),
            .PADOUT(N__34073),
            .PADIN(N__34072),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31958),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__34065),
            .DIN(N__34064),
            .DOUT(N__34063),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__34065),
            .PADOUT(N__34064),
            .PADIN(N__34063),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__34056),
            .DIN(N__34055),
            .DOUT(N__34054),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__34056),
            .PADOUT(N__34055),
            .PADIN(N__34054),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__34047),
            .DIN(N__34046),
            .DOUT(N__34045),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__34047),
            .PADOUT(N__34046),
            .PADIN(N__34045),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__34038),
            .DIN(N__34037),
            .DOUT(N__34036),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__34038),
            .PADOUT(N__34037),
            .PADIN(N__34036),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__34029),
            .DIN(N__34028),
            .DOUT(N__34027),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__34029),
            .PADOUT(N__34028),
            .PADIN(N__34027),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22406),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__34020),
            .DIN(N__34019),
            .DOUT(N__34018),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__34020),
            .PADOUT(N__34019),
            .PADIN(N__34018),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__34011),
            .DIN(N__34010),
            .DOUT(N__34009),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__34011),
            .PADOUT(N__34010),
            .PADIN(N__34009),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30275),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__34002),
            .DIN(N__34001),
            .DOUT(N__34000),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__34002),
            .PADOUT(N__34001),
            .PADIN(N__34000),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30335),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__33993),
            .DIN(N__33992),
            .DOUT(N__33991),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__33993),
            .PADOUT(N__33992),
            .PADIN(N__33991),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__33984),
            .DIN(N__33983),
            .DOUT(N__33982),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__33984),
            .PADOUT(N__33983),
            .PADIN(N__33982),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__33975),
            .DIN(N__33974),
            .DOUT(N__33973),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__33975),
            .PADOUT(N__33974),
            .PADIN(N__33973),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__33966),
            .DIN(N__33965),
            .DOUT(N__33964),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__33966),
            .PADOUT(N__33965),
            .PADIN(N__33964),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__33957),
            .DIN(N__33956),
            .DOUT(N__33955),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__33957),
            .PADOUT(N__33956),
            .PADIN(N__33955),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27460),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__33948),
            .DIN(N__33947),
            .DOUT(N__33946),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__33948),
            .PADOUT(N__33947),
            .PADIN(N__33946),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20366),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__33939),
            .DIN(N__33938),
            .DOUT(N__33937),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__33939),
            .PADOUT(N__33938),
            .PADIN(N__33937),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__33930),
            .DIN(N__33929),
            .DOUT(N__33928),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__33930),
            .PADOUT(N__33929),
            .PADIN(N__33928),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29288),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__33921),
            .DIN(N__33920),
            .DOUT(N__33919),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__33921),
            .PADOUT(N__33920),
            .PADIN(N__33919),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__33912),
            .DIN(N__33911),
            .DOUT(N__33910),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__33912),
            .PADOUT(N__33911),
            .PADIN(N__33910),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__33903),
            .DIN(N__33902),
            .DOUT(N__33901),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__33903),
            .PADOUT(N__33902),
            .PADIN(N__33901),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__33894),
            .DIN(N__33893),
            .DOUT(N__33892),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__33894),
            .PADOUT(N__33893),
            .PADIN(N__33892),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__33885),
            .DIN(N__33884),
            .DOUT(N__33883),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__33885),
            .PADOUT(N__33884),
            .PADIN(N__33883),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16223),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__33876),
            .DIN(N__33875),
            .DOUT(N__33874),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__33876),
            .PADOUT(N__33875),
            .PADIN(N__33874),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__33867),
            .DIN(N__33866),
            .DOUT(N__33865),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__33867),
            .PADOUT(N__33866),
            .PADIN(N__33865),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16337),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__33858),
            .DIN(N__33857),
            .DOUT(N__33856),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__33858),
            .PADOUT(N__33857),
            .PADIN(N__33856),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__33849),
            .DIN(N__33848),
            .DOUT(N__33847),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__33849),
            .PADOUT(N__33848),
            .PADIN(N__33847),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30385),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__33840),
            .DIN(N__33839),
            .DOUT(N__33838),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__33840),
            .PADOUT(N__33839),
            .PADIN(N__33838),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16307),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__33831),
            .DIN(N__33830),
            .DOUT(N__33829),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__33831),
            .PADOUT(N__33830),
            .PADIN(N__33829),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__33822),
            .DIN(N__33821),
            .DOUT(N__33820),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__33822),
            .PADOUT(N__33821),
            .PADIN(N__33820),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__33813),
            .DIN(N__33812),
            .DOUT(N__33811),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__33813),
            .PADOUT(N__33812),
            .PADIN(N__33811),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__33804),
            .DIN(N__33803),
            .DOUT(N__33802),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__33804),
            .PADOUT(N__33803),
            .PADIN(N__33802),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__33795),
            .DIN(N__33794),
            .DOUT(N__33793),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__33795),
            .PADOUT(N__33794),
            .PADIN(N__33793),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30356),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__33786),
            .DIN(N__33785),
            .DOUT(N__33784),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__33786),
            .PADOUT(N__33785),
            .PADIN(N__33784),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__33777),
            .DIN(N__33776),
            .DOUT(N__33775),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__33777),
            .PADOUT(N__33776),
            .PADIN(N__33775),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__33768),
            .DIN(N__33767),
            .DOUT(N__33766),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__33768),
            .PADOUT(N__33767),
            .PADIN(N__33766),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__33759),
            .DIN(N__33758),
            .DOUT(N__33757),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__33759),
            .PADOUT(N__33758),
            .PADIN(N__33757),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__33750),
            .DIN(N__33749),
            .DOUT(N__33748),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__33750),
            .PADOUT(N__33749),
            .PADIN(N__33748),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__33741),
            .DIN(N__33740),
            .DOUT(N__33739),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__33741),
            .PADOUT(N__33740),
            .PADIN(N__33739),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__33732),
            .DIN(N__33731),
            .DOUT(N__33730),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__33732),
            .PADOUT(N__33731),
            .PADIN(N__33730),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30306),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__33723),
            .DIN(N__33722),
            .DOUT(N__33721),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__33723),
            .PADOUT(N__33722),
            .PADIN(N__33721),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    CascadeMux I__7867 (
            .O(N__33704),
            .I(N__33700));
    InMux I__7866 (
            .O(N__33703),
            .I(N__33695));
    InMux I__7865 (
            .O(N__33700),
            .I(N__33695));
    LocalMux I__7864 (
            .O(N__33695),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ));
    InMux I__7863 (
            .O(N__33692),
            .I(N__33689));
    LocalMux I__7862 (
            .O(N__33689),
            .I(\VPP_VDDQ.count_2_1_10 ));
    InMux I__7861 (
            .O(N__33686),
            .I(N__33682));
    InMux I__7860 (
            .O(N__33685),
            .I(N__33679));
    LocalMux I__7859 (
            .O(N__33682),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    LocalMux I__7858 (
            .O(N__33679),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    CascadeMux I__7857 (
            .O(N__33674),
            .I(\VPP_VDDQ.count_2_1_10_cascade_ ));
    InMux I__7856 (
            .O(N__33671),
            .I(N__33668));
    LocalMux I__7855 (
            .O(N__33668),
            .I(\VPP_VDDQ.un1_count_2_1_axb_10 ));
    CascadeMux I__7854 (
            .O(N__33665),
            .I(N__33651));
    CascadeMux I__7853 (
            .O(N__33664),
            .I(N__33648));
    CascadeMux I__7852 (
            .O(N__33663),
            .I(N__33644));
    CascadeMux I__7851 (
            .O(N__33662),
            .I(N__33641));
    InMux I__7850 (
            .O(N__33661),
            .I(N__33638));
    InMux I__7849 (
            .O(N__33660),
            .I(N__33635));
    CascadeMux I__7848 (
            .O(N__33659),
            .I(N__33627));
    CascadeMux I__7847 (
            .O(N__33658),
            .I(N__33622));
    CascadeMux I__7846 (
            .O(N__33657),
            .I(N__33612));
    InMux I__7845 (
            .O(N__33656),
            .I(N__33609));
    InMux I__7844 (
            .O(N__33655),
            .I(N__33598));
    InMux I__7843 (
            .O(N__33654),
            .I(N__33598));
    InMux I__7842 (
            .O(N__33651),
            .I(N__33598));
    InMux I__7841 (
            .O(N__33648),
            .I(N__33598));
    InMux I__7840 (
            .O(N__33647),
            .I(N__33598));
    InMux I__7839 (
            .O(N__33644),
            .I(N__33593));
    InMux I__7838 (
            .O(N__33641),
            .I(N__33593));
    LocalMux I__7837 (
            .O(N__33638),
            .I(N__33588));
    LocalMux I__7836 (
            .O(N__33635),
            .I(N__33588));
    InMux I__7835 (
            .O(N__33634),
            .I(N__33577));
    InMux I__7834 (
            .O(N__33633),
            .I(N__33577));
    InMux I__7833 (
            .O(N__33632),
            .I(N__33577));
    InMux I__7832 (
            .O(N__33631),
            .I(N__33577));
    InMux I__7831 (
            .O(N__33630),
            .I(N__33577));
    InMux I__7830 (
            .O(N__33627),
            .I(N__33568));
    InMux I__7829 (
            .O(N__33626),
            .I(N__33568));
    InMux I__7828 (
            .O(N__33625),
            .I(N__33568));
    InMux I__7827 (
            .O(N__33622),
            .I(N__33568));
    CascadeMux I__7826 (
            .O(N__33621),
            .I(N__33564));
    CascadeMux I__7825 (
            .O(N__33620),
            .I(N__33561));
    CascadeMux I__7824 (
            .O(N__33619),
            .I(N__33551));
    CascadeMux I__7823 (
            .O(N__33618),
            .I(N__33548));
    InMux I__7822 (
            .O(N__33617),
            .I(N__33538));
    InMux I__7821 (
            .O(N__33616),
            .I(N__33538));
    InMux I__7820 (
            .O(N__33615),
            .I(N__33538));
    InMux I__7819 (
            .O(N__33612),
            .I(N__33535));
    LocalMux I__7818 (
            .O(N__33609),
            .I(N__33522));
    LocalMux I__7817 (
            .O(N__33598),
            .I(N__33522));
    LocalMux I__7816 (
            .O(N__33593),
            .I(N__33522));
    Span4Mux_v I__7815 (
            .O(N__33588),
            .I(N__33522));
    LocalMux I__7814 (
            .O(N__33577),
            .I(N__33522));
    LocalMux I__7813 (
            .O(N__33568),
            .I(N__33522));
    InMux I__7812 (
            .O(N__33567),
            .I(N__33507));
    InMux I__7811 (
            .O(N__33564),
            .I(N__33507));
    InMux I__7810 (
            .O(N__33561),
            .I(N__33507));
    InMux I__7809 (
            .O(N__33560),
            .I(N__33507));
    InMux I__7808 (
            .O(N__33559),
            .I(N__33507));
    InMux I__7807 (
            .O(N__33558),
            .I(N__33507));
    InMux I__7806 (
            .O(N__33557),
            .I(N__33507));
    InMux I__7805 (
            .O(N__33556),
            .I(N__33502));
    InMux I__7804 (
            .O(N__33555),
            .I(N__33502));
    InMux I__7803 (
            .O(N__33554),
            .I(N__33495));
    InMux I__7802 (
            .O(N__33551),
            .I(N__33495));
    InMux I__7801 (
            .O(N__33548),
            .I(N__33495));
    InMux I__7800 (
            .O(N__33547),
            .I(N__33488));
    InMux I__7799 (
            .O(N__33546),
            .I(N__33488));
    InMux I__7798 (
            .O(N__33545),
            .I(N__33488));
    LocalMux I__7797 (
            .O(N__33538),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7796 (
            .O(N__33535),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__7795 (
            .O(N__33522),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7794 (
            .O(N__33507),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7793 (
            .O(N__33502),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7792 (
            .O(N__33495),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7791 (
            .O(N__33488),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    CascadeMux I__7790 (
            .O(N__33473),
            .I(N__33467));
    CascadeMux I__7789 (
            .O(N__33472),
            .I(N__33461));
    InMux I__7788 (
            .O(N__33471),
            .I(N__33447));
    InMux I__7787 (
            .O(N__33470),
            .I(N__33436));
    InMux I__7786 (
            .O(N__33467),
            .I(N__33436));
    InMux I__7785 (
            .O(N__33466),
            .I(N__33436));
    InMux I__7784 (
            .O(N__33465),
            .I(N__33436));
    InMux I__7783 (
            .O(N__33464),
            .I(N__33436));
    InMux I__7782 (
            .O(N__33461),
            .I(N__33419));
    InMux I__7781 (
            .O(N__33460),
            .I(N__33419));
    InMux I__7780 (
            .O(N__33459),
            .I(N__33419));
    InMux I__7779 (
            .O(N__33458),
            .I(N__33419));
    InMux I__7778 (
            .O(N__33457),
            .I(N__33406));
    InMux I__7777 (
            .O(N__33456),
            .I(N__33406));
    InMux I__7776 (
            .O(N__33455),
            .I(N__33406));
    InMux I__7775 (
            .O(N__33454),
            .I(N__33406));
    InMux I__7774 (
            .O(N__33453),
            .I(N__33406));
    InMux I__7773 (
            .O(N__33452),
            .I(N__33406));
    CascadeMux I__7772 (
            .O(N__33451),
            .I(N__33403));
    CascadeMux I__7771 (
            .O(N__33450),
            .I(N__33394));
    LocalMux I__7770 (
            .O(N__33447),
            .I(N__33386));
    LocalMux I__7769 (
            .O(N__33436),
            .I(N__33386));
    InMux I__7768 (
            .O(N__33435),
            .I(N__33377));
    InMux I__7767 (
            .O(N__33434),
            .I(N__33377));
    InMux I__7766 (
            .O(N__33433),
            .I(N__33377));
    InMux I__7765 (
            .O(N__33432),
            .I(N__33377));
    InMux I__7764 (
            .O(N__33431),
            .I(N__33374));
    InMux I__7763 (
            .O(N__33430),
            .I(N__33369));
    InMux I__7762 (
            .O(N__33429),
            .I(N__33369));
    InMux I__7761 (
            .O(N__33428),
            .I(N__33366));
    LocalMux I__7760 (
            .O(N__33419),
            .I(N__33361));
    LocalMux I__7759 (
            .O(N__33406),
            .I(N__33361));
    InMux I__7758 (
            .O(N__33403),
            .I(N__33346));
    InMux I__7757 (
            .O(N__33402),
            .I(N__33346));
    InMux I__7756 (
            .O(N__33401),
            .I(N__33346));
    InMux I__7755 (
            .O(N__33400),
            .I(N__33346));
    InMux I__7754 (
            .O(N__33399),
            .I(N__33346));
    InMux I__7753 (
            .O(N__33398),
            .I(N__33346));
    InMux I__7752 (
            .O(N__33397),
            .I(N__33346));
    InMux I__7751 (
            .O(N__33394),
            .I(N__33337));
    InMux I__7750 (
            .O(N__33393),
            .I(N__33337));
    InMux I__7749 (
            .O(N__33392),
            .I(N__33337));
    InMux I__7748 (
            .O(N__33391),
            .I(N__33337));
    Span4Mux_v I__7747 (
            .O(N__33386),
            .I(N__33332));
    LocalMux I__7746 (
            .O(N__33377),
            .I(N__33332));
    LocalMux I__7745 (
            .O(N__33374),
            .I(N__33329));
    LocalMux I__7744 (
            .O(N__33369),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7743 (
            .O(N__33366),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv12 I__7742 (
            .O(N__33361),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7741 (
            .O(N__33346),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7740 (
            .O(N__33337),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7739 (
            .O(N__33332),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7738 (
            .O(N__33329),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    CascadeMux I__7737 (
            .O(N__33314),
            .I(N__33310));
    InMux I__7736 (
            .O(N__33313),
            .I(N__33307));
    InMux I__7735 (
            .O(N__33310),
            .I(N__33304));
    LocalMux I__7734 (
            .O(N__33307),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ));
    LocalMux I__7733 (
            .O(N__33304),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ));
    CascadeMux I__7732 (
            .O(N__33299),
            .I(N__33294));
    CascadeMux I__7731 (
            .O(N__33298),
            .I(N__33287));
    CascadeMux I__7730 (
            .O(N__33297),
            .I(N__33274));
    InMux I__7729 (
            .O(N__33294),
            .I(N__33257));
    InMux I__7728 (
            .O(N__33293),
            .I(N__33257));
    InMux I__7727 (
            .O(N__33292),
            .I(N__33257));
    InMux I__7726 (
            .O(N__33291),
            .I(N__33257));
    InMux I__7725 (
            .O(N__33290),
            .I(N__33257));
    InMux I__7724 (
            .O(N__33287),
            .I(N__33254));
    InMux I__7723 (
            .O(N__33286),
            .I(N__33245));
    InMux I__7722 (
            .O(N__33285),
            .I(N__33245));
    InMux I__7721 (
            .O(N__33284),
            .I(N__33245));
    InMux I__7720 (
            .O(N__33283),
            .I(N__33245));
    InMux I__7719 (
            .O(N__33282),
            .I(N__33225));
    InMux I__7718 (
            .O(N__33281),
            .I(N__33225));
    InMux I__7717 (
            .O(N__33280),
            .I(N__33225));
    InMux I__7716 (
            .O(N__33279),
            .I(N__33225));
    InMux I__7715 (
            .O(N__33278),
            .I(N__33225));
    InMux I__7714 (
            .O(N__33277),
            .I(N__33220));
    InMux I__7713 (
            .O(N__33274),
            .I(N__33220));
    InMux I__7712 (
            .O(N__33273),
            .I(N__33209));
    InMux I__7711 (
            .O(N__33272),
            .I(N__33209));
    InMux I__7710 (
            .O(N__33271),
            .I(N__33209));
    InMux I__7709 (
            .O(N__33270),
            .I(N__33209));
    InMux I__7708 (
            .O(N__33269),
            .I(N__33209));
    InMux I__7707 (
            .O(N__33268),
            .I(N__33204));
    LocalMux I__7706 (
            .O(N__33257),
            .I(N__33197));
    LocalMux I__7705 (
            .O(N__33254),
            .I(N__33197));
    LocalMux I__7704 (
            .O(N__33245),
            .I(N__33197));
    InMux I__7703 (
            .O(N__33244),
            .I(N__33184));
    InMux I__7702 (
            .O(N__33243),
            .I(N__33184));
    InMux I__7701 (
            .O(N__33242),
            .I(N__33184));
    InMux I__7700 (
            .O(N__33241),
            .I(N__33184));
    InMux I__7699 (
            .O(N__33240),
            .I(N__33184));
    InMux I__7698 (
            .O(N__33239),
            .I(N__33184));
    InMux I__7697 (
            .O(N__33238),
            .I(N__33177));
    InMux I__7696 (
            .O(N__33237),
            .I(N__33177));
    InMux I__7695 (
            .O(N__33236),
            .I(N__33177));
    LocalMux I__7694 (
            .O(N__33225),
            .I(N__33170));
    LocalMux I__7693 (
            .O(N__33220),
            .I(N__33170));
    LocalMux I__7692 (
            .O(N__33209),
            .I(N__33170));
    InMux I__7691 (
            .O(N__33208),
            .I(N__33165));
    InMux I__7690 (
            .O(N__33207),
            .I(N__33165));
    LocalMux I__7689 (
            .O(N__33204),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7688 (
            .O(N__33197),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7687 (
            .O(N__33184),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7686 (
            .O(N__33177),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7685 (
            .O(N__33170),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7684 (
            .O(N__33165),
            .I(\VPP_VDDQ.N_1_i ));
    InMux I__7683 (
            .O(N__33152),
            .I(N__33149));
    LocalMux I__7682 (
            .O(N__33149),
            .I(\VPP_VDDQ.count_2_0_12 ));
    ClkMux I__7681 (
            .O(N__33146),
            .I(N__33143));
    LocalMux I__7680 (
            .O(N__33143),
            .I(N__33132));
    ClkMux I__7679 (
            .O(N__33142),
            .I(N__33129));
    ClkMux I__7678 (
            .O(N__33141),
            .I(N__33124));
    ClkMux I__7677 (
            .O(N__33140),
            .I(N__33120));
    ClkMux I__7676 (
            .O(N__33139),
            .I(N__33117));
    ClkMux I__7675 (
            .O(N__33138),
            .I(N__33114));
    ClkMux I__7674 (
            .O(N__33137),
            .I(N__33107));
    ClkMux I__7673 (
            .O(N__33136),
            .I(N__33104));
    ClkMux I__7672 (
            .O(N__33135),
            .I(N__33101));
    Span4Mux_s2_h I__7671 (
            .O(N__33132),
            .I(N__33094));
    LocalMux I__7670 (
            .O(N__33129),
            .I(N__33094));
    ClkMux I__7669 (
            .O(N__33128),
            .I(N__33091));
    ClkMux I__7668 (
            .O(N__33127),
            .I(N__33087));
    LocalMux I__7667 (
            .O(N__33124),
            .I(N__33082));
    ClkMux I__7666 (
            .O(N__33123),
            .I(N__33079));
    LocalMux I__7665 (
            .O(N__33120),
            .I(N__33072));
    LocalMux I__7664 (
            .O(N__33117),
            .I(N__33072));
    LocalMux I__7663 (
            .O(N__33114),
            .I(N__33063));
    ClkMux I__7662 (
            .O(N__33113),
            .I(N__33060));
    ClkMux I__7661 (
            .O(N__33112),
            .I(N__33056));
    ClkMux I__7660 (
            .O(N__33111),
            .I(N__33053));
    ClkMux I__7659 (
            .O(N__33110),
            .I(N__33045));
    LocalMux I__7658 (
            .O(N__33107),
            .I(N__33042));
    LocalMux I__7657 (
            .O(N__33104),
            .I(N__33039));
    LocalMux I__7656 (
            .O(N__33101),
            .I(N__33036));
    ClkMux I__7655 (
            .O(N__33100),
            .I(N__33033));
    ClkMux I__7654 (
            .O(N__33099),
            .I(N__33030));
    Span4Mux_v I__7653 (
            .O(N__33094),
            .I(N__33023));
    LocalMux I__7652 (
            .O(N__33091),
            .I(N__33023));
    ClkMux I__7651 (
            .O(N__33090),
            .I(N__33020));
    LocalMux I__7650 (
            .O(N__33087),
            .I(N__33017));
    ClkMux I__7649 (
            .O(N__33086),
            .I(N__33013));
    ClkMux I__7648 (
            .O(N__33085),
            .I(N__33010));
    Span4Mux_s2_h I__7647 (
            .O(N__33082),
            .I(N__33005));
    LocalMux I__7646 (
            .O(N__33079),
            .I(N__33005));
    ClkMux I__7645 (
            .O(N__33078),
            .I(N__33002));
    ClkMux I__7644 (
            .O(N__33077),
            .I(N__32999));
    Span4Mux_h I__7643 (
            .O(N__33072),
            .I(N__32996));
    ClkMux I__7642 (
            .O(N__33071),
            .I(N__32993));
    ClkMux I__7641 (
            .O(N__33070),
            .I(N__32990));
    ClkMux I__7640 (
            .O(N__33069),
            .I(N__32986));
    ClkMux I__7639 (
            .O(N__33068),
            .I(N__32982));
    ClkMux I__7638 (
            .O(N__33067),
            .I(N__32978));
    ClkMux I__7637 (
            .O(N__33066),
            .I(N__32975));
    Span4Mux_v I__7636 (
            .O(N__33063),
            .I(N__32968));
    LocalMux I__7635 (
            .O(N__33060),
            .I(N__32965));
    ClkMux I__7634 (
            .O(N__33059),
            .I(N__32960));
    LocalMux I__7633 (
            .O(N__33056),
            .I(N__32956));
    LocalMux I__7632 (
            .O(N__33053),
            .I(N__32953));
    ClkMux I__7631 (
            .O(N__33052),
            .I(N__32950));
    ClkMux I__7630 (
            .O(N__33051),
            .I(N__32945));
    ClkMux I__7629 (
            .O(N__33050),
            .I(N__32939));
    ClkMux I__7628 (
            .O(N__33049),
            .I(N__32936));
    ClkMux I__7627 (
            .O(N__33048),
            .I(N__32932));
    LocalMux I__7626 (
            .O(N__33045),
            .I(N__32929));
    Span4Mux_v I__7625 (
            .O(N__33042),
            .I(N__32918));
    Span4Mux_v I__7624 (
            .O(N__33039),
            .I(N__32918));
    Span4Mux_s1_h I__7623 (
            .O(N__33036),
            .I(N__32918));
    LocalMux I__7622 (
            .O(N__33033),
            .I(N__32918));
    LocalMux I__7621 (
            .O(N__33030),
            .I(N__32915));
    ClkMux I__7620 (
            .O(N__33029),
            .I(N__32912));
    ClkMux I__7619 (
            .O(N__33028),
            .I(N__32908));
    Span4Mux_h I__7618 (
            .O(N__33023),
            .I(N__32901));
    LocalMux I__7617 (
            .O(N__33020),
            .I(N__32901));
    Span4Mux_s2_h I__7616 (
            .O(N__33017),
            .I(N__32896));
    ClkMux I__7615 (
            .O(N__33016),
            .I(N__32893));
    LocalMux I__7614 (
            .O(N__33013),
            .I(N__32888));
    LocalMux I__7613 (
            .O(N__33010),
            .I(N__32888));
    Span4Mux_h I__7612 (
            .O(N__33005),
            .I(N__32884));
    LocalMux I__7611 (
            .O(N__33002),
            .I(N__32879));
    LocalMux I__7610 (
            .O(N__32999),
            .I(N__32879));
    Span4Mux_v I__7609 (
            .O(N__32996),
            .I(N__32872));
    LocalMux I__7608 (
            .O(N__32993),
            .I(N__32872));
    LocalMux I__7607 (
            .O(N__32990),
            .I(N__32872));
    ClkMux I__7606 (
            .O(N__32989),
            .I(N__32869));
    LocalMux I__7605 (
            .O(N__32986),
            .I(N__32866));
    ClkMux I__7604 (
            .O(N__32985),
            .I(N__32863));
    LocalMux I__7603 (
            .O(N__32982),
            .I(N__32860));
    ClkMux I__7602 (
            .O(N__32981),
            .I(N__32857));
    LocalMux I__7601 (
            .O(N__32978),
            .I(N__32854));
    LocalMux I__7600 (
            .O(N__32975),
            .I(N__32851));
    ClkMux I__7599 (
            .O(N__32974),
            .I(N__32848));
    ClkMux I__7598 (
            .O(N__32973),
            .I(N__32845));
    ClkMux I__7597 (
            .O(N__32972),
            .I(N__32840));
    ClkMux I__7596 (
            .O(N__32971),
            .I(N__32837));
    Span4Mux_h I__7595 (
            .O(N__32968),
            .I(N__32832));
    Span4Mux_v I__7594 (
            .O(N__32965),
            .I(N__32832));
    ClkMux I__7593 (
            .O(N__32964),
            .I(N__32829));
    ClkMux I__7592 (
            .O(N__32963),
            .I(N__32826));
    LocalMux I__7591 (
            .O(N__32960),
            .I(N__32823));
    ClkMux I__7590 (
            .O(N__32959),
            .I(N__32820));
    Span4Mux_v I__7589 (
            .O(N__32956),
            .I(N__32814));
    Span4Mux_s1_h I__7588 (
            .O(N__32953),
            .I(N__32814));
    LocalMux I__7587 (
            .O(N__32950),
            .I(N__32811));
    ClkMux I__7586 (
            .O(N__32949),
            .I(N__32808));
    ClkMux I__7585 (
            .O(N__32948),
            .I(N__32805));
    LocalMux I__7584 (
            .O(N__32945),
            .I(N__32802));
    ClkMux I__7583 (
            .O(N__32944),
            .I(N__32799));
    ClkMux I__7582 (
            .O(N__32943),
            .I(N__32795));
    ClkMux I__7581 (
            .O(N__32942),
            .I(N__32791));
    LocalMux I__7580 (
            .O(N__32939),
            .I(N__32788));
    LocalMux I__7579 (
            .O(N__32936),
            .I(N__32785));
    ClkMux I__7578 (
            .O(N__32935),
            .I(N__32782));
    LocalMux I__7577 (
            .O(N__32932),
            .I(N__32777));
    Span4Mux_h I__7576 (
            .O(N__32929),
            .I(N__32777));
    ClkMux I__7575 (
            .O(N__32928),
            .I(N__32773));
    ClkMux I__7574 (
            .O(N__32927),
            .I(N__32770));
    Span4Mux_v I__7573 (
            .O(N__32918),
            .I(N__32764));
    Span4Mux_h I__7572 (
            .O(N__32915),
            .I(N__32764));
    LocalMux I__7571 (
            .O(N__32912),
            .I(N__32761));
    ClkMux I__7570 (
            .O(N__32911),
            .I(N__32758));
    LocalMux I__7569 (
            .O(N__32908),
            .I(N__32755));
    ClkMux I__7568 (
            .O(N__32907),
            .I(N__32752));
    ClkMux I__7567 (
            .O(N__32906),
            .I(N__32749));
    Span4Mux_v I__7566 (
            .O(N__32901),
            .I(N__32744));
    ClkMux I__7565 (
            .O(N__32900),
            .I(N__32741));
    ClkMux I__7564 (
            .O(N__32899),
            .I(N__32738));
    Span4Mux_h I__7563 (
            .O(N__32896),
            .I(N__32731));
    LocalMux I__7562 (
            .O(N__32893),
            .I(N__32731));
    Span4Mux_h I__7561 (
            .O(N__32888),
            .I(N__32731));
    ClkMux I__7560 (
            .O(N__32887),
            .I(N__32728));
    Span4Mux_v I__7559 (
            .O(N__32884),
            .I(N__32719));
    Span4Mux_v I__7558 (
            .O(N__32879),
            .I(N__32719));
    Span4Mux_v I__7557 (
            .O(N__32872),
            .I(N__32719));
    LocalMux I__7556 (
            .O(N__32869),
            .I(N__32719));
    Span4Mux_v I__7555 (
            .O(N__32866),
            .I(N__32714));
    LocalMux I__7554 (
            .O(N__32863),
            .I(N__32714));
    Span4Mux_s2_h I__7553 (
            .O(N__32860),
            .I(N__32709));
    LocalMux I__7552 (
            .O(N__32857),
            .I(N__32709));
    Span4Mux_v I__7551 (
            .O(N__32854),
            .I(N__32700));
    Span4Mux_v I__7550 (
            .O(N__32851),
            .I(N__32700));
    LocalMux I__7549 (
            .O(N__32848),
            .I(N__32700));
    LocalMux I__7548 (
            .O(N__32845),
            .I(N__32700));
    ClkMux I__7547 (
            .O(N__32844),
            .I(N__32697));
    ClkMux I__7546 (
            .O(N__32843),
            .I(N__32694));
    LocalMux I__7545 (
            .O(N__32840),
            .I(N__32690));
    LocalMux I__7544 (
            .O(N__32837),
            .I(N__32687));
    Span4Mux_v I__7543 (
            .O(N__32832),
            .I(N__32680));
    LocalMux I__7542 (
            .O(N__32829),
            .I(N__32680));
    LocalMux I__7541 (
            .O(N__32826),
            .I(N__32677));
    Span4Mux_v I__7540 (
            .O(N__32823),
            .I(N__32672));
    LocalMux I__7539 (
            .O(N__32820),
            .I(N__32672));
    ClkMux I__7538 (
            .O(N__32819),
            .I(N__32669));
    Span4Mux_h I__7537 (
            .O(N__32814),
            .I(N__32660));
    Span4Mux_v I__7536 (
            .O(N__32811),
            .I(N__32660));
    LocalMux I__7535 (
            .O(N__32808),
            .I(N__32660));
    LocalMux I__7534 (
            .O(N__32805),
            .I(N__32660));
    Span4Mux_s1_h I__7533 (
            .O(N__32802),
            .I(N__32655));
    LocalMux I__7532 (
            .O(N__32799),
            .I(N__32655));
    ClkMux I__7531 (
            .O(N__32798),
            .I(N__32652));
    LocalMux I__7530 (
            .O(N__32795),
            .I(N__32649));
    ClkMux I__7529 (
            .O(N__32794),
            .I(N__32646));
    LocalMux I__7528 (
            .O(N__32791),
            .I(N__32643));
    Span4Mux_v I__7527 (
            .O(N__32788),
            .I(N__32640));
    Span4Mux_s1_h I__7526 (
            .O(N__32785),
            .I(N__32635));
    LocalMux I__7525 (
            .O(N__32782),
            .I(N__32635));
    Span4Mux_v I__7524 (
            .O(N__32777),
            .I(N__32631));
    ClkMux I__7523 (
            .O(N__32776),
            .I(N__32628));
    LocalMux I__7522 (
            .O(N__32773),
            .I(N__32625));
    LocalMux I__7521 (
            .O(N__32770),
            .I(N__32622));
    ClkMux I__7520 (
            .O(N__32769),
            .I(N__32619));
    Span4Mux_v I__7519 (
            .O(N__32764),
            .I(N__32612));
    Span4Mux_v I__7518 (
            .O(N__32761),
            .I(N__32612));
    LocalMux I__7517 (
            .O(N__32758),
            .I(N__32612));
    Span4Mux_s1_h I__7516 (
            .O(N__32755),
            .I(N__32605));
    LocalMux I__7515 (
            .O(N__32752),
            .I(N__32605));
    LocalMux I__7514 (
            .O(N__32749),
            .I(N__32605));
    ClkMux I__7513 (
            .O(N__32748),
            .I(N__32602));
    ClkMux I__7512 (
            .O(N__32747),
            .I(N__32599));
    Span4Mux_v I__7511 (
            .O(N__32744),
            .I(N__32592));
    LocalMux I__7510 (
            .O(N__32741),
            .I(N__32592));
    LocalMux I__7509 (
            .O(N__32738),
            .I(N__32592));
    Span4Mux_v I__7508 (
            .O(N__32731),
            .I(N__32587));
    LocalMux I__7507 (
            .O(N__32728),
            .I(N__32587));
    Span4Mux_v I__7506 (
            .O(N__32719),
            .I(N__32580));
    Span4Mux_h I__7505 (
            .O(N__32714),
            .I(N__32580));
    Span4Mux_h I__7504 (
            .O(N__32709),
            .I(N__32580));
    Span4Mux_v I__7503 (
            .O(N__32700),
            .I(N__32573));
    LocalMux I__7502 (
            .O(N__32697),
            .I(N__32573));
    LocalMux I__7501 (
            .O(N__32694),
            .I(N__32573));
    ClkMux I__7500 (
            .O(N__32693),
            .I(N__32570));
    Span4Mux_h I__7499 (
            .O(N__32690),
            .I(N__32564));
    Span4Mux_h I__7498 (
            .O(N__32687),
            .I(N__32564));
    ClkMux I__7497 (
            .O(N__32686),
            .I(N__32561));
    ClkMux I__7496 (
            .O(N__32685),
            .I(N__32558));
    Span4Mux_v I__7495 (
            .O(N__32680),
            .I(N__32555));
    Span4Mux_v I__7494 (
            .O(N__32677),
            .I(N__32548));
    Span4Mux_s2_h I__7493 (
            .O(N__32672),
            .I(N__32548));
    LocalMux I__7492 (
            .O(N__32669),
            .I(N__32548));
    Span4Mux_v I__7491 (
            .O(N__32660),
            .I(N__32541));
    Span4Mux_h I__7490 (
            .O(N__32655),
            .I(N__32541));
    LocalMux I__7489 (
            .O(N__32652),
            .I(N__32541));
    Span4Mux_h I__7488 (
            .O(N__32649),
            .I(N__32534));
    LocalMux I__7487 (
            .O(N__32646),
            .I(N__32534));
    Span4Mux_h I__7486 (
            .O(N__32643),
            .I(N__32534));
    Span4Mux_v I__7485 (
            .O(N__32640),
            .I(N__32529));
    Span4Mux_h I__7484 (
            .O(N__32635),
            .I(N__32529));
    ClkMux I__7483 (
            .O(N__32634),
            .I(N__32526));
    Span4Mux_h I__7482 (
            .O(N__32631),
            .I(N__32521));
    LocalMux I__7481 (
            .O(N__32628),
            .I(N__32521));
    Span4Mux_s2_h I__7480 (
            .O(N__32625),
            .I(N__32512));
    Span4Mux_s2_h I__7479 (
            .O(N__32622),
            .I(N__32512));
    LocalMux I__7478 (
            .O(N__32619),
            .I(N__32512));
    Span4Mux_h I__7477 (
            .O(N__32612),
            .I(N__32512));
    Span4Mux_v I__7476 (
            .O(N__32605),
            .I(N__32507));
    LocalMux I__7475 (
            .O(N__32602),
            .I(N__32507));
    LocalMux I__7474 (
            .O(N__32599),
            .I(N__32504));
    Span4Mux_v I__7473 (
            .O(N__32592),
            .I(N__32493));
    Span4Mux_v I__7472 (
            .O(N__32587),
            .I(N__32493));
    IoSpan4Mux I__7471 (
            .O(N__32580),
            .I(N__32493));
    Span4Mux_h I__7470 (
            .O(N__32573),
            .I(N__32493));
    LocalMux I__7469 (
            .O(N__32570),
            .I(N__32493));
    ClkMux I__7468 (
            .O(N__32569),
            .I(N__32490));
    Span4Mux_v I__7467 (
            .O(N__32564),
            .I(N__32482));
    LocalMux I__7466 (
            .O(N__32561),
            .I(N__32482));
    LocalMux I__7465 (
            .O(N__32558),
            .I(N__32482));
    IoSpan4Mux I__7464 (
            .O(N__32555),
            .I(N__32479));
    Span4Mux_h I__7463 (
            .O(N__32548),
            .I(N__32472));
    Span4Mux_v I__7462 (
            .O(N__32541),
            .I(N__32472));
    Span4Mux_v I__7461 (
            .O(N__32534),
            .I(N__32472));
    Span4Mux_v I__7460 (
            .O(N__32529),
            .I(N__32467));
    LocalMux I__7459 (
            .O(N__32526),
            .I(N__32467));
    Span4Mux_v I__7458 (
            .O(N__32521),
            .I(N__32460));
    Span4Mux_h I__7457 (
            .O(N__32512),
            .I(N__32460));
    Span4Mux_h I__7456 (
            .O(N__32507),
            .I(N__32460));
    IoSpan4Mux I__7455 (
            .O(N__32504),
            .I(N__32455));
    IoSpan4Mux I__7454 (
            .O(N__32493),
            .I(N__32455));
    LocalMux I__7453 (
            .O(N__32490),
            .I(N__32452));
    ClkMux I__7452 (
            .O(N__32489),
            .I(N__32449));
    Span4Mux_v I__7451 (
            .O(N__32482),
            .I(N__32446));
    Odrv4 I__7450 (
            .O(N__32479),
            .I(fpga_osc));
    Odrv4 I__7449 (
            .O(N__32472),
            .I(fpga_osc));
    Odrv4 I__7448 (
            .O(N__32467),
            .I(fpga_osc));
    Odrv4 I__7447 (
            .O(N__32460),
            .I(fpga_osc));
    Odrv4 I__7446 (
            .O(N__32455),
            .I(fpga_osc));
    Odrv4 I__7445 (
            .O(N__32452),
            .I(fpga_osc));
    LocalMux I__7444 (
            .O(N__32449),
            .I(fpga_osc));
    Odrv4 I__7443 (
            .O(N__32446),
            .I(fpga_osc));
    CEMux I__7442 (
            .O(N__32429),
            .I(N__32426));
    LocalMux I__7441 (
            .O(N__32426),
            .I(N__32422));
    CEMux I__7440 (
            .O(N__32425),
            .I(N__32419));
    Span4Mux_v I__7439 (
            .O(N__32422),
            .I(N__32413));
    LocalMux I__7438 (
            .O(N__32419),
            .I(N__32413));
    CEMux I__7437 (
            .O(N__32418),
            .I(N__32410));
    Span4Mux_v I__7436 (
            .O(N__32413),
            .I(N__32404));
    LocalMux I__7435 (
            .O(N__32410),
            .I(N__32404));
    CEMux I__7434 (
            .O(N__32409),
            .I(N__32397));
    Span4Mux_h I__7433 (
            .O(N__32404),
            .I(N__32394));
    CEMux I__7432 (
            .O(N__32403),
            .I(N__32391));
    InMux I__7431 (
            .O(N__32402),
            .I(N__32388));
    InMux I__7430 (
            .O(N__32401),
            .I(N__32383));
    InMux I__7429 (
            .O(N__32400),
            .I(N__32383));
    LocalMux I__7428 (
            .O(N__32397),
            .I(N__32369));
    Span4Mux_s0_h I__7427 (
            .O(N__32394),
            .I(N__32369));
    LocalMux I__7426 (
            .O(N__32391),
            .I(N__32369));
    LocalMux I__7425 (
            .O(N__32388),
            .I(N__32364));
    LocalMux I__7424 (
            .O(N__32383),
            .I(N__32364));
    InMux I__7423 (
            .O(N__32382),
            .I(N__32351));
    InMux I__7422 (
            .O(N__32381),
            .I(N__32351));
    InMux I__7421 (
            .O(N__32380),
            .I(N__32346));
    InMux I__7420 (
            .O(N__32379),
            .I(N__32346));
    InMux I__7419 (
            .O(N__32378),
            .I(N__32339));
    InMux I__7418 (
            .O(N__32377),
            .I(N__32339));
    InMux I__7417 (
            .O(N__32376),
            .I(N__32339));
    Span4Mux_v I__7416 (
            .O(N__32369),
            .I(N__32334));
    Span4Mux_h I__7415 (
            .O(N__32364),
            .I(N__32334));
    InMux I__7414 (
            .O(N__32363),
            .I(N__32328));
    InMux I__7413 (
            .O(N__32362),
            .I(N__32325));
    InMux I__7412 (
            .O(N__32361),
            .I(N__32312));
    InMux I__7411 (
            .O(N__32360),
            .I(N__32312));
    InMux I__7410 (
            .O(N__32359),
            .I(N__32312));
    InMux I__7409 (
            .O(N__32358),
            .I(N__32312));
    InMux I__7408 (
            .O(N__32357),
            .I(N__32312));
    InMux I__7407 (
            .O(N__32356),
            .I(N__32312));
    LocalMux I__7406 (
            .O(N__32351),
            .I(N__32303));
    LocalMux I__7405 (
            .O(N__32346),
            .I(N__32303));
    LocalMux I__7404 (
            .O(N__32339),
            .I(N__32303));
    Span4Mux_v I__7403 (
            .O(N__32334),
            .I(N__32303));
    InMux I__7402 (
            .O(N__32333),
            .I(N__32296));
    InMux I__7401 (
            .O(N__32332),
            .I(N__32296));
    InMux I__7400 (
            .O(N__32331),
            .I(N__32296));
    LocalMux I__7399 (
            .O(N__32328),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    LocalMux I__7398 (
            .O(N__32325),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    LocalMux I__7397 (
            .O(N__32312),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    Odrv4 I__7396 (
            .O(N__32303),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    LocalMux I__7395 (
            .O(N__32296),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    CascadeMux I__7394 (
            .O(N__32285),
            .I(N__32282));
    InMux I__7393 (
            .O(N__32282),
            .I(N__32278));
    InMux I__7392 (
            .O(N__32281),
            .I(N__32275));
    LocalMux I__7391 (
            .O(N__32278),
            .I(N__32272));
    LocalMux I__7390 (
            .O(N__32275),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    Odrv4 I__7389 (
            .O(N__32272),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    InMux I__7388 (
            .O(N__32267),
            .I(N__32264));
    LocalMux I__7387 (
            .O(N__32264),
            .I(N__32261));
    Odrv12 I__7386 (
            .O(N__32261),
            .I(\VPP_VDDQ.count_2_0_3 ));
    CascadeMux I__7385 (
            .O(N__32258),
            .I(N__32255));
    InMux I__7384 (
            .O(N__32255),
            .I(N__32251));
    InMux I__7383 (
            .O(N__32254),
            .I(N__32248));
    LocalMux I__7382 (
            .O(N__32251),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7 ));
    LocalMux I__7381 (
            .O(N__32248),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7 ));
    InMux I__7380 (
            .O(N__32243),
            .I(N__32240));
    LocalMux I__7379 (
            .O(N__32240),
            .I(N__32237));
    Odrv4 I__7378 (
            .O(N__32237),
            .I(\VPP_VDDQ.count_2_0_6 ));
    InMux I__7377 (
            .O(N__32234),
            .I(N__32231));
    LocalMux I__7376 (
            .O(N__32231),
            .I(N__32228));
    Span4Mux_h I__7375 (
            .O(N__32228),
            .I(N__32225));
    Span4Mux_v I__7374 (
            .O(N__32225),
            .I(N__32222));
    Odrv4 I__7373 (
            .O(N__32222),
            .I(\VPP_VDDQ.count_2_0_8 ));
    CascadeMux I__7372 (
            .O(N__32219),
            .I(N__32215));
    InMux I__7371 (
            .O(N__32218),
            .I(N__32210));
    InMux I__7370 (
            .O(N__32215),
            .I(N__32210));
    LocalMux I__7369 (
            .O(N__32210),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ));
    InMux I__7368 (
            .O(N__32207),
            .I(N__32204));
    LocalMux I__7367 (
            .O(N__32204),
            .I(N__32201));
    Span12Mux_s11_v I__7366 (
            .O(N__32201),
            .I(N__32198));
    Odrv12 I__7365 (
            .O(N__32198),
            .I(\VPP_VDDQ.count_2_1_8 ));
    CascadeMux I__7364 (
            .O(N__32195),
            .I(\VPP_VDDQ.count_2_1_11_cascade_ ));
    InMux I__7363 (
            .O(N__32192),
            .I(N__32189));
    LocalMux I__7362 (
            .O(N__32189),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    CascadeMux I__7361 (
            .O(N__32186),
            .I(\VPP_VDDQ.count_2Z0Z_11_cascade_ ));
    InMux I__7360 (
            .O(N__32183),
            .I(N__32180));
    LocalMux I__7359 (
            .O(N__32180),
            .I(N__32177));
    Odrv12 I__7358 (
            .O(N__32177),
            .I(\VPP_VDDQ.un9_clk_100khz_5 ));
    CascadeMux I__7357 (
            .O(N__32174),
            .I(N__32170));
    InMux I__7356 (
            .O(N__32173),
            .I(N__32165));
    InMux I__7355 (
            .O(N__32170),
            .I(N__32165));
    LocalMux I__7354 (
            .O(N__32165),
            .I(N__32162));
    Odrv4 I__7353 (
            .O(N__32162),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ));
    InMux I__7352 (
            .O(N__32159),
            .I(N__32156));
    LocalMux I__7351 (
            .O(N__32156),
            .I(\VPP_VDDQ.count_2_0_11 ));
    CascadeMux I__7350 (
            .O(N__32153),
            .I(\VPP_VDDQ.N_1_i_cascade_ ));
    InMux I__7349 (
            .O(N__32150),
            .I(N__32146));
    InMux I__7348 (
            .O(N__32149),
            .I(N__32143));
    LocalMux I__7347 (
            .O(N__32146),
            .I(N__32138));
    LocalMux I__7346 (
            .O(N__32143),
            .I(N__32138));
    Span4Mux_h I__7345 (
            .O(N__32138),
            .I(N__32132));
    InMux I__7344 (
            .O(N__32137),
            .I(N__32127));
    InMux I__7343 (
            .O(N__32136),
            .I(N__32127));
    InMux I__7342 (
            .O(N__32135),
            .I(N__32124));
    Span4Mux_v I__7341 (
            .O(N__32132),
            .I(N__32121));
    LocalMux I__7340 (
            .O(N__32127),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__7339 (
            .O(N__32124),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    Odrv4 I__7338 (
            .O(N__32121),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    InMux I__7337 (
            .O(N__32114),
            .I(N__32111));
    LocalMux I__7336 (
            .O(N__32111),
            .I(\VPP_VDDQ.count_2_0_0 ));
    CascadeMux I__7335 (
            .O(N__32108),
            .I(N__32105));
    InMux I__7334 (
            .O(N__32105),
            .I(N__32099));
    InMux I__7333 (
            .O(N__32104),
            .I(N__32099));
    LocalMux I__7332 (
            .O(N__32099),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ));
    InMux I__7331 (
            .O(N__32096),
            .I(N__32093));
    LocalMux I__7330 (
            .O(N__32093),
            .I(\VPP_VDDQ.count_2_1_7 ));
    CascadeMux I__7329 (
            .O(N__32090),
            .I(N__32087));
    InMux I__7328 (
            .O(N__32087),
            .I(N__32081));
    InMux I__7327 (
            .O(N__32086),
            .I(N__32081));
    LocalMux I__7326 (
            .O(N__32081),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    CascadeMux I__7325 (
            .O(N__32078),
            .I(\VPP_VDDQ.count_2_1_7_cascade_ ));
    InMux I__7324 (
            .O(N__32075),
            .I(N__32072));
    LocalMux I__7323 (
            .O(N__32072),
            .I(\VPP_VDDQ.un1_count_2_1_axb_7 ));
    CascadeMux I__7322 (
            .O(N__32069),
            .I(\VPP_VDDQ.count_2_1_12_cascade_ ));
    InMux I__7321 (
            .O(N__32066),
            .I(N__32060));
    InMux I__7320 (
            .O(N__32065),
            .I(N__32060));
    LocalMux I__7319 (
            .O(N__32060),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    CascadeMux I__7318 (
            .O(N__32057),
            .I(N__32053));
    CascadeMux I__7317 (
            .O(N__32056),
            .I(N__32050));
    InMux I__7316 (
            .O(N__32053),
            .I(N__32047));
    InMux I__7315 (
            .O(N__32050),
            .I(N__32044));
    LocalMux I__7314 (
            .O(N__32047),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    LocalMux I__7313 (
            .O(N__32044),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    InMux I__7312 (
            .O(N__32039),
            .I(N__32036));
    LocalMux I__7311 (
            .O(N__32036),
            .I(\VPP_VDDQ.count_2_0_14 ));
    CascadeMux I__7310 (
            .O(N__32033),
            .I(\VPP_VDDQ.count_2_1_14_cascade_ ));
    InMux I__7309 (
            .O(N__32030),
            .I(N__32026));
    InMux I__7308 (
            .O(N__32029),
            .I(N__32023));
    LocalMux I__7307 (
            .O(N__32026),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    LocalMux I__7306 (
            .O(N__32023),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    InMux I__7305 (
            .O(N__32018),
            .I(N__32015));
    LocalMux I__7304 (
            .O(N__32015),
            .I(\VPP_VDDQ.curr_state_2_0_0 ));
    CascadeMux I__7303 (
            .O(N__32012),
            .I(\VPP_VDDQ.m4_0_cascade_ ));
    InMux I__7302 (
            .O(N__32009),
            .I(N__32005));
    InMux I__7301 (
            .O(N__32008),
            .I(N__31982));
    LocalMux I__7300 (
            .O(N__32005),
            .I(N__31979));
    InMux I__7299 (
            .O(N__32004),
            .I(N__31976));
    InMux I__7298 (
            .O(N__32003),
            .I(N__31973));
    InMux I__7297 (
            .O(N__32002),
            .I(N__31970));
    InMux I__7296 (
            .O(N__32001),
            .I(N__31964));
    InMux I__7295 (
            .O(N__32000),
            .I(N__31961));
    InMux I__7294 (
            .O(N__31999),
            .I(N__31955));
    InMux I__7293 (
            .O(N__31998),
            .I(N__31952));
    InMux I__7292 (
            .O(N__31997),
            .I(N__31943));
    InMux I__7291 (
            .O(N__31996),
            .I(N__31943));
    InMux I__7290 (
            .O(N__31995),
            .I(N__31943));
    InMux I__7289 (
            .O(N__31994),
            .I(N__31943));
    InMux I__7288 (
            .O(N__31993),
            .I(N__31938));
    InMux I__7287 (
            .O(N__31992),
            .I(N__31938));
    InMux I__7286 (
            .O(N__31991),
            .I(N__31931));
    InMux I__7285 (
            .O(N__31990),
            .I(N__31931));
    InMux I__7284 (
            .O(N__31989),
            .I(N__31931));
    InMux I__7283 (
            .O(N__31988),
            .I(N__31928));
    InMux I__7282 (
            .O(N__31987),
            .I(N__31921));
    InMux I__7281 (
            .O(N__31986),
            .I(N__31921));
    InMux I__7280 (
            .O(N__31985),
            .I(N__31921));
    LocalMux I__7279 (
            .O(N__31982),
            .I(N__31916));
    Span4Mux_s1_h I__7278 (
            .O(N__31979),
            .I(N__31916));
    LocalMux I__7277 (
            .O(N__31976),
            .I(N__31913));
    LocalMux I__7276 (
            .O(N__31973),
            .I(N__31908));
    LocalMux I__7275 (
            .O(N__31970),
            .I(N__31908));
    InMux I__7274 (
            .O(N__31969),
            .I(N__31901));
    InMux I__7273 (
            .O(N__31968),
            .I(N__31901));
    InMux I__7272 (
            .O(N__31967),
            .I(N__31901));
    LocalMux I__7271 (
            .O(N__31964),
            .I(N__31896));
    LocalMux I__7270 (
            .O(N__31961),
            .I(N__31896));
    InMux I__7269 (
            .O(N__31960),
            .I(N__31891));
    InMux I__7268 (
            .O(N__31959),
            .I(N__31891));
    IoInMux I__7267 (
            .O(N__31958),
            .I(N__31886));
    LocalMux I__7266 (
            .O(N__31955),
            .I(N__31882));
    LocalMux I__7265 (
            .O(N__31952),
            .I(N__31879));
    LocalMux I__7264 (
            .O(N__31943),
            .I(N__31872));
    LocalMux I__7263 (
            .O(N__31938),
            .I(N__31872));
    LocalMux I__7262 (
            .O(N__31931),
            .I(N__31872));
    LocalMux I__7261 (
            .O(N__31928),
            .I(N__31865));
    LocalMux I__7260 (
            .O(N__31921),
            .I(N__31865));
    Span4Mux_h I__7259 (
            .O(N__31916),
            .I(N__31865));
    Span4Mux_s1_v I__7258 (
            .O(N__31913),
            .I(N__31862));
    Span4Mux_v I__7257 (
            .O(N__31908),
            .I(N__31857));
    LocalMux I__7256 (
            .O(N__31901),
            .I(N__31857));
    Span4Mux_v I__7255 (
            .O(N__31896),
            .I(N__31854));
    LocalMux I__7254 (
            .O(N__31891),
            .I(N__31851));
    InMux I__7253 (
            .O(N__31890),
            .I(N__31846));
    InMux I__7252 (
            .O(N__31889),
            .I(N__31846));
    LocalMux I__7251 (
            .O(N__31886),
            .I(N__31843));
    InMux I__7250 (
            .O(N__31885),
            .I(N__31840));
    Span4Mux_v I__7249 (
            .O(N__31882),
            .I(N__31835));
    Span4Mux_v I__7248 (
            .O(N__31879),
            .I(N__31835));
    Span12Mux_v I__7247 (
            .O(N__31872),
            .I(N__31832));
    Span4Mux_v I__7246 (
            .O(N__31865),
            .I(N__31827));
    Span4Mux_h I__7245 (
            .O(N__31862),
            .I(N__31827));
    Span4Mux_h I__7244 (
            .O(N__31857),
            .I(N__31818));
    Span4Mux_h I__7243 (
            .O(N__31854),
            .I(N__31818));
    Span4Mux_h I__7242 (
            .O(N__31851),
            .I(N__31818));
    LocalMux I__7241 (
            .O(N__31846),
            .I(N__31818));
    Odrv12 I__7240 (
            .O(N__31843),
            .I(suswarn_n));
    LocalMux I__7239 (
            .O(N__31840),
            .I(suswarn_n));
    Odrv4 I__7238 (
            .O(N__31835),
            .I(suswarn_n));
    Odrv12 I__7237 (
            .O(N__31832),
            .I(suswarn_n));
    Odrv4 I__7236 (
            .O(N__31827),
            .I(suswarn_n));
    Odrv4 I__7235 (
            .O(N__31818),
            .I(suswarn_n));
    CascadeMux I__7234 (
            .O(N__31805),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ));
    CascadeMux I__7233 (
            .O(N__31802),
            .I(N__31796));
    InMux I__7232 (
            .O(N__31801),
            .I(N__31790));
    InMux I__7231 (
            .O(N__31800),
            .I(N__31787));
    InMux I__7230 (
            .O(N__31799),
            .I(N__31784));
    InMux I__7229 (
            .O(N__31796),
            .I(N__31779));
    InMux I__7228 (
            .O(N__31795),
            .I(N__31779));
    InMux I__7227 (
            .O(N__31794),
            .I(N__31776));
    InMux I__7226 (
            .O(N__31793),
            .I(N__31773));
    LocalMux I__7225 (
            .O(N__31790),
            .I(N__31760));
    LocalMux I__7224 (
            .O(N__31787),
            .I(N__31757));
    LocalMux I__7223 (
            .O(N__31784),
            .I(N__31754));
    LocalMux I__7222 (
            .O(N__31779),
            .I(N__31751));
    LocalMux I__7221 (
            .O(N__31776),
            .I(N__31748));
    LocalMux I__7220 (
            .O(N__31773),
            .I(N__31745));
    CEMux I__7219 (
            .O(N__31772),
            .I(N__31712));
    CEMux I__7218 (
            .O(N__31771),
            .I(N__31712));
    CEMux I__7217 (
            .O(N__31770),
            .I(N__31712));
    CEMux I__7216 (
            .O(N__31769),
            .I(N__31712));
    CEMux I__7215 (
            .O(N__31768),
            .I(N__31712));
    CEMux I__7214 (
            .O(N__31767),
            .I(N__31712));
    CEMux I__7213 (
            .O(N__31766),
            .I(N__31712));
    CEMux I__7212 (
            .O(N__31765),
            .I(N__31712));
    CEMux I__7211 (
            .O(N__31764),
            .I(N__31712));
    CEMux I__7210 (
            .O(N__31763),
            .I(N__31712));
    Glb2LocalMux I__7209 (
            .O(N__31760),
            .I(N__31712));
    Glb2LocalMux I__7208 (
            .O(N__31757),
            .I(N__31712));
    Glb2LocalMux I__7207 (
            .O(N__31754),
            .I(N__31712));
    Glb2LocalMux I__7206 (
            .O(N__31751),
            .I(N__31712));
    Glb2LocalMux I__7205 (
            .O(N__31748),
            .I(N__31712));
    Glb2LocalMux I__7204 (
            .O(N__31745),
            .I(N__31712));
    GlobalMux I__7203 (
            .O(N__31712),
            .I(N__31709));
    gio2CtrlBuf I__7202 (
            .O(N__31709),
            .I(N_579_g));
    CascadeMux I__7201 (
            .O(N__31706),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_ ));
    CascadeMux I__7200 (
            .O(N__31703),
            .I(N__31700));
    InMux I__7199 (
            .O(N__31700),
            .I(N__31697));
    LocalMux I__7198 (
            .O(N__31697),
            .I(N__31693));
    InMux I__7197 (
            .O(N__31696),
            .I(N__31690));
    Odrv4 I__7196 (
            .O(N__31693),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    LocalMux I__7195 (
            .O(N__31690),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    InMux I__7194 (
            .O(N__31685),
            .I(N__31682));
    LocalMux I__7193 (
            .O(N__31682),
            .I(\VPP_VDDQ.count_2_1_6 ));
    InMux I__7192 (
            .O(N__31679),
            .I(N__31667));
    InMux I__7191 (
            .O(N__31678),
            .I(N__31667));
    InMux I__7190 (
            .O(N__31677),
            .I(N__31667));
    InMux I__7189 (
            .O(N__31676),
            .I(N__31667));
    LocalMux I__7188 (
            .O(N__31667),
            .I(N__31664));
    Odrv4 I__7187 (
            .O(N__31664),
            .I(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ));
    CascadeMux I__7186 (
            .O(N__31661),
            .I(N__31655));
    CascadeMux I__7185 (
            .O(N__31660),
            .I(N__31650));
    InMux I__7184 (
            .O(N__31659),
            .I(N__31643));
    InMux I__7183 (
            .O(N__31658),
            .I(N__31643));
    InMux I__7182 (
            .O(N__31655),
            .I(N__31643));
    InMux I__7181 (
            .O(N__31654),
            .I(N__31636));
    InMux I__7180 (
            .O(N__31653),
            .I(N__31636));
    InMux I__7179 (
            .O(N__31650),
            .I(N__31636));
    LocalMux I__7178 (
            .O(N__31643),
            .I(N__31633));
    LocalMux I__7177 (
            .O(N__31636),
            .I(N__31630));
    Span4Mux_v I__7176 (
            .O(N__31633),
            .I(N__31626));
    Span4Mux_s1_h I__7175 (
            .O(N__31630),
            .I(N__31623));
    InMux I__7174 (
            .O(N__31629),
            .I(N__31620));
    Span4Mux_v I__7173 (
            .O(N__31626),
            .I(N__31617));
    Span4Mux_v I__7172 (
            .O(N__31623),
            .I(N__31612));
    LocalMux I__7171 (
            .O(N__31620),
            .I(N__31612));
    Odrv4 I__7170 (
            .O(N__31617),
            .I(vddq_ok));
    Odrv4 I__7169 (
            .O(N__31612),
            .I(vddq_ok));
    InMux I__7168 (
            .O(N__31607),
            .I(N__31604));
    LocalMux I__7167 (
            .O(N__31604),
            .I(N__31600));
    CascadeMux I__7166 (
            .O(N__31603),
            .I(N__31596));
    Span4Mux_v I__7165 (
            .O(N__31600),
            .I(N__31592));
    InMux I__7164 (
            .O(N__31599),
            .I(N__31587));
    InMux I__7163 (
            .O(N__31596),
            .I(N__31587));
    InMux I__7162 (
            .O(N__31595),
            .I(N__31584));
    Odrv4 I__7161 (
            .O(N__31592),
            .I(N_362));
    LocalMux I__7160 (
            .O(N__31587),
            .I(N_362));
    LocalMux I__7159 (
            .O(N__31584),
            .I(N_362));
    CascadeMux I__7158 (
            .O(N__31577),
            .I(\VPP_VDDQ.count_2_1_0_cascade_ ));
    InMux I__7157 (
            .O(N__31574),
            .I(N__31570));
    InMux I__7156 (
            .O(N__31573),
            .I(N__31567));
    LocalMux I__7155 (
            .O(N__31570),
            .I(N__31562));
    LocalMux I__7154 (
            .O(N__31567),
            .I(N__31562));
    Odrv4 I__7153 (
            .O(N__31562),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    InMux I__7152 (
            .O(N__31559),
            .I(N__31556));
    LocalMux I__7151 (
            .O(N__31556),
            .I(\VPP_VDDQ.un9_clk_100khz_12 ));
    CascadeMux I__7150 (
            .O(N__31553),
            .I(\VPP_VDDQ.un9_clk_100khz_4_cascade_ ));
    InMux I__7149 (
            .O(N__31550),
            .I(N__31547));
    LocalMux I__7148 (
            .O(N__31547),
            .I(\VPP_VDDQ.un9_clk_100khz_11 ));
    CascadeMux I__7147 (
            .O(N__31544),
            .I(\VPP_VDDQ.N_47_cascade_ ));
    InMux I__7146 (
            .O(N__31541),
            .I(N__31537));
    InMux I__7145 (
            .O(N__31540),
            .I(N__31534));
    LocalMux I__7144 (
            .O(N__31537),
            .I(N__31529));
    LocalMux I__7143 (
            .O(N__31534),
            .I(N__31529));
    Span4Mux_s2_h I__7142 (
            .O(N__31529),
            .I(N__31526));
    Span4Mux_v I__7141 (
            .O(N__31526),
            .I(N__31523));
    Odrv4 I__7140 (
            .O(N__31523),
            .I(\VPP_VDDQ.count_2_RNIZ0Z_1 ));
    CascadeMux I__7139 (
            .O(N__31520),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ));
    CascadeMux I__7138 (
            .O(N__31517),
            .I(N__31514));
    InMux I__7137 (
            .O(N__31514),
            .I(N__31511));
    LocalMux I__7136 (
            .O(N__31511),
            .I(N__31507));
    InMux I__7135 (
            .O(N__31510),
            .I(N__31504));
    Span4Mux_h I__7134 (
            .O(N__31507),
            .I(N__31499));
    LocalMux I__7133 (
            .O(N__31504),
            .I(N__31499));
    Span4Mux_s3_h I__7132 (
            .O(N__31499),
            .I(N__31496));
    Span4Mux_v I__7131 (
            .O(N__31496),
            .I(N__31493));
    Odrv4 I__7130 (
            .O(N__31493),
            .I(\VPP_VDDQ.count_2_1_1 ));
    InMux I__7129 (
            .O(N__31490),
            .I(N__31487));
    LocalMux I__7128 (
            .O(N__31487),
            .I(\VPP_VDDQ.curr_state_2_0_1 ));
    CascadeMux I__7127 (
            .O(N__31484),
            .I(N__31480));
    CascadeMux I__7126 (
            .O(N__31483),
            .I(N__31477));
    InMux I__7125 (
            .O(N__31480),
            .I(N__31474));
    InMux I__7124 (
            .O(N__31477),
            .I(N__31471));
    LocalMux I__7123 (
            .O(N__31474),
            .I(N__31468));
    LocalMux I__7122 (
            .O(N__31471),
            .I(N__31465));
    Odrv4 I__7121 (
            .O(N__31468),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ));
    Odrv4 I__7120 (
            .O(N__31465),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ));
    InMux I__7119 (
            .O(N__31460),
            .I(N__31454));
    InMux I__7118 (
            .O(N__31459),
            .I(N__31454));
    LocalMux I__7117 (
            .O(N__31454),
            .I(\VPP_VDDQ.count_2_1_2 ));
    CascadeMux I__7116 (
            .O(N__31451),
            .I(\VPP_VDDQ.count_2_1_3_cascade_ ));
    InMux I__7115 (
            .O(N__31448),
            .I(N__31444));
    InMux I__7114 (
            .O(N__31447),
            .I(N__31441));
    LocalMux I__7113 (
            .O(N__31444),
            .I(N__31438));
    LocalMux I__7112 (
            .O(N__31441),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    Odrv4 I__7111 (
            .O(N__31438),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    InMux I__7110 (
            .O(N__31433),
            .I(N__31430));
    LocalMux I__7109 (
            .O(N__31430),
            .I(\VPP_VDDQ.N_385 ));
    CascadeMux I__7108 (
            .O(N__31427),
            .I(\VPP_VDDQ.N_385_cascade_ ));
    InMux I__7107 (
            .O(N__31424),
            .I(N__31420));
    InMux I__7106 (
            .O(N__31423),
            .I(N__31417));
    LocalMux I__7105 (
            .O(N__31420),
            .I(N__31414));
    LocalMux I__7104 (
            .O(N__31417),
            .I(\POWERLED.count_clkZ0Z_11 ));
    Odrv12 I__7103 (
            .O(N__31414),
            .I(\POWERLED.count_clkZ0Z_11 ));
    CascadeMux I__7102 (
            .O(N__31409),
            .I(N__31406));
    InMux I__7101 (
            .O(N__31406),
            .I(N__31400));
    InMux I__7100 (
            .O(N__31405),
            .I(N__31400));
    LocalMux I__7099 (
            .O(N__31400),
            .I(N__31397));
    Odrv4 I__7098 (
            .O(N__31397),
            .I(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ));
    InMux I__7097 (
            .O(N__31394),
            .I(N__31391));
    LocalMux I__7096 (
            .O(N__31391),
            .I(\POWERLED.count_clk_0_11 ));
    InMux I__7095 (
            .O(N__31388),
            .I(N__31385));
    LocalMux I__7094 (
            .O(N__31385),
            .I(\POWERLED.count_clk_0_12 ));
    CascadeMux I__7093 (
            .O(N__31382),
            .I(N__31379));
    InMux I__7092 (
            .O(N__31379),
            .I(N__31373));
    InMux I__7091 (
            .O(N__31378),
            .I(N__31373));
    LocalMux I__7090 (
            .O(N__31373),
            .I(N__31370));
    Odrv4 I__7089 (
            .O(N__31370),
            .I(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ));
    InMux I__7088 (
            .O(N__31367),
            .I(N__31363));
    InMux I__7087 (
            .O(N__31366),
            .I(N__31360));
    LocalMux I__7086 (
            .O(N__31363),
            .I(N__31355));
    LocalMux I__7085 (
            .O(N__31360),
            .I(N__31355));
    Odrv12 I__7084 (
            .O(N__31355),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__7083 (
            .O(N__31352),
            .I(N__31349));
    LocalMux I__7082 (
            .O(N__31349),
            .I(N__31342));
    InMux I__7081 (
            .O(N__31348),
            .I(N__31339));
    InMux I__7080 (
            .O(N__31347),
            .I(N__31332));
    InMux I__7079 (
            .O(N__31346),
            .I(N__31332));
    InMux I__7078 (
            .O(N__31345),
            .I(N__31332));
    Span4Mux_h I__7077 (
            .O(N__31342),
            .I(N__31329));
    LocalMux I__7076 (
            .O(N__31339),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__7075 (
            .O(N__31332),
            .I(\POWERLED.count_clkZ0Z_0 ));
    Odrv4 I__7074 (
            .O(N__31329),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__7073 (
            .O(N__31322),
            .I(N__31304));
    InMux I__7072 (
            .O(N__31321),
            .I(N__31304));
    InMux I__7071 (
            .O(N__31320),
            .I(N__31299));
    InMux I__7070 (
            .O(N__31319),
            .I(N__31299));
    InMux I__7069 (
            .O(N__31318),
            .I(N__31290));
    InMux I__7068 (
            .O(N__31317),
            .I(N__31290));
    InMux I__7067 (
            .O(N__31316),
            .I(N__31290));
    InMux I__7066 (
            .O(N__31315),
            .I(N__31290));
    CascadeMux I__7065 (
            .O(N__31314),
            .I(N__31287));
    InMux I__7064 (
            .O(N__31313),
            .I(N__31272));
    InMux I__7063 (
            .O(N__31312),
            .I(N__31272));
    InMux I__7062 (
            .O(N__31311),
            .I(N__31272));
    InMux I__7061 (
            .O(N__31310),
            .I(N__31272));
    InMux I__7060 (
            .O(N__31309),
            .I(N__31272));
    LocalMux I__7059 (
            .O(N__31304),
            .I(N__31265));
    LocalMux I__7058 (
            .O(N__31299),
            .I(N__31265));
    LocalMux I__7057 (
            .O(N__31290),
            .I(N__31265));
    InMux I__7056 (
            .O(N__31287),
            .I(N__31254));
    InMux I__7055 (
            .O(N__31286),
            .I(N__31254));
    InMux I__7054 (
            .O(N__31285),
            .I(N__31254));
    InMux I__7053 (
            .O(N__31284),
            .I(N__31254));
    InMux I__7052 (
            .O(N__31283),
            .I(N__31254));
    LocalMux I__7051 (
            .O(N__31272),
            .I(N__31244));
    Span4Mux_v I__7050 (
            .O(N__31265),
            .I(N__31244));
    LocalMux I__7049 (
            .O(N__31254),
            .I(N__31244));
    InMux I__7048 (
            .O(N__31253),
            .I(N__31237));
    InMux I__7047 (
            .O(N__31252),
            .I(N__31237));
    InMux I__7046 (
            .O(N__31251),
            .I(N__31237));
    Span4Mux_s3_h I__7045 (
            .O(N__31244),
            .I(N__31234));
    LocalMux I__7044 (
            .O(N__31237),
            .I(\POWERLED.func_state_RNICAC53_0_0 ));
    Odrv4 I__7043 (
            .O(N__31234),
            .I(\POWERLED.func_state_RNICAC53_0_0 ));
    InMux I__7042 (
            .O(N__31229),
            .I(N__31226));
    LocalMux I__7041 (
            .O(N__31226),
            .I(\POWERLED.count_clk_0_1 ));
    CEMux I__7040 (
            .O(N__31223),
            .I(N__31220));
    LocalMux I__7039 (
            .O(N__31220),
            .I(N__31214));
    CEMux I__7038 (
            .O(N__31219),
            .I(N__31211));
    CEMux I__7037 (
            .O(N__31218),
            .I(N__31208));
    CEMux I__7036 (
            .O(N__31217),
            .I(N__31198));
    Span4Mux_v I__7035 (
            .O(N__31214),
            .I(N__31193));
    LocalMux I__7034 (
            .O(N__31211),
            .I(N__31193));
    LocalMux I__7033 (
            .O(N__31208),
            .I(N__31188));
    CEMux I__7032 (
            .O(N__31207),
            .I(N__31183));
    InMux I__7031 (
            .O(N__31206),
            .I(N__31183));
    InMux I__7030 (
            .O(N__31205),
            .I(N__31174));
    InMux I__7029 (
            .O(N__31204),
            .I(N__31174));
    InMux I__7028 (
            .O(N__31203),
            .I(N__31174));
    InMux I__7027 (
            .O(N__31202),
            .I(N__31174));
    CEMux I__7026 (
            .O(N__31201),
            .I(N__31171));
    LocalMux I__7025 (
            .O(N__31198),
            .I(N__31166));
    Span4Mux_s2_h I__7024 (
            .O(N__31193),
            .I(N__31166));
    InMux I__7023 (
            .O(N__31192),
            .I(N__31163));
    CascadeMux I__7022 (
            .O(N__31191),
            .I(N__31157));
    Span4Mux_v I__7021 (
            .O(N__31188),
            .I(N__31152));
    LocalMux I__7020 (
            .O(N__31183),
            .I(N__31152));
    LocalMux I__7019 (
            .O(N__31174),
            .I(N__31149));
    LocalMux I__7018 (
            .O(N__31171),
            .I(N__31136));
    Span4Mux_h I__7017 (
            .O(N__31166),
            .I(N__31136));
    LocalMux I__7016 (
            .O(N__31163),
            .I(N__31136));
    InMux I__7015 (
            .O(N__31162),
            .I(N__31131));
    InMux I__7014 (
            .O(N__31161),
            .I(N__31131));
    InMux I__7013 (
            .O(N__31160),
            .I(N__31126));
    InMux I__7012 (
            .O(N__31157),
            .I(N__31126));
    Span4Mux_h I__7011 (
            .O(N__31152),
            .I(N__31123));
    Span4Mux_h I__7010 (
            .O(N__31149),
            .I(N__31120));
    InMux I__7009 (
            .O(N__31148),
            .I(N__31107));
    InMux I__7008 (
            .O(N__31147),
            .I(N__31107));
    InMux I__7007 (
            .O(N__31146),
            .I(N__31107));
    InMux I__7006 (
            .O(N__31145),
            .I(N__31107));
    InMux I__7005 (
            .O(N__31144),
            .I(N__31107));
    InMux I__7004 (
            .O(N__31143),
            .I(N__31107));
    Sp12to4 I__7003 (
            .O(N__31136),
            .I(N__31100));
    LocalMux I__7002 (
            .O(N__31131),
            .I(N__31100));
    LocalMux I__7001 (
            .O(N__31126),
            .I(N__31100));
    Odrv4 I__7000 (
            .O(N__31123),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__6999 (
            .O(N__31120),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__6998 (
            .O(N__31107),
            .I(\POWERLED.count_clk_en ));
    Odrv12 I__6997 (
            .O(N__31100),
            .I(\POWERLED.count_clk_en ));
    InMux I__6996 (
            .O(N__31091),
            .I(N__31088));
    LocalMux I__6995 (
            .O(N__31088),
            .I(\POWERLED.count_clk_RNIZ0Z_0 ));
    CascadeMux I__6994 (
            .O(N__31085),
            .I(N__31082));
    InMux I__6993 (
            .O(N__31082),
            .I(N__31079));
    LocalMux I__6992 (
            .O(N__31079),
            .I(N__31073));
    InMux I__6991 (
            .O(N__31078),
            .I(N__31070));
    InMux I__6990 (
            .O(N__31077),
            .I(N__31067));
    InMux I__6989 (
            .O(N__31076),
            .I(N__31064));
    Span4Mux_h I__6988 (
            .O(N__31073),
            .I(N__31061));
    LocalMux I__6987 (
            .O(N__31070),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__6986 (
            .O(N__31067),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__6985 (
            .O(N__31064),
            .I(\POWERLED.count_clkZ0Z_1 ));
    Odrv4 I__6984 (
            .O(N__31061),
            .I(\POWERLED.count_clkZ0Z_1 ));
    InMux I__6983 (
            .O(N__31052),
            .I(N__31048));
    InMux I__6982 (
            .O(N__31051),
            .I(N__31045));
    LocalMux I__6981 (
            .O(N__31048),
            .I(\POWERLED.N_163 ));
    LocalMux I__6980 (
            .O(N__31045),
            .I(\POWERLED.N_163 ));
    InMux I__6979 (
            .O(N__31040),
            .I(N__31036));
    InMux I__6978 (
            .O(N__31039),
            .I(N__31033));
    LocalMux I__6977 (
            .O(N__31036),
            .I(N__31029));
    LocalMux I__6976 (
            .O(N__31033),
            .I(N__31026));
    CascadeMux I__6975 (
            .O(N__31032),
            .I(N__31023));
    Span4Mux_s3_h I__6974 (
            .O(N__31029),
            .I(N__31020));
    Span4Mux_s2_h I__6973 (
            .O(N__31026),
            .I(N__31017));
    InMux I__6972 (
            .O(N__31023),
            .I(N__31014));
    Odrv4 I__6971 (
            .O(N__31020),
            .I(\POWERLED.count_clkZ0Z_5 ));
    Odrv4 I__6970 (
            .O(N__31017),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__6969 (
            .O(N__31014),
            .I(\POWERLED.count_clkZ0Z_5 ));
    CascadeMux I__6968 (
            .O(N__31007),
            .I(\POWERLED.count_clkZ0Z_1_cascade_ ));
    InMux I__6967 (
            .O(N__31004),
            .I(N__30999));
    InMux I__6966 (
            .O(N__31003),
            .I(N__30996));
    CascadeMux I__6965 (
            .O(N__31002),
            .I(N__30993));
    LocalMux I__6964 (
            .O(N__30999),
            .I(N__30990));
    LocalMux I__6963 (
            .O(N__30996),
            .I(N__30987));
    InMux I__6962 (
            .O(N__30993),
            .I(N__30984));
    Span4Mux_v I__6961 (
            .O(N__30990),
            .I(N__30981));
    Span4Mux_s2_h I__6960 (
            .O(N__30987),
            .I(N__30978));
    LocalMux I__6959 (
            .O(N__30984),
            .I(N__30975));
    Odrv4 I__6958 (
            .O(N__30981),
            .I(\POWERLED.count_clkZ0Z_9 ));
    Odrv4 I__6957 (
            .O(N__30978),
            .I(\POWERLED.count_clkZ0Z_9 ));
    Odrv4 I__6956 (
            .O(N__30975),
            .I(\POWERLED.count_clkZ0Z_9 ));
    InMux I__6955 (
            .O(N__30968),
            .I(N__30962));
    InMux I__6954 (
            .O(N__30967),
            .I(N__30962));
    LocalMux I__6953 (
            .O(N__30962),
            .I(\POWERLED.N_176 ));
    CascadeMux I__6952 (
            .O(N__30959),
            .I(\POWERLED.count_offZ0Z_0_cascade_ ));
    InMux I__6951 (
            .O(N__30956),
            .I(N__30953));
    LocalMux I__6950 (
            .O(N__30953),
            .I(\POWERLED.count_off_0_0 ));
    CascadeMux I__6949 (
            .O(N__30950),
            .I(N__30947));
    InMux I__6948 (
            .O(N__30947),
            .I(N__30943));
    InMux I__6947 (
            .O(N__30946),
            .I(N__30940));
    LocalMux I__6946 (
            .O(N__30943),
            .I(N__30935));
    LocalMux I__6945 (
            .O(N__30940),
            .I(N__30935));
    Odrv4 I__6944 (
            .O(N__30935),
            .I(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ));
    CascadeMux I__6943 (
            .O(N__30932),
            .I(N__30926));
    InMux I__6942 (
            .O(N__30931),
            .I(N__30903));
    InMux I__6941 (
            .O(N__30930),
            .I(N__30903));
    InMux I__6940 (
            .O(N__30929),
            .I(N__30903));
    InMux I__6939 (
            .O(N__30926),
            .I(N__30894));
    InMux I__6938 (
            .O(N__30925),
            .I(N__30894));
    InMux I__6937 (
            .O(N__30924),
            .I(N__30894));
    InMux I__6936 (
            .O(N__30923),
            .I(N__30894));
    InMux I__6935 (
            .O(N__30922),
            .I(N__30889));
    InMux I__6934 (
            .O(N__30921),
            .I(N__30889));
    InMux I__6933 (
            .O(N__30920),
            .I(N__30877));
    InMux I__6932 (
            .O(N__30919),
            .I(N__30877));
    InMux I__6931 (
            .O(N__30918),
            .I(N__30877));
    InMux I__6930 (
            .O(N__30917),
            .I(N__30877));
    InMux I__6929 (
            .O(N__30916),
            .I(N__30877));
    InMux I__6928 (
            .O(N__30915),
            .I(N__30864));
    InMux I__6927 (
            .O(N__30914),
            .I(N__30864));
    InMux I__6926 (
            .O(N__30913),
            .I(N__30864));
    InMux I__6925 (
            .O(N__30912),
            .I(N__30864));
    InMux I__6924 (
            .O(N__30911),
            .I(N__30864));
    InMux I__6923 (
            .O(N__30910),
            .I(N__30864));
    LocalMux I__6922 (
            .O(N__30903),
            .I(N__30848));
    LocalMux I__6921 (
            .O(N__30894),
            .I(N__30848));
    LocalMux I__6920 (
            .O(N__30889),
            .I(N__30845));
    InMux I__6919 (
            .O(N__30888),
            .I(N__30842));
    LocalMux I__6918 (
            .O(N__30877),
            .I(N__30839));
    LocalMux I__6917 (
            .O(N__30864),
            .I(N__30836));
    InMux I__6916 (
            .O(N__30863),
            .I(N__30823));
    InMux I__6915 (
            .O(N__30862),
            .I(N__30823));
    InMux I__6914 (
            .O(N__30861),
            .I(N__30823));
    InMux I__6913 (
            .O(N__30860),
            .I(N__30823));
    InMux I__6912 (
            .O(N__30859),
            .I(N__30823));
    InMux I__6911 (
            .O(N__30858),
            .I(N__30823));
    InMux I__6910 (
            .O(N__30857),
            .I(N__30812));
    InMux I__6909 (
            .O(N__30856),
            .I(N__30812));
    InMux I__6908 (
            .O(N__30855),
            .I(N__30812));
    InMux I__6907 (
            .O(N__30854),
            .I(N__30812));
    InMux I__6906 (
            .O(N__30853),
            .I(N__30812));
    Span4Mux_h I__6905 (
            .O(N__30848),
            .I(N__30809));
    Odrv12 I__6904 (
            .O(N__30845),
            .I(\POWERLED.N_116 ));
    LocalMux I__6903 (
            .O(N__30842),
            .I(\POWERLED.N_116 ));
    Odrv4 I__6902 (
            .O(N__30839),
            .I(\POWERLED.N_116 ));
    Odrv4 I__6901 (
            .O(N__30836),
            .I(\POWERLED.N_116 ));
    LocalMux I__6900 (
            .O(N__30823),
            .I(\POWERLED.N_116 ));
    LocalMux I__6899 (
            .O(N__30812),
            .I(\POWERLED.N_116 ));
    Odrv4 I__6898 (
            .O(N__30809),
            .I(\POWERLED.N_116 ));
    InMux I__6897 (
            .O(N__30794),
            .I(N__30791));
    LocalMux I__6896 (
            .O(N__30791),
            .I(\POWERLED.count_off_0_4 ));
    CEMux I__6895 (
            .O(N__30788),
            .I(N__30779));
    InMux I__6894 (
            .O(N__30787),
            .I(N__30768));
    CEMux I__6893 (
            .O(N__30786),
            .I(N__30768));
    CascadeMux I__6892 (
            .O(N__30785),
            .I(N__30762));
    CascadeMux I__6891 (
            .O(N__30784),
            .I(N__30758));
    CEMux I__6890 (
            .O(N__30783),
            .I(N__30748));
    CEMux I__6889 (
            .O(N__30782),
            .I(N__30745));
    LocalMux I__6888 (
            .O(N__30779),
            .I(N__30742));
    CascadeMux I__6887 (
            .O(N__30778),
            .I(N__30739));
    CascadeMux I__6886 (
            .O(N__30777),
            .I(N__30736));
    InMux I__6885 (
            .O(N__30776),
            .I(N__30727));
    InMux I__6884 (
            .O(N__30775),
            .I(N__30727));
    InMux I__6883 (
            .O(N__30774),
            .I(N__30727));
    InMux I__6882 (
            .O(N__30773),
            .I(N__30724));
    LocalMux I__6881 (
            .O(N__30768),
            .I(N__30721));
    InMux I__6880 (
            .O(N__30767),
            .I(N__30716));
    InMux I__6879 (
            .O(N__30766),
            .I(N__30716));
    CEMux I__6878 (
            .O(N__30765),
            .I(N__30711));
    InMux I__6877 (
            .O(N__30762),
            .I(N__30704));
    InMux I__6876 (
            .O(N__30761),
            .I(N__30704));
    InMux I__6875 (
            .O(N__30758),
            .I(N__30704));
    InMux I__6874 (
            .O(N__30757),
            .I(N__30695));
    InMux I__6873 (
            .O(N__30756),
            .I(N__30695));
    InMux I__6872 (
            .O(N__30755),
            .I(N__30695));
    InMux I__6871 (
            .O(N__30754),
            .I(N__30695));
    InMux I__6870 (
            .O(N__30753),
            .I(N__30688));
    InMux I__6869 (
            .O(N__30752),
            .I(N__30688));
    CEMux I__6868 (
            .O(N__30751),
            .I(N__30688));
    LocalMux I__6867 (
            .O(N__30748),
            .I(N__30683));
    LocalMux I__6866 (
            .O(N__30745),
            .I(N__30683));
    Span4Mux_v I__6865 (
            .O(N__30742),
            .I(N__30680));
    InMux I__6864 (
            .O(N__30739),
            .I(N__30671));
    InMux I__6863 (
            .O(N__30736),
            .I(N__30671));
    InMux I__6862 (
            .O(N__30735),
            .I(N__30671));
    InMux I__6861 (
            .O(N__30734),
            .I(N__30671));
    LocalMux I__6860 (
            .O(N__30727),
            .I(N__30668));
    LocalMux I__6859 (
            .O(N__30724),
            .I(N__30665));
    Span4Mux_v I__6858 (
            .O(N__30721),
            .I(N__30662));
    LocalMux I__6857 (
            .O(N__30716),
            .I(N__30659));
    InMux I__6856 (
            .O(N__30715),
            .I(N__30654));
    InMux I__6855 (
            .O(N__30714),
            .I(N__30654));
    LocalMux I__6854 (
            .O(N__30711),
            .I(N__30649));
    LocalMux I__6853 (
            .O(N__30704),
            .I(N__30649));
    LocalMux I__6852 (
            .O(N__30695),
            .I(N__30646));
    LocalMux I__6851 (
            .O(N__30688),
            .I(N__30643));
    Span4Mux_s3_v I__6850 (
            .O(N__30683),
            .I(N__30632));
    Span4Mux_s0_h I__6849 (
            .O(N__30680),
            .I(N__30632));
    LocalMux I__6848 (
            .O(N__30671),
            .I(N__30632));
    Span4Mux_s3_v I__6847 (
            .O(N__30668),
            .I(N__30632));
    Span4Mux_v I__6846 (
            .O(N__30665),
            .I(N__30632));
    Span4Mux_s1_h I__6845 (
            .O(N__30662),
            .I(N__30623));
    Span4Mux_v I__6844 (
            .O(N__30659),
            .I(N__30623));
    LocalMux I__6843 (
            .O(N__30654),
            .I(N__30623));
    Span4Mux_s3_v I__6842 (
            .O(N__30649),
            .I(N__30623));
    Span4Mux_s3_h I__6841 (
            .O(N__30646),
            .I(N__30620));
    Odrv12 I__6840 (
            .O(N__30643),
            .I(\POWERLED.count_off_enZ0 ));
    Odrv4 I__6839 (
            .O(N__30632),
            .I(\POWERLED.count_off_enZ0 ));
    Odrv4 I__6838 (
            .O(N__30623),
            .I(\POWERLED.count_off_enZ0 ));
    Odrv4 I__6837 (
            .O(N__30620),
            .I(\POWERLED.count_off_enZ0 ));
    InMux I__6836 (
            .O(N__30611),
            .I(N__30608));
    LocalMux I__6835 (
            .O(N__30608),
            .I(N__30605));
    Span12Mux_v I__6834 (
            .O(N__30605),
            .I(N__30602));
    Odrv12 I__6833 (
            .O(N__30602),
            .I(v33s_ok));
    InMux I__6832 (
            .O(N__30599),
            .I(N__30596));
    LocalMux I__6831 (
            .O(N__30596),
            .I(N__30593));
    Span4Mux_v I__6830 (
            .O(N__30593),
            .I(N__30590));
    Odrv4 I__6829 (
            .O(N__30590),
            .I(vccst_cpu_ok));
    CascadeMux I__6828 (
            .O(N__30587),
            .I(N__30580));
    CascadeMux I__6827 (
            .O(N__30586),
            .I(N__30577));
    InMux I__6826 (
            .O(N__30585),
            .I(N__30571));
    InMux I__6825 (
            .O(N__30584),
            .I(N__30571));
    InMux I__6824 (
            .O(N__30583),
            .I(N__30568));
    InMux I__6823 (
            .O(N__30580),
            .I(N__30565));
    InMux I__6822 (
            .O(N__30577),
            .I(N__30562));
    InMux I__6821 (
            .O(N__30576),
            .I(N__30559));
    LocalMux I__6820 (
            .O(N__30571),
            .I(N__30556));
    LocalMux I__6819 (
            .O(N__30568),
            .I(N__30551));
    LocalMux I__6818 (
            .O(N__30565),
            .I(N__30543));
    LocalMux I__6817 (
            .O(N__30562),
            .I(N__30536));
    LocalMux I__6816 (
            .O(N__30559),
            .I(N__30536));
    Span4Mux_s3_h I__6815 (
            .O(N__30556),
            .I(N__30536));
    InMux I__6814 (
            .O(N__30555),
            .I(N__30531));
    InMux I__6813 (
            .O(N__30554),
            .I(N__30531));
    Span4Mux_v I__6812 (
            .O(N__30551),
            .I(N__30528));
    InMux I__6811 (
            .O(N__30550),
            .I(N__30525));
    InMux I__6810 (
            .O(N__30549),
            .I(N__30516));
    InMux I__6809 (
            .O(N__30548),
            .I(N__30516));
    InMux I__6808 (
            .O(N__30547),
            .I(N__30510));
    InMux I__6807 (
            .O(N__30546),
            .I(N__30510));
    Span4Mux_v I__6806 (
            .O(N__30543),
            .I(N__30506));
    Span4Mux_h I__6805 (
            .O(N__30536),
            .I(N__30501));
    LocalMux I__6804 (
            .O(N__30531),
            .I(N__30501));
    Span4Mux_v I__6803 (
            .O(N__30528),
            .I(N__30498));
    LocalMux I__6802 (
            .O(N__30525),
            .I(N__30495));
    InMux I__6801 (
            .O(N__30524),
            .I(N__30488));
    InMux I__6800 (
            .O(N__30523),
            .I(N__30488));
    InMux I__6799 (
            .O(N__30522),
            .I(N__30488));
    CascadeMux I__6798 (
            .O(N__30521),
            .I(N__30485));
    LocalMux I__6797 (
            .O(N__30516),
            .I(N__30479));
    InMux I__6796 (
            .O(N__30515),
            .I(N__30476));
    LocalMux I__6795 (
            .O(N__30510),
            .I(N__30473));
    InMux I__6794 (
            .O(N__30509),
            .I(N__30470));
    Span4Mux_h I__6793 (
            .O(N__30506),
            .I(N__30465));
    Span4Mux_v I__6792 (
            .O(N__30501),
            .I(N__30465));
    Span4Mux_h I__6791 (
            .O(N__30498),
            .I(N__30458));
    Span4Mux_v I__6790 (
            .O(N__30495),
            .I(N__30458));
    LocalMux I__6789 (
            .O(N__30488),
            .I(N__30458));
    InMux I__6788 (
            .O(N__30485),
            .I(N__30453));
    InMux I__6787 (
            .O(N__30484),
            .I(N__30453));
    InMux I__6786 (
            .O(N__30483),
            .I(N__30448));
    InMux I__6785 (
            .O(N__30482),
            .I(N__30448));
    Span12Mux_s7_h I__6784 (
            .O(N__30479),
            .I(N__30441));
    LocalMux I__6783 (
            .O(N__30476),
            .I(N__30441));
    Span12Mux_s4_h I__6782 (
            .O(N__30473),
            .I(N__30441));
    LocalMux I__6781 (
            .O(N__30470),
            .I(slp_s3n_signal));
    Odrv4 I__6780 (
            .O(N__30465),
            .I(slp_s3n_signal));
    Odrv4 I__6779 (
            .O(N__30458),
            .I(slp_s3n_signal));
    LocalMux I__6778 (
            .O(N__30453),
            .I(slp_s3n_signal));
    LocalMux I__6777 (
            .O(N__30448),
            .I(slp_s3n_signal));
    Odrv12 I__6776 (
            .O(N__30441),
            .I(slp_s3n_signal));
    InMux I__6775 (
            .O(N__30428),
            .I(N__30425));
    LocalMux I__6774 (
            .O(N__30425),
            .I(N__30422));
    Span4Mux_s3_h I__6773 (
            .O(N__30422),
            .I(N__30419));
    Span4Mux_h I__6772 (
            .O(N__30419),
            .I(N__30412));
    InMux I__6771 (
            .O(N__30418),
            .I(N__30403));
    InMux I__6770 (
            .O(N__30417),
            .I(N__30403));
    InMux I__6769 (
            .O(N__30416),
            .I(N__30403));
    InMux I__6768 (
            .O(N__30415),
            .I(N__30403));
    Odrv4 I__6767 (
            .O(N__30412),
            .I(rsmrst_pwrgd_signal));
    LocalMux I__6766 (
            .O(N__30403),
            .I(rsmrst_pwrgd_signal));
    InMux I__6765 (
            .O(N__30398),
            .I(N__30395));
    LocalMux I__6764 (
            .O(N__30395),
            .I(v5s_ok));
    CascadeMux I__6763 (
            .O(N__30392),
            .I(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ));
    InMux I__6762 (
            .O(N__30389),
            .I(N__30386));
    LocalMux I__6761 (
            .O(N__30386),
            .I(N__30382));
    IoInMux I__6760 (
            .O(N__30385),
            .I(N__30379));
    Span4Mux_v I__6759 (
            .O(N__30382),
            .I(N__30376));
    LocalMux I__6758 (
            .O(N__30379),
            .I(N__30373));
    Sp12to4 I__6757 (
            .O(N__30376),
            .I(N__30370));
    Span4Mux_s0_h I__6756 (
            .O(N__30373),
            .I(N__30367));
    Span12Mux_s4_h I__6755 (
            .O(N__30370),
            .I(N__30364));
    Span4Mux_v I__6754 (
            .O(N__30367),
            .I(N__30361));
    Odrv12 I__6753 (
            .O(N__30364),
            .I(dsw_pwrok));
    Odrv4 I__6752 (
            .O(N__30361),
            .I(dsw_pwrok));
    IoInMux I__6751 (
            .O(N__30356),
            .I(N__30353));
    LocalMux I__6750 (
            .O(N__30353),
            .I(N__30350));
    Span4Mux_s1_v I__6749 (
            .O(N__30350),
            .I(N__30347));
    Span4Mux_v I__6748 (
            .O(N__30347),
            .I(N__30344));
    Span4Mux_v I__6747 (
            .O(N__30344),
            .I(N__30341));
    Odrv4 I__6746 (
            .O(N__30341),
            .I(vccin_en));
    CascadeMux I__6745 (
            .O(N__30338),
            .I(\VPP_VDDQ.delayed_vddq_okZ0_cascade_ ));
    IoInMux I__6744 (
            .O(N__30335),
            .I(N__30332));
    LocalMux I__6743 (
            .O(N__30332),
            .I(N__30329));
    Span4Mux_s2_h I__6742 (
            .O(N__30329),
            .I(N__30325));
    InMux I__6741 (
            .O(N__30328),
            .I(N__30322));
    Span4Mux_v I__6740 (
            .O(N__30325),
            .I(N__30319));
    LocalMux I__6739 (
            .O(N__30322),
            .I(N__30316));
    Span4Mux_v I__6738 (
            .O(N__30319),
            .I(N__30311));
    Span4Mux_s2_h I__6737 (
            .O(N__30316),
            .I(N__30311));
    Span4Mux_h I__6736 (
            .O(N__30311),
            .I(N__30307));
    CascadeMux I__6735 (
            .O(N__30310),
            .I(N__30303));
    Span4Mux_h I__6734 (
            .O(N__30307),
            .I(N__30299));
    IoInMux I__6733 (
            .O(N__30306),
            .I(N__30296));
    InMux I__6732 (
            .O(N__30303),
            .I(N__30293));
    InMux I__6731 (
            .O(N__30302),
            .I(N__30290));
    Span4Mux_v I__6730 (
            .O(N__30299),
            .I(N__30287));
    LocalMux I__6729 (
            .O(N__30296),
            .I(N__30280));
    LocalMux I__6728 (
            .O(N__30293),
            .I(N__30280));
    LocalMux I__6727 (
            .O(N__30290),
            .I(N__30280));
    Odrv4 I__6726 (
            .O(N__30287),
            .I(pch_pwrok));
    Odrv12 I__6725 (
            .O(N__30280),
            .I(pch_pwrok));
    IoInMux I__6724 (
            .O(N__30275),
            .I(N__30272));
    LocalMux I__6723 (
            .O(N__30272),
            .I(N__30269));
    IoSpan4Mux I__6722 (
            .O(N__30269),
            .I(N__30266));
    Span4Mux_s2_v I__6721 (
            .O(N__30266),
            .I(N__30263));
    Span4Mux_v I__6720 (
            .O(N__30263),
            .I(N__30260));
    Span4Mux_h I__6719 (
            .O(N__30260),
            .I(N__30257));
    Odrv4 I__6718 (
            .O(N__30257),
            .I(vccst_pwrgd));
    InMux I__6717 (
            .O(N__30254),
            .I(N__30251));
    LocalMux I__6716 (
            .O(N__30251),
            .I(\VPP_VDDQ.delayed_vddq_ok_en ));
    CascadeMux I__6715 (
            .O(N__30248),
            .I(\VPP_VDDQ.delayed_vddq_ok_en_cascade_ ));
    CascadeMux I__6714 (
            .O(N__30245),
            .I(N__30242));
    InMux I__6713 (
            .O(N__30242),
            .I(N__30236));
    InMux I__6712 (
            .O(N__30241),
            .I(N__30236));
    LocalMux I__6711 (
            .O(N__30236),
            .I(N__30233));
    Odrv4 I__6710 (
            .O(N__30233),
            .I(\VPP_VDDQ.delayed_vddq_ok_0 ));
    InMux I__6709 (
            .O(N__30230),
            .I(N__30218));
    InMux I__6708 (
            .O(N__30229),
            .I(N__30218));
    InMux I__6707 (
            .O(N__30228),
            .I(N__30218));
    InMux I__6706 (
            .O(N__30227),
            .I(N__30218));
    LocalMux I__6705 (
            .O(N__30218),
            .I(\VPP_VDDQ.N_53 ));
    SRMux I__6704 (
            .O(N__30215),
            .I(N__30212));
    LocalMux I__6703 (
            .O(N__30212),
            .I(N__30209));
    Sp12to4 I__6702 (
            .O(N__30209),
            .I(N__30206));
    Odrv12 I__6701 (
            .O(N__30206),
            .I(\VPP_VDDQ.N_53_i ));
    InMux I__6700 (
            .O(N__30203),
            .I(N__30200));
    LocalMux I__6699 (
            .O(N__30200),
            .I(N__30196));
    InMux I__6698 (
            .O(N__30199),
            .I(N__30193));
    Odrv4 I__6697 (
            .O(N__30196),
            .I(\POWERLED.count_offZ0Z_15 ));
    LocalMux I__6696 (
            .O(N__30193),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__6695 (
            .O(N__30188),
            .I(\POWERLED.un3_count_off_1_cry_14 ));
    InMux I__6694 (
            .O(N__30185),
            .I(N__30179));
    InMux I__6693 (
            .O(N__30184),
            .I(N__30179));
    LocalMux I__6692 (
            .O(N__30179),
            .I(N__30176));
    Odrv4 I__6691 (
            .O(N__30176),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNIB6QDZ0 ));
    InMux I__6690 (
            .O(N__30173),
            .I(N__30170));
    LocalMux I__6689 (
            .O(N__30170),
            .I(N__30167));
    Span4Mux_v I__6688 (
            .O(N__30167),
            .I(N__30164));
    Odrv4 I__6687 (
            .O(N__30164),
            .I(\POWERLED.count_off_0_14 ));
    CascadeMux I__6686 (
            .O(N__30161),
            .I(N__30157));
    InMux I__6685 (
            .O(N__30160),
            .I(N__30154));
    InMux I__6684 (
            .O(N__30157),
            .I(N__30151));
    LocalMux I__6683 (
            .O(N__30154),
            .I(N__30148));
    LocalMux I__6682 (
            .O(N__30151),
            .I(\POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0 ));
    Odrv4 I__6681 (
            .O(N__30148),
            .I(\POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0 ));
    InMux I__6680 (
            .O(N__30143),
            .I(N__30140));
    LocalMux I__6679 (
            .O(N__30140),
            .I(N__30136));
    InMux I__6678 (
            .O(N__30139),
            .I(N__30133));
    Odrv12 I__6677 (
            .O(N__30136),
            .I(\POWERLED.count_offZ0Z_14 ));
    LocalMux I__6676 (
            .O(N__30133),
            .I(\POWERLED.count_offZ0Z_14 ));
    InMux I__6675 (
            .O(N__30128),
            .I(N__30125));
    LocalMux I__6674 (
            .O(N__30125),
            .I(N__30122));
    Odrv12 I__6673 (
            .O(N__30122),
            .I(\POWERLED.count_offZ0Z_4 ));
    CascadeMux I__6672 (
            .O(N__30119),
            .I(\POWERLED.count_offZ0Z_4_cascade_ ));
    InMux I__6671 (
            .O(N__30116),
            .I(N__30113));
    LocalMux I__6670 (
            .O(N__30113),
            .I(N__30110));
    Odrv4 I__6669 (
            .O(N__30110),
            .I(\POWERLED.un34_clk_100khz_2 ));
    InMux I__6668 (
            .O(N__30107),
            .I(N__30101));
    InMux I__6667 (
            .O(N__30106),
            .I(N__30101));
    LocalMux I__6666 (
            .O(N__30101),
            .I(N__30098));
    Odrv4 I__6665 (
            .O(N__30098),
            .I(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ));
    InMux I__6664 (
            .O(N__30095),
            .I(N__30092));
    LocalMux I__6663 (
            .O(N__30092),
            .I(\POWERLED.count_off_1_3 ));
    CascadeMux I__6662 (
            .O(N__30089),
            .I(\POWERLED.count_off_1_3_cascade_ ));
    InMux I__6661 (
            .O(N__30086),
            .I(N__30080));
    InMux I__6660 (
            .O(N__30085),
            .I(N__30080));
    LocalMux I__6659 (
            .O(N__30080),
            .I(\POWERLED.count_offZ0Z_3 ));
    InMux I__6658 (
            .O(N__30077),
            .I(N__30074));
    LocalMux I__6657 (
            .O(N__30074),
            .I(N__30071));
    Odrv12 I__6656 (
            .O(N__30071),
            .I(\POWERLED.un3_count_off_1_axb_3 ));
    CascadeMux I__6655 (
            .O(N__30068),
            .I(N__30062));
    CascadeMux I__6654 (
            .O(N__30067),
            .I(N__30059));
    InMux I__6653 (
            .O(N__30066),
            .I(N__30054));
    InMux I__6652 (
            .O(N__30065),
            .I(N__30054));
    InMux I__6651 (
            .O(N__30062),
            .I(N__30051));
    InMux I__6650 (
            .O(N__30059),
            .I(N__30048));
    LocalMux I__6649 (
            .O(N__30054),
            .I(N__30043));
    LocalMux I__6648 (
            .O(N__30051),
            .I(N__30043));
    LocalMux I__6647 (
            .O(N__30048),
            .I(\POWERLED.count_offZ0Z_0 ));
    Odrv4 I__6646 (
            .O(N__30043),
            .I(\POWERLED.count_offZ0Z_0 ));
    InMux I__6645 (
            .O(N__30038),
            .I(N__30035));
    LocalMux I__6644 (
            .O(N__30035),
            .I(\POWERLED.un3_count_off_1_axb_7 ));
    InMux I__6643 (
            .O(N__30032),
            .I(N__30026));
    InMux I__6642 (
            .O(N__30031),
            .I(N__30026));
    LocalMux I__6641 (
            .O(N__30026),
            .I(\POWERLED.un3_count_off_1_cry_6_c_RNISH5FZ0 ));
    InMux I__6640 (
            .O(N__30023),
            .I(\POWERLED.un3_count_off_1_cry_6 ));
    InMux I__6639 (
            .O(N__30020),
            .I(N__30017));
    LocalMux I__6638 (
            .O(N__30017),
            .I(N__30013));
    InMux I__6637 (
            .O(N__30016),
            .I(N__30010));
    Odrv4 I__6636 (
            .O(N__30013),
            .I(\POWERLED.count_offZ0Z_8 ));
    LocalMux I__6635 (
            .O(N__30010),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__6634 (
            .O(N__30005),
            .I(N__29999));
    InMux I__6633 (
            .O(N__30004),
            .I(N__29999));
    LocalMux I__6632 (
            .O(N__29999),
            .I(\POWERLED.un3_count_off_1_cry_7_c_RNITJ6FZ0 ));
    InMux I__6631 (
            .O(N__29996),
            .I(\POWERLED.un3_count_off_1_cry_7 ));
    InMux I__6630 (
            .O(N__29993),
            .I(N__29990));
    LocalMux I__6629 (
            .O(N__29990),
            .I(N__29987));
    Span4Mux_s2_h I__6628 (
            .O(N__29987),
            .I(N__29984));
    Odrv4 I__6627 (
            .O(N__29984),
            .I(\POWERLED.un3_count_off_1_axb_9 ));
    InMux I__6626 (
            .O(N__29981),
            .I(N__29975));
    InMux I__6625 (
            .O(N__29980),
            .I(N__29975));
    LocalMux I__6624 (
            .O(N__29975),
            .I(N__29972));
    Span4Mux_v I__6623 (
            .O(N__29972),
            .I(N__29969));
    Odrv4 I__6622 (
            .O(N__29969),
            .I(\POWERLED.un3_count_off_1_cry_8_c_RNIUL7FZ0 ));
    InMux I__6621 (
            .O(N__29966),
            .I(bfn_12_5_0_));
    InMux I__6620 (
            .O(N__29963),
            .I(N__29960));
    LocalMux I__6619 (
            .O(N__29960),
            .I(N__29957));
    Span4Mux_v I__6618 (
            .O(N__29957),
            .I(N__29954));
    Sp12to4 I__6617 (
            .O(N__29954),
            .I(N__29951));
    Odrv12 I__6616 (
            .O(N__29951),
            .I(\POWERLED.count_offZ0Z_10 ));
    CascadeMux I__6615 (
            .O(N__29948),
            .I(N__29945));
    InMux I__6614 (
            .O(N__29945),
            .I(N__29939));
    InMux I__6613 (
            .O(N__29944),
            .I(N__29939));
    LocalMux I__6612 (
            .O(N__29939),
            .I(N__29936));
    Span4Mux_v I__6611 (
            .O(N__29936),
            .I(N__29933));
    Odrv4 I__6610 (
            .O(N__29933),
            .I(\POWERLED.un3_count_off_1_cry_9_c_RNIVN8FZ0 ));
    InMux I__6609 (
            .O(N__29930),
            .I(\POWERLED.un3_count_off_1_cry_9 ));
    InMux I__6608 (
            .O(N__29927),
            .I(N__29924));
    LocalMux I__6607 (
            .O(N__29924),
            .I(\POWERLED.un3_count_off_1_axb_11 ));
    InMux I__6606 (
            .O(N__29921),
            .I(N__29915));
    InMux I__6605 (
            .O(N__29920),
            .I(N__29915));
    LocalMux I__6604 (
            .O(N__29915),
            .I(\POWERLED.un3_count_off_1_cry_10_c_RNI7ULDZ0 ));
    InMux I__6603 (
            .O(N__29912),
            .I(\POWERLED.un3_count_off_1_cry_10 ));
    InMux I__6602 (
            .O(N__29909),
            .I(N__29906));
    LocalMux I__6601 (
            .O(N__29906),
            .I(N__29902));
    InMux I__6600 (
            .O(N__29905),
            .I(N__29899));
    Span4Mux_v I__6599 (
            .O(N__29902),
            .I(N__29896));
    LocalMux I__6598 (
            .O(N__29899),
            .I(N__29893));
    Odrv4 I__6597 (
            .O(N__29896),
            .I(\POWERLED.count_offZ0Z_12 ));
    Odrv4 I__6596 (
            .O(N__29893),
            .I(\POWERLED.count_offZ0Z_12 ));
    CascadeMux I__6595 (
            .O(N__29888),
            .I(N__29885));
    InMux I__6594 (
            .O(N__29885),
            .I(N__29879));
    InMux I__6593 (
            .O(N__29884),
            .I(N__29879));
    LocalMux I__6592 (
            .O(N__29879),
            .I(N__29876));
    Odrv4 I__6591 (
            .O(N__29876),
            .I(\POWERLED.un3_count_off_1_cry_11_c_RNI80NDZ0 ));
    InMux I__6590 (
            .O(N__29873),
            .I(\POWERLED.un3_count_off_1_cry_11 ));
    InMux I__6589 (
            .O(N__29870),
            .I(N__29867));
    LocalMux I__6588 (
            .O(N__29867),
            .I(N__29864));
    Odrv4 I__6587 (
            .O(N__29864),
            .I(\POWERLED.count_offZ0Z_13 ));
    CascadeMux I__6586 (
            .O(N__29861),
            .I(N__29858));
    InMux I__6585 (
            .O(N__29858),
            .I(N__29852));
    InMux I__6584 (
            .O(N__29857),
            .I(N__29852));
    LocalMux I__6583 (
            .O(N__29852),
            .I(N__29849));
    Odrv12 I__6582 (
            .O(N__29849),
            .I(\POWERLED.un3_count_off_1_cry_12_c_RNI92ODZ0 ));
    InMux I__6581 (
            .O(N__29846),
            .I(\POWERLED.un3_count_off_1_cry_12 ));
    InMux I__6580 (
            .O(N__29843),
            .I(\POWERLED.un3_count_off_1_cry_13 ));
    InMux I__6579 (
            .O(N__29840),
            .I(N__29837));
    LocalMux I__6578 (
            .O(N__29837),
            .I(\POWERLED.count_off_0_13 ));
    CascadeMux I__6577 (
            .O(N__29834),
            .I(\POWERLED.count_offZ0Z_13_cascade_ ));
    InMux I__6576 (
            .O(N__29831),
            .I(N__29828));
    LocalMux I__6575 (
            .O(N__29828),
            .I(N__29825));
    Span4Mux_h I__6574 (
            .O(N__29825),
            .I(N__29822));
    Odrv4 I__6573 (
            .O(N__29822),
            .I(\POWERLED.un34_clk_100khz_11 ));
    InMux I__6572 (
            .O(N__29819),
            .I(N__29814));
    InMux I__6571 (
            .O(N__29818),
            .I(N__29811));
    InMux I__6570 (
            .O(N__29817),
            .I(N__29808));
    LocalMux I__6569 (
            .O(N__29814),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__6568 (
            .O(N__29811),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__6567 (
            .O(N__29808),
            .I(\POWERLED.count_offZ0Z_1 ));
    InMux I__6566 (
            .O(N__29801),
            .I(N__29798));
    LocalMux I__6565 (
            .O(N__29798),
            .I(\POWERLED.un3_count_off_1_axb_2 ));
    InMux I__6564 (
            .O(N__29795),
            .I(N__29789));
    InMux I__6563 (
            .O(N__29794),
            .I(N__29789));
    LocalMux I__6562 (
            .O(N__29789),
            .I(\POWERLED.un3_count_off_1_cry_1_c_RNIN70FZ0 ));
    InMux I__6561 (
            .O(N__29786),
            .I(\POWERLED.un3_count_off_1_cry_1 ));
    InMux I__6560 (
            .O(N__29783),
            .I(\POWERLED.un3_count_off_1_cry_2 ));
    InMux I__6559 (
            .O(N__29780),
            .I(\POWERLED.un3_count_off_1_cry_3 ));
    CascadeMux I__6558 (
            .O(N__29777),
            .I(N__29773));
    InMux I__6557 (
            .O(N__29776),
            .I(N__29770));
    InMux I__6556 (
            .O(N__29773),
            .I(N__29767));
    LocalMux I__6555 (
            .O(N__29770),
            .I(\POWERLED.count_offZ0Z_5 ));
    LocalMux I__6554 (
            .O(N__29767),
            .I(\POWERLED.count_offZ0Z_5 ));
    CascadeMux I__6553 (
            .O(N__29762),
            .I(N__29758));
    InMux I__6552 (
            .O(N__29761),
            .I(N__29753));
    InMux I__6551 (
            .O(N__29758),
            .I(N__29753));
    LocalMux I__6550 (
            .O(N__29753),
            .I(\POWERLED.un3_count_off_1_cry_4_c_RNIQD3FZ0 ));
    InMux I__6549 (
            .O(N__29750),
            .I(\POWERLED.un3_count_off_1_cry_4 ));
    InMux I__6548 (
            .O(N__29747),
            .I(N__29744));
    LocalMux I__6547 (
            .O(N__29744),
            .I(\POWERLED.un3_count_off_1_axb_6 ));
    InMux I__6546 (
            .O(N__29741),
            .I(N__29737));
    InMux I__6545 (
            .O(N__29740),
            .I(N__29734));
    LocalMux I__6544 (
            .O(N__29737),
            .I(\POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0 ));
    LocalMux I__6543 (
            .O(N__29734),
            .I(\POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0 ));
    InMux I__6542 (
            .O(N__29729),
            .I(\POWERLED.un3_count_off_1_cry_5 ));
    InMux I__6541 (
            .O(N__29726),
            .I(N__29722));
    InMux I__6540 (
            .O(N__29725),
            .I(N__29719));
    LocalMux I__6539 (
            .O(N__29722),
            .I(\VPP_VDDQ.N_186 ));
    LocalMux I__6538 (
            .O(N__29719),
            .I(\VPP_VDDQ.N_186 ));
    CascadeMux I__6537 (
            .O(N__29714),
            .I(N__29711));
    InMux I__6536 (
            .O(N__29711),
            .I(N__29708));
    LocalMux I__6535 (
            .O(N__29708),
            .I(\VPP_VDDQ.N_214 ));
    InMux I__6534 (
            .O(N__29705),
            .I(N__29701));
    InMux I__6533 (
            .O(N__29704),
            .I(N__29698));
    LocalMux I__6532 (
            .O(N__29701),
            .I(N__29695));
    LocalMux I__6531 (
            .O(N__29698),
            .I(N__29692));
    Span4Mux_v I__6530 (
            .O(N__29695),
            .I(N__29689));
    Span4Mux_s3_h I__6529 (
            .O(N__29692),
            .I(N__29686));
    Odrv4 I__6528 (
            .O(N__29689),
            .I(\VPP_VDDQ.un6_count ));
    Odrv4 I__6527 (
            .O(N__29686),
            .I(\VPP_VDDQ.un6_count ));
    InMux I__6526 (
            .O(N__29681),
            .I(N__29676));
    InMux I__6525 (
            .O(N__29680),
            .I(N__29668));
    InMux I__6524 (
            .O(N__29679),
            .I(N__29668));
    LocalMux I__6523 (
            .O(N__29676),
            .I(N__29665));
    InMux I__6522 (
            .O(N__29675),
            .I(N__29658));
    InMux I__6521 (
            .O(N__29674),
            .I(N__29658));
    InMux I__6520 (
            .O(N__29673),
            .I(N__29658));
    LocalMux I__6519 (
            .O(N__29668),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    Odrv4 I__6518 (
            .O(N__29665),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__6517 (
            .O(N__29658),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    CascadeMux I__6516 (
            .O(N__29651),
            .I(N__29647));
    InMux I__6515 (
            .O(N__29650),
            .I(N__29641));
    InMux I__6514 (
            .O(N__29647),
            .I(N__29641));
    InMux I__6513 (
            .O(N__29646),
            .I(N__29637));
    LocalMux I__6512 (
            .O(N__29641),
            .I(N__29634));
    InMux I__6511 (
            .O(N__29640),
            .I(N__29631));
    LocalMux I__6510 (
            .O(N__29637),
            .I(\VPP_VDDQ.N_360 ));
    Odrv4 I__6509 (
            .O(N__29634),
            .I(\VPP_VDDQ.N_360 ));
    LocalMux I__6508 (
            .O(N__29631),
            .I(\VPP_VDDQ.N_360 ));
    CascadeMux I__6507 (
            .O(N__29624),
            .I(N__29621));
    InMux I__6506 (
            .O(N__29621),
            .I(N__29611));
    InMux I__6505 (
            .O(N__29620),
            .I(N__29611));
    InMux I__6504 (
            .O(N__29619),
            .I(N__29608));
    InMux I__6503 (
            .O(N__29618),
            .I(N__29601));
    InMux I__6502 (
            .O(N__29617),
            .I(N__29601));
    InMux I__6501 (
            .O(N__29616),
            .I(N__29601));
    LocalMux I__6500 (
            .O(N__29611),
            .I(N__29598));
    LocalMux I__6499 (
            .O(N__29608),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__6498 (
            .O(N__29601),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    Odrv4 I__6497 (
            .O(N__29598),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    InMux I__6496 (
            .O(N__29591),
            .I(N__29530));
    InMux I__6495 (
            .O(N__29590),
            .I(N__29530));
    InMux I__6494 (
            .O(N__29589),
            .I(N__29530));
    InMux I__6493 (
            .O(N__29588),
            .I(N__29530));
    InMux I__6492 (
            .O(N__29587),
            .I(N__29521));
    InMux I__6491 (
            .O(N__29586),
            .I(N__29521));
    InMux I__6490 (
            .O(N__29585),
            .I(N__29521));
    InMux I__6489 (
            .O(N__29584),
            .I(N__29521));
    InMux I__6488 (
            .O(N__29583),
            .I(N__29512));
    InMux I__6487 (
            .O(N__29582),
            .I(N__29512));
    InMux I__6486 (
            .O(N__29581),
            .I(N__29512));
    InMux I__6485 (
            .O(N__29580),
            .I(N__29512));
    InMux I__6484 (
            .O(N__29579),
            .I(N__29505));
    InMux I__6483 (
            .O(N__29578),
            .I(N__29505));
    InMux I__6482 (
            .O(N__29577),
            .I(N__29505));
    InMux I__6481 (
            .O(N__29576),
            .I(N__29500));
    InMux I__6480 (
            .O(N__29575),
            .I(N__29500));
    InMux I__6479 (
            .O(N__29574),
            .I(N__29491));
    InMux I__6478 (
            .O(N__29573),
            .I(N__29491));
    InMux I__6477 (
            .O(N__29572),
            .I(N__29491));
    InMux I__6476 (
            .O(N__29571),
            .I(N__29491));
    InMux I__6475 (
            .O(N__29570),
            .I(N__29484));
    InMux I__6474 (
            .O(N__29569),
            .I(N__29484));
    InMux I__6473 (
            .O(N__29568),
            .I(N__29484));
    InMux I__6472 (
            .O(N__29567),
            .I(N__29475));
    InMux I__6471 (
            .O(N__29566),
            .I(N__29475));
    InMux I__6470 (
            .O(N__29565),
            .I(N__29475));
    InMux I__6469 (
            .O(N__29564),
            .I(N__29475));
    InMux I__6468 (
            .O(N__29563),
            .I(N__29468));
    InMux I__6467 (
            .O(N__29562),
            .I(N__29468));
    InMux I__6466 (
            .O(N__29561),
            .I(N__29468));
    InMux I__6465 (
            .O(N__29560),
            .I(N__29459));
    InMux I__6464 (
            .O(N__29559),
            .I(N__29459));
    InMux I__6463 (
            .O(N__29558),
            .I(N__29459));
    InMux I__6462 (
            .O(N__29557),
            .I(N__29459));
    InMux I__6461 (
            .O(N__29556),
            .I(N__29450));
    InMux I__6460 (
            .O(N__29555),
            .I(N__29450));
    InMux I__6459 (
            .O(N__29554),
            .I(N__29450));
    InMux I__6458 (
            .O(N__29553),
            .I(N__29450));
    InMux I__6457 (
            .O(N__29552),
            .I(N__29441));
    InMux I__6456 (
            .O(N__29551),
            .I(N__29441));
    InMux I__6455 (
            .O(N__29550),
            .I(N__29441));
    InMux I__6454 (
            .O(N__29549),
            .I(N__29441));
    InMux I__6453 (
            .O(N__29548),
            .I(N__29436));
    InMux I__6452 (
            .O(N__29547),
            .I(N__29436));
    InMux I__6451 (
            .O(N__29546),
            .I(N__29427));
    InMux I__6450 (
            .O(N__29545),
            .I(N__29427));
    InMux I__6449 (
            .O(N__29544),
            .I(N__29427));
    InMux I__6448 (
            .O(N__29543),
            .I(N__29427));
    InMux I__6447 (
            .O(N__29542),
            .I(N__29422));
    InMux I__6446 (
            .O(N__29541),
            .I(N__29422));
    InMux I__6445 (
            .O(N__29540),
            .I(N__29417));
    InMux I__6444 (
            .O(N__29539),
            .I(N__29417));
    LocalMux I__6443 (
            .O(N__29530),
            .I(N__29412));
    LocalMux I__6442 (
            .O(N__29521),
            .I(N__29409));
    LocalMux I__6441 (
            .O(N__29512),
            .I(N__29405));
    LocalMux I__6440 (
            .O(N__29505),
            .I(N__29402));
    LocalMux I__6439 (
            .O(N__29500),
            .I(N__29398));
    LocalMux I__6438 (
            .O(N__29491),
            .I(N__29392));
    LocalMux I__6437 (
            .O(N__29484),
            .I(N__29389));
    LocalMux I__6436 (
            .O(N__29475),
            .I(N__29386));
    LocalMux I__6435 (
            .O(N__29468),
            .I(N__29383));
    LocalMux I__6434 (
            .O(N__29459),
            .I(N__29380));
    LocalMux I__6433 (
            .O(N__29450),
            .I(N__29377));
    LocalMux I__6432 (
            .O(N__29441),
            .I(N__29374));
    LocalMux I__6431 (
            .O(N__29436),
            .I(N__29371));
    LocalMux I__6430 (
            .O(N__29427),
            .I(N__29368));
    LocalMux I__6429 (
            .O(N__29422),
            .I(N__29365));
    LocalMux I__6428 (
            .O(N__29417),
            .I(N__29362));
    CEMux I__6427 (
            .O(N__29416),
            .I(N__29315));
    CEMux I__6426 (
            .O(N__29415),
            .I(N__29315));
    Glb2LocalMux I__6425 (
            .O(N__29412),
            .I(N__29315));
    Glb2LocalMux I__6424 (
            .O(N__29409),
            .I(N__29315));
    CEMux I__6423 (
            .O(N__29408),
            .I(N__29315));
    Glb2LocalMux I__6422 (
            .O(N__29405),
            .I(N__29315));
    Glb2LocalMux I__6421 (
            .O(N__29402),
            .I(N__29315));
    CEMux I__6420 (
            .O(N__29401),
            .I(N__29315));
    Glb2LocalMux I__6419 (
            .O(N__29398),
            .I(N__29315));
    CEMux I__6418 (
            .O(N__29397),
            .I(N__29315));
    CEMux I__6417 (
            .O(N__29396),
            .I(N__29315));
    CEMux I__6416 (
            .O(N__29395),
            .I(N__29315));
    Glb2LocalMux I__6415 (
            .O(N__29392),
            .I(N__29315));
    Glb2LocalMux I__6414 (
            .O(N__29389),
            .I(N__29315));
    Glb2LocalMux I__6413 (
            .O(N__29386),
            .I(N__29315));
    Glb2LocalMux I__6412 (
            .O(N__29383),
            .I(N__29315));
    Glb2LocalMux I__6411 (
            .O(N__29380),
            .I(N__29315));
    Glb2LocalMux I__6410 (
            .O(N__29377),
            .I(N__29315));
    Glb2LocalMux I__6409 (
            .O(N__29374),
            .I(N__29315));
    Glb2LocalMux I__6408 (
            .O(N__29371),
            .I(N__29315));
    Glb2LocalMux I__6407 (
            .O(N__29368),
            .I(N__29315));
    Glb2LocalMux I__6406 (
            .O(N__29365),
            .I(N__29315));
    Glb2LocalMux I__6405 (
            .O(N__29362),
            .I(N__29315));
    GlobalMux I__6404 (
            .O(N__29315),
            .I(N__29312));
    gio2CtrlBuf I__6403 (
            .O(N__29312),
            .I(N_27_g));
    CascadeMux I__6402 (
            .O(N__29309),
            .I(\POWERLED.count_off_RNIZ0Z_1_cascade_ ));
    InMux I__6401 (
            .O(N__29306),
            .I(N__29303));
    LocalMux I__6400 (
            .O(N__29303),
            .I(\POWERLED.count_off_0_12 ));
    InMux I__6399 (
            .O(N__29300),
            .I(N__29297));
    LocalMux I__6398 (
            .O(N__29297),
            .I(\POWERLED.count_off_RNIZ0Z_1 ));
    InMux I__6397 (
            .O(N__29294),
            .I(N__29291));
    LocalMux I__6396 (
            .O(N__29291),
            .I(\POWERLED.count_off_0_1 ));
    IoInMux I__6395 (
            .O(N__29288),
            .I(N__29285));
    LocalMux I__6394 (
            .O(N__29285),
            .I(N__29282));
    IoSpan4Mux I__6393 (
            .O(N__29282),
            .I(N__29279));
    Odrv4 I__6392 (
            .O(N__29279),
            .I(vpp_en));
    InMux I__6391 (
            .O(N__29276),
            .I(N__29273));
    LocalMux I__6390 (
            .O(N__29273),
            .I(N__29270));
    Span4Mux_v I__6389 (
            .O(N__29270),
            .I(N__29264));
    IoInMux I__6388 (
            .O(N__29269),
            .I(N__29261));
    InMux I__6387 (
            .O(N__29268),
            .I(N__29256));
    InMux I__6386 (
            .O(N__29267),
            .I(N__29256));
    IoSpan4Mux I__6385 (
            .O(N__29264),
            .I(N__29251));
    LocalMux I__6384 (
            .O(N__29261),
            .I(N__29251));
    LocalMux I__6383 (
            .O(N__29256),
            .I(N__29246));
    IoSpan4Mux I__6382 (
            .O(N__29251),
            .I(N__29243));
    CascadeMux I__6381 (
            .O(N__29250),
            .I(N__29239));
    InMux I__6380 (
            .O(N__29249),
            .I(N__29235));
    Span4Mux_s3_v I__6379 (
            .O(N__29246),
            .I(N__29232));
    Span4Mux_s0_h I__6378 (
            .O(N__29243),
            .I(N__29228));
    InMux I__6377 (
            .O(N__29242),
            .I(N__29225));
    InMux I__6376 (
            .O(N__29239),
            .I(N__29222));
    CascadeMux I__6375 (
            .O(N__29238),
            .I(N__29219));
    LocalMux I__6374 (
            .O(N__29235),
            .I(N__29216));
    Span4Mux_v I__6373 (
            .O(N__29232),
            .I(N__29213));
    InMux I__6372 (
            .O(N__29231),
            .I(N__29210));
    Span4Mux_h I__6371 (
            .O(N__29228),
            .I(N__29207));
    LocalMux I__6370 (
            .O(N__29225),
            .I(N__29202));
    LocalMux I__6369 (
            .O(N__29222),
            .I(N__29202));
    InMux I__6368 (
            .O(N__29219),
            .I(N__29197));
    Span4Mux_v I__6367 (
            .O(N__29216),
            .I(N__29190));
    Span4Mux_v I__6366 (
            .O(N__29213),
            .I(N__29190));
    LocalMux I__6365 (
            .O(N__29210),
            .I(N__29190));
    Span4Mux_h I__6364 (
            .O(N__29207),
            .I(N__29185));
    Span4Mux_h I__6363 (
            .O(N__29202),
            .I(N__29185));
    InMux I__6362 (
            .O(N__29201),
            .I(N__29182));
    InMux I__6361 (
            .O(N__29200),
            .I(N__29179));
    LocalMux I__6360 (
            .O(N__29197),
            .I(N__29176));
    Odrv4 I__6359 (
            .O(N__29190),
            .I(vccst_en));
    Odrv4 I__6358 (
            .O(N__29185),
            .I(vccst_en));
    LocalMux I__6357 (
            .O(N__29182),
            .I(vccst_en));
    LocalMux I__6356 (
            .O(N__29179),
            .I(vccst_en));
    Odrv4 I__6355 (
            .O(N__29176),
            .I(vccst_en));
    CascadeMux I__6354 (
            .O(N__29165),
            .I(\VPP_VDDQ.N_360_cascade_ ));
    CascadeMux I__6353 (
            .O(N__29162),
            .I(N__29158));
    InMux I__6352 (
            .O(N__29161),
            .I(N__29155));
    InMux I__6351 (
            .O(N__29158),
            .I(N__29152));
    LocalMux I__6350 (
            .O(N__29155),
            .I(N__29147));
    LocalMux I__6349 (
            .O(N__29152),
            .I(N__29147));
    Span4Mux_h I__6348 (
            .O(N__29147),
            .I(N__29144));
    Odrv4 I__6347 (
            .O(N__29144),
            .I(\VPP_VDDQ.N_264_i ));
    CascadeMux I__6346 (
            .O(N__29141),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ));
    InMux I__6345 (
            .O(N__29138),
            .I(N__29132));
    InMux I__6344 (
            .O(N__29137),
            .I(N__29132));
    LocalMux I__6343 (
            .O(N__29132),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    SRMux I__6342 (
            .O(N__29129),
            .I(N__29125));
    SRMux I__6341 (
            .O(N__29128),
            .I(N__29122));
    LocalMux I__6340 (
            .O(N__29125),
            .I(N__29118));
    LocalMux I__6339 (
            .O(N__29122),
            .I(N__29115));
    SRMux I__6338 (
            .O(N__29121),
            .I(N__29112));
    Span4Mux_h I__6337 (
            .O(N__29118),
            .I(N__29109));
    Span4Mux_v I__6336 (
            .O(N__29115),
            .I(N__29106));
    LocalMux I__6335 (
            .O(N__29112),
            .I(N__29103));
    Odrv4 I__6334 (
            .O(N__29109),
            .I(\VPP_VDDQ.curr_state_RNITROD7Z0Z_0 ));
    Odrv4 I__6333 (
            .O(N__29106),
            .I(\VPP_VDDQ.curr_state_RNITROD7Z0Z_0 ));
    Odrv12 I__6332 (
            .O(N__29103),
            .I(\VPP_VDDQ.curr_state_RNITROD7Z0Z_0 ));
    CascadeMux I__6331 (
            .O(N__29096),
            .I(\VPP_VDDQ.curr_state_RNITROD7Z0Z_0_cascade_ ));
    CEMux I__6330 (
            .O(N__29093),
            .I(N__29090));
    LocalMux I__6329 (
            .O(N__29090),
            .I(N__29087));
    Odrv4 I__6328 (
            .O(N__29087),
            .I(\VPP_VDDQ.N_27_0 ));
    InMux I__6327 (
            .O(N__29084),
            .I(N__29081));
    LocalMux I__6326 (
            .O(N__29081),
            .I(\VPP_VDDQ.N_382 ));
    InMux I__6325 (
            .O(N__29078),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13 ));
    InMux I__6324 (
            .O(N__29075),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14 ));
    InMux I__6323 (
            .O(N__29072),
            .I(N__29066));
    InMux I__6322 (
            .O(N__29071),
            .I(N__29066));
    LocalMux I__6321 (
            .O(N__29066),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    CascadeMux I__6320 (
            .O(N__29063),
            .I(\VPP_VDDQ.count_2_1_13_cascade_ ));
    InMux I__6319 (
            .O(N__29060),
            .I(N__29057));
    LocalMux I__6318 (
            .O(N__29057),
            .I(\VPP_VDDQ.count_2_0_13 ));
    CascadeMux I__6317 (
            .O(N__29054),
            .I(N__29050));
    InMux I__6316 (
            .O(N__29053),
            .I(N__29045));
    InMux I__6315 (
            .O(N__29050),
            .I(N__29045));
    LocalMux I__6314 (
            .O(N__29045),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    CascadeMux I__6313 (
            .O(N__29042),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ));
    CascadeMux I__6312 (
            .O(N__29039),
            .I(N__29035));
    InMux I__6311 (
            .O(N__29038),
            .I(N__29030));
    InMux I__6310 (
            .O(N__29035),
            .I(N__29030));
    LocalMux I__6309 (
            .O(N__29030),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    InMux I__6308 (
            .O(N__29027),
            .I(N__29021));
    InMux I__6307 (
            .O(N__29026),
            .I(N__29021));
    LocalMux I__6306 (
            .O(N__29021),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ));
    InMux I__6305 (
            .O(N__29018),
            .I(N__29015));
    LocalMux I__6304 (
            .O(N__29015),
            .I(\VPP_VDDQ.count_2_0_15 ));
    InMux I__6303 (
            .O(N__29012),
            .I(N__29009));
    LocalMux I__6302 (
            .O(N__29009),
            .I(\VPP_VDDQ.un1_count_2_1_axb_5 ));
    InMux I__6301 (
            .O(N__29006),
            .I(N__29003));
    LocalMux I__6300 (
            .O(N__29003),
            .I(N__28999));
    InMux I__6299 (
            .O(N__29002),
            .I(N__28996));
    Odrv4 I__6298 (
            .O(N__28999),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ));
    LocalMux I__6297 (
            .O(N__28996),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ));
    InMux I__6296 (
            .O(N__28991),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4 ));
    InMux I__6295 (
            .O(N__28988),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5 ));
    InMux I__6294 (
            .O(N__28985),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6 ));
    InMux I__6293 (
            .O(N__28982),
            .I(N__28978));
    InMux I__6292 (
            .O(N__28981),
            .I(N__28975));
    LocalMux I__6291 (
            .O(N__28978),
            .I(N__28972));
    LocalMux I__6290 (
            .O(N__28975),
            .I(N__28969));
    Span4Mux_s2_h I__6289 (
            .O(N__28972),
            .I(N__28966));
    Span4Mux_s2_h I__6288 (
            .O(N__28969),
            .I(N__28963));
    Span4Mux_v I__6287 (
            .O(N__28966),
            .I(N__28960));
    Span4Mux_v I__6286 (
            .O(N__28963),
            .I(N__28957));
    Odrv4 I__6285 (
            .O(N__28960),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    Odrv4 I__6284 (
            .O(N__28957),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    InMux I__6283 (
            .O(N__28952),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7 ));
    CascadeMux I__6282 (
            .O(N__28949),
            .I(N__28945));
    InMux I__6281 (
            .O(N__28948),
            .I(N__28940));
    InMux I__6280 (
            .O(N__28945),
            .I(N__28940));
    LocalMux I__6279 (
            .O(N__28940),
            .I(N__28937));
    Odrv4 I__6278 (
            .O(N__28937),
            .I(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ));
    InMux I__6277 (
            .O(N__28934),
            .I(bfn_11_12_0_));
    InMux I__6276 (
            .O(N__28931),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9 ));
    InMux I__6275 (
            .O(N__28928),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10 ));
    InMux I__6274 (
            .O(N__28925),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11 ));
    InMux I__6273 (
            .O(N__28922),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12 ));
    CascadeMux I__6272 (
            .O(N__28919),
            .I(N__28915));
    InMux I__6271 (
            .O(N__28918),
            .I(N__28910));
    InMux I__6270 (
            .O(N__28915),
            .I(N__28910));
    LocalMux I__6269 (
            .O(N__28910),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    InMux I__6268 (
            .O(N__28907),
            .I(N__28901));
    InMux I__6267 (
            .O(N__28906),
            .I(N__28901));
    LocalMux I__6266 (
            .O(N__28901),
            .I(\VPP_VDDQ.count_2_1_4 ));
    InMux I__6265 (
            .O(N__28898),
            .I(N__28895));
    LocalMux I__6264 (
            .O(N__28895),
            .I(\VPP_VDDQ.count_2_1_5 ));
    CascadeMux I__6263 (
            .O(N__28892),
            .I(\VPP_VDDQ.count_2_1_5_cascade_ ));
    CascadeMux I__6262 (
            .O(N__28889),
            .I(N__28886));
    InMux I__6261 (
            .O(N__28886),
            .I(N__28880));
    InMux I__6260 (
            .O(N__28885),
            .I(N__28880));
    LocalMux I__6259 (
            .O(N__28880),
            .I(N__28877));
    Odrv12 I__6258 (
            .O(N__28877),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    CascadeMux I__6257 (
            .O(N__28874),
            .I(N__28871));
    InMux I__6256 (
            .O(N__28871),
            .I(N__28865));
    InMux I__6255 (
            .O(N__28870),
            .I(N__28865));
    LocalMux I__6254 (
            .O(N__28865),
            .I(\VPP_VDDQ.count_2Z0Z_2 ));
    CascadeMux I__6253 (
            .O(N__28862),
            .I(N__28859));
    InMux I__6252 (
            .O(N__28859),
            .I(N__28856));
    LocalMux I__6251 (
            .O(N__28856),
            .I(N__28853));
    Span4Mux_v I__6250 (
            .O(N__28853),
            .I(N__28850));
    Span4Mux_v I__6249 (
            .O(N__28850),
            .I(N__28847));
    Odrv4 I__6248 (
            .O(N__28847),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    InMux I__6247 (
            .O(N__28844),
            .I(N__28841));
    LocalMux I__6246 (
            .O(N__28841),
            .I(\VPP_VDDQ.un1_count_2_1_axb_2 ));
    InMux I__6245 (
            .O(N__28838),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1 ));
    InMux I__6244 (
            .O(N__28835),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2 ));
    InMux I__6243 (
            .O(N__28832),
            .I(N__28829));
    LocalMux I__6242 (
            .O(N__28829),
            .I(\VPP_VDDQ.un1_count_2_1_axb_4 ));
    CascadeMux I__6241 (
            .O(N__28826),
            .I(N__28823));
    InMux I__6240 (
            .O(N__28823),
            .I(N__28817));
    InMux I__6239 (
            .O(N__28822),
            .I(N__28817));
    LocalMux I__6238 (
            .O(N__28817),
            .I(N__28814));
    Odrv4 I__6237 (
            .O(N__28814),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ));
    InMux I__6236 (
            .O(N__28811),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3 ));
    CascadeMux I__6235 (
            .O(N__28808),
            .I(\VPP_VDDQ.count_2_1_9_cascade_ ));
    InMux I__6234 (
            .O(N__28805),
            .I(N__28802));
    LocalMux I__6233 (
            .O(N__28802),
            .I(\VPP_VDDQ.count_2_0_9 ));
    InMux I__6232 (
            .O(N__28799),
            .I(N__28796));
    LocalMux I__6231 (
            .O(N__28796),
            .I(N__28792));
    InMux I__6230 (
            .O(N__28795),
            .I(N__28789));
    Span4Mux_v I__6229 (
            .O(N__28792),
            .I(N__28784));
    LocalMux I__6228 (
            .O(N__28789),
            .I(N__28784));
    Span4Mux_h I__6227 (
            .O(N__28784),
            .I(N__28781));
    Span4Mux_s0_h I__6226 (
            .O(N__28781),
            .I(N__28778));
    Odrv4 I__6225 (
            .O(N__28778),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    InMux I__6224 (
            .O(N__28775),
            .I(N__28772));
    LocalMux I__6223 (
            .O(N__28772),
            .I(N__28769));
    Span4Mux_v I__6222 (
            .O(N__28769),
            .I(N__28766));
    Span4Mux_v I__6221 (
            .O(N__28766),
            .I(N__28763));
    Odrv4 I__6220 (
            .O(N__28763),
            .I(\VPP_VDDQ.un9_clk_100khz_2 ));
    InMux I__6219 (
            .O(N__28760),
            .I(N__28757));
    LocalMux I__6218 (
            .O(N__28757),
            .I(\VPP_VDDQ.un9_clk_100khz_0 ));
    CascadeMux I__6217 (
            .O(N__28754),
            .I(\VPP_VDDQ.un9_clk_100khz_1_cascade_ ));
    InMux I__6216 (
            .O(N__28751),
            .I(N__28748));
    LocalMux I__6215 (
            .O(N__28748),
            .I(\VPP_VDDQ.un9_clk_100khz_3 ));
    CascadeMux I__6214 (
            .O(N__28745),
            .I(N__28742));
    InMux I__6213 (
            .O(N__28742),
            .I(N__28739));
    LocalMux I__6212 (
            .O(N__28739),
            .I(\POWERLED.count_clk_0_10 ));
    InMux I__6211 (
            .O(N__28736),
            .I(N__28730));
    InMux I__6210 (
            .O(N__28735),
            .I(N__28730));
    LocalMux I__6209 (
            .O(N__28730),
            .I(N__28727));
    Odrv4 I__6208 (
            .O(N__28727),
            .I(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ));
    CascadeMux I__6207 (
            .O(N__28724),
            .I(N__28721));
    InMux I__6206 (
            .O(N__28721),
            .I(N__28718));
    LocalMux I__6205 (
            .O(N__28718),
            .I(N__28715));
    Odrv4 I__6204 (
            .O(N__28715),
            .I(\POWERLED.count_clkZ0Z_10 ));
    CascadeMux I__6203 (
            .O(N__28712),
            .I(\POWERLED.count_clkZ0Z_10_cascade_ ));
    InMux I__6202 (
            .O(N__28709),
            .I(N__28705));
    InMux I__6201 (
            .O(N__28708),
            .I(N__28702));
    LocalMux I__6200 (
            .O(N__28705),
            .I(N__28699));
    LocalMux I__6199 (
            .O(N__28702),
            .I(\POWERLED.count_clkZ0Z_15 ));
    Odrv4 I__6198 (
            .O(N__28699),
            .I(\POWERLED.count_clkZ0Z_15 ));
    InMux I__6197 (
            .O(N__28694),
            .I(N__28690));
    CascadeMux I__6196 (
            .O(N__28693),
            .I(N__28687));
    LocalMux I__6195 (
            .O(N__28690),
            .I(N__28684));
    InMux I__6194 (
            .O(N__28687),
            .I(N__28681));
    Odrv4 I__6193 (
            .O(N__28684),
            .I(\POWERLED.count_clkZ0Z_13 ));
    LocalMux I__6192 (
            .O(N__28681),
            .I(\POWERLED.count_clkZ0Z_13 ));
    CascadeMux I__6191 (
            .O(N__28676),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_4_cascade_ ));
    InMux I__6190 (
            .O(N__28673),
            .I(N__28669));
    CascadeMux I__6189 (
            .O(N__28672),
            .I(N__28666));
    LocalMux I__6188 (
            .O(N__28669),
            .I(N__28663));
    InMux I__6187 (
            .O(N__28666),
            .I(N__28660));
    Odrv4 I__6186 (
            .O(N__28663),
            .I(\POWERLED.count_clkZ0Z_14 ));
    LocalMux I__6185 (
            .O(N__28660),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__6184 (
            .O(N__28655),
            .I(N__28652));
    LocalMux I__6183 (
            .O(N__28652),
            .I(\POWERLED.count_clk_0_0 ));
    CascadeMux I__6182 (
            .O(N__28649),
            .I(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ));
    CascadeMux I__6181 (
            .O(N__28646),
            .I(\POWERLED.count_clkZ0Z_0_cascade_ ));
    CascadeMux I__6180 (
            .O(N__28643),
            .I(\POWERLED.N_352_cascade_ ));
    InMux I__6179 (
            .O(N__28640),
            .I(N__28637));
    LocalMux I__6178 (
            .O(N__28637),
            .I(N__28634));
    Span4Mux_h I__6177 (
            .O(N__28634),
            .I(N__28629));
    InMux I__6176 (
            .O(N__28633),
            .I(N__28626));
    InMux I__6175 (
            .O(N__28632),
            .I(N__28623));
    Odrv4 I__6174 (
            .O(N__28629),
            .I(\POWERLED.N_394 ));
    LocalMux I__6173 (
            .O(N__28626),
            .I(\POWERLED.N_394 ));
    LocalMux I__6172 (
            .O(N__28623),
            .I(\POWERLED.N_394 ));
    InMux I__6171 (
            .O(N__28616),
            .I(N__28610));
    InMux I__6170 (
            .O(N__28615),
            .I(N__28610));
    LocalMux I__6169 (
            .O(N__28610),
            .I(N__28606));
    CascadeMux I__6168 (
            .O(N__28609),
            .I(N__28603));
    Span4Mux_s3_h I__6167 (
            .O(N__28606),
            .I(N__28600));
    InMux I__6166 (
            .O(N__28603),
            .I(N__28597));
    Odrv4 I__6165 (
            .O(N__28600),
            .I(\POWERLED.count_clkZ0Z_2 ));
    LocalMux I__6164 (
            .O(N__28597),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__6163 (
            .O(N__28592),
            .I(N__28586));
    InMux I__6162 (
            .O(N__28591),
            .I(N__28586));
    LocalMux I__6161 (
            .O(N__28586),
            .I(N__28582));
    CascadeMux I__6160 (
            .O(N__28585),
            .I(N__28579));
    Span4Mux_s3_h I__6159 (
            .O(N__28582),
            .I(N__28576));
    InMux I__6158 (
            .O(N__28579),
            .I(N__28573));
    Odrv4 I__6157 (
            .O(N__28576),
            .I(\POWERLED.count_clkZ0Z_3 ));
    LocalMux I__6156 (
            .O(N__28573),
            .I(\POWERLED.count_clkZ0Z_3 ));
    CascadeMux I__6155 (
            .O(N__28568),
            .I(N__28565));
    InMux I__6154 (
            .O(N__28565),
            .I(N__28562));
    LocalMux I__6153 (
            .O(N__28562),
            .I(N__28557));
    InMux I__6152 (
            .O(N__28561),
            .I(N__28554));
    CascadeMux I__6151 (
            .O(N__28560),
            .I(N__28551));
    Span4Mux_s2_h I__6150 (
            .O(N__28557),
            .I(N__28548));
    LocalMux I__6149 (
            .O(N__28554),
            .I(N__28545));
    InMux I__6148 (
            .O(N__28551),
            .I(N__28542));
    Odrv4 I__6147 (
            .O(N__28548),
            .I(\POWERLED.count_clkZ0Z_6 ));
    Odrv4 I__6146 (
            .O(N__28545),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__6145 (
            .O(N__28542),
            .I(\POWERLED.count_clkZ0Z_6 ));
    InMux I__6144 (
            .O(N__28535),
            .I(N__28529));
    InMux I__6143 (
            .O(N__28534),
            .I(N__28529));
    LocalMux I__6142 (
            .O(N__28529),
            .I(N__28525));
    CascadeMux I__6141 (
            .O(N__28528),
            .I(N__28522));
    Span4Mux_v I__6140 (
            .O(N__28525),
            .I(N__28519));
    InMux I__6139 (
            .O(N__28522),
            .I(N__28516));
    Odrv4 I__6138 (
            .O(N__28519),
            .I(\POWERLED.count_clkZ0Z_8 ));
    LocalMux I__6137 (
            .O(N__28516),
            .I(\POWERLED.count_clkZ0Z_8 ));
    InMux I__6136 (
            .O(N__28511),
            .I(N__28507));
    InMux I__6135 (
            .O(N__28510),
            .I(N__28504));
    LocalMux I__6134 (
            .O(N__28507),
            .I(N__28500));
    LocalMux I__6133 (
            .O(N__28504),
            .I(N__28497));
    CascadeMux I__6132 (
            .O(N__28503),
            .I(N__28494));
    Span4Mux_h I__6131 (
            .O(N__28500),
            .I(N__28491));
    Span4Mux_s3_h I__6130 (
            .O(N__28497),
            .I(N__28488));
    InMux I__6129 (
            .O(N__28494),
            .I(N__28485));
    Odrv4 I__6128 (
            .O(N__28491),
            .I(\POWERLED.count_clkZ0Z_4 ));
    Odrv4 I__6127 (
            .O(N__28488),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__6126 (
            .O(N__28485),
            .I(\POWERLED.count_clkZ0Z_4 ));
    CascadeMux I__6125 (
            .O(N__28478),
            .I(\POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ));
    CascadeMux I__6124 (
            .O(N__28475),
            .I(N__28467));
    CascadeMux I__6123 (
            .O(N__28474),
            .I(N__28463));
    InMux I__6122 (
            .O(N__28473),
            .I(N__28457));
    InMux I__6121 (
            .O(N__28472),
            .I(N__28453));
    InMux I__6120 (
            .O(N__28471),
            .I(N__28450));
    InMux I__6119 (
            .O(N__28470),
            .I(N__28439));
    InMux I__6118 (
            .O(N__28467),
            .I(N__28439));
    InMux I__6117 (
            .O(N__28466),
            .I(N__28439));
    InMux I__6116 (
            .O(N__28463),
            .I(N__28436));
    CascadeMux I__6115 (
            .O(N__28462),
            .I(N__28433));
    CascadeMux I__6114 (
            .O(N__28461),
            .I(N__28430));
    InMux I__6113 (
            .O(N__28460),
            .I(N__28425));
    LocalMux I__6112 (
            .O(N__28457),
            .I(N__28421));
    InMux I__6111 (
            .O(N__28456),
            .I(N__28418));
    LocalMux I__6110 (
            .O(N__28453),
            .I(N__28415));
    LocalMux I__6109 (
            .O(N__28450),
            .I(N__28412));
    InMux I__6108 (
            .O(N__28449),
            .I(N__28409));
    InMux I__6107 (
            .O(N__28448),
            .I(N__28404));
    InMux I__6106 (
            .O(N__28447),
            .I(N__28404));
    InMux I__6105 (
            .O(N__28446),
            .I(N__28401));
    LocalMux I__6104 (
            .O(N__28439),
            .I(N__28398));
    LocalMux I__6103 (
            .O(N__28436),
            .I(N__28395));
    InMux I__6102 (
            .O(N__28433),
            .I(N__28388));
    InMux I__6101 (
            .O(N__28430),
            .I(N__28388));
    InMux I__6100 (
            .O(N__28429),
            .I(N__28388));
    InMux I__6099 (
            .O(N__28428),
            .I(N__28385));
    LocalMux I__6098 (
            .O(N__28425),
            .I(N__28382));
    InMux I__6097 (
            .O(N__28424),
            .I(N__28379));
    Span4Mux_h I__6096 (
            .O(N__28421),
            .I(N__28368));
    LocalMux I__6095 (
            .O(N__28418),
            .I(N__28368));
    Span4Mux_h I__6094 (
            .O(N__28415),
            .I(N__28368));
    Span4Mux_v I__6093 (
            .O(N__28412),
            .I(N__28368));
    LocalMux I__6092 (
            .O(N__28409),
            .I(N__28368));
    LocalMux I__6091 (
            .O(N__28404),
            .I(N__28365));
    LocalMux I__6090 (
            .O(N__28401),
            .I(N__28360));
    Span4Mux_s2_v I__6089 (
            .O(N__28398),
            .I(N__28360));
    Span4Mux_v I__6088 (
            .O(N__28395),
            .I(N__28349));
    LocalMux I__6087 (
            .O(N__28388),
            .I(N__28349));
    LocalMux I__6086 (
            .O(N__28385),
            .I(N__28349));
    Span4Mux_v I__6085 (
            .O(N__28382),
            .I(N__28349));
    LocalMux I__6084 (
            .O(N__28379),
            .I(N__28349));
    Span4Mux_v I__6083 (
            .O(N__28368),
            .I(N__28346));
    Span4Mux_h I__6082 (
            .O(N__28365),
            .I(N__28341));
    Span4Mux_h I__6081 (
            .O(N__28360),
            .I(N__28341));
    Span4Mux_v I__6080 (
            .O(N__28349),
            .I(N__28337));
    Span4Mux_h I__6079 (
            .O(N__28346),
            .I(N__28332));
    Span4Mux_v I__6078 (
            .O(N__28341),
            .I(N__28332));
    InMux I__6077 (
            .O(N__28340),
            .I(N__28329));
    Odrv4 I__6076 (
            .O(N__28337),
            .I(\POWERLED.N_2182_i ));
    Odrv4 I__6075 (
            .O(N__28332),
            .I(\POWERLED.N_2182_i ));
    LocalMux I__6074 (
            .O(N__28329),
            .I(\POWERLED.N_2182_i ));
    InMux I__6073 (
            .O(N__28322),
            .I(N__28319));
    LocalMux I__6072 (
            .O(N__28319),
            .I(\POWERLED.N_352 ));
    InMux I__6071 (
            .O(N__28316),
            .I(N__28306));
    InMux I__6070 (
            .O(N__28315),
            .I(N__28306));
    InMux I__6069 (
            .O(N__28314),
            .I(N__28306));
    CascadeMux I__6068 (
            .O(N__28313),
            .I(N__28303));
    LocalMux I__6067 (
            .O(N__28306),
            .I(N__28300));
    InMux I__6066 (
            .O(N__28303),
            .I(N__28297));
    Span4Mux_s2_h I__6065 (
            .O(N__28300),
            .I(N__28294));
    LocalMux I__6064 (
            .O(N__28297),
            .I(N__28291));
    Odrv4 I__6063 (
            .O(N__28294),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__6062 (
            .O(N__28291),
            .I(\POWERLED.count_clkZ0Z_7 ));
    CascadeMux I__6061 (
            .O(N__28286),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_2_2_cascade_ ));
    InMux I__6060 (
            .O(N__28283),
            .I(N__28274));
    InMux I__6059 (
            .O(N__28282),
            .I(N__28274));
    InMux I__6058 (
            .O(N__28281),
            .I(N__28274));
    LocalMux I__6057 (
            .O(N__28274),
            .I(\POWERLED.count_clk_RNIZ0Z_9 ));
    InMux I__6056 (
            .O(N__28271),
            .I(N__28265));
    InMux I__6055 (
            .O(N__28270),
            .I(N__28265));
    LocalMux I__6054 (
            .O(N__28265),
            .I(\POWERLED.count_offZ0Z_6 ));
    InMux I__6053 (
            .O(N__28262),
            .I(N__28259));
    LocalMux I__6052 (
            .O(N__28259),
            .I(N__28256));
    Span4Mux_v I__6051 (
            .O(N__28256),
            .I(N__28253));
    Odrv4 I__6050 (
            .O(N__28253),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a3_0 ));
    CascadeMux I__6049 (
            .O(N__28250),
            .I(N__28246));
    InMux I__6048 (
            .O(N__28249),
            .I(N__28243));
    InMux I__6047 (
            .O(N__28246),
            .I(N__28238));
    LocalMux I__6046 (
            .O(N__28243),
            .I(N__28235));
    InMux I__6045 (
            .O(N__28242),
            .I(N__28232));
    InMux I__6044 (
            .O(N__28241),
            .I(N__28229));
    LocalMux I__6043 (
            .O(N__28238),
            .I(N__28226));
    Span4Mux_h I__6042 (
            .O(N__28235),
            .I(N__28221));
    LocalMux I__6041 (
            .O(N__28232),
            .I(N__28221));
    LocalMux I__6040 (
            .O(N__28229),
            .I(N__28218));
    Odrv4 I__6039 (
            .O(N__28226),
            .I(\POWERLED.func_state_RNI_2Z0Z_1 ));
    Odrv4 I__6038 (
            .O(N__28221),
            .I(\POWERLED.func_state_RNI_2Z0Z_1 ));
    Odrv12 I__6037 (
            .O(N__28218),
            .I(\POWERLED.func_state_RNI_2Z0Z_1 ));
    CascadeMux I__6036 (
            .O(N__28211),
            .I(\POWERLED.N_289_cascade_ ));
    InMux I__6035 (
            .O(N__28208),
            .I(N__28204));
    InMux I__6034 (
            .O(N__28207),
            .I(N__28201));
    LocalMux I__6033 (
            .O(N__28204),
            .I(N__28197));
    LocalMux I__6032 (
            .O(N__28201),
            .I(N__28194));
    InMux I__6031 (
            .O(N__28200),
            .I(N__28191));
    Span4Mux_v I__6030 (
            .O(N__28197),
            .I(N__28188));
    Span4Mux_v I__6029 (
            .O(N__28194),
            .I(N__28185));
    LocalMux I__6028 (
            .O(N__28191),
            .I(\POWERLED.func_state_RNIBVNS_2Z0Z_0 ));
    Odrv4 I__6027 (
            .O(N__28188),
            .I(\POWERLED.func_state_RNIBVNS_2Z0Z_0 ));
    Odrv4 I__6026 (
            .O(N__28185),
            .I(\POWERLED.func_state_RNIBVNS_2Z0Z_0 ));
    InMux I__6025 (
            .O(N__28178),
            .I(N__28174));
    InMux I__6024 (
            .O(N__28177),
            .I(N__28171));
    LocalMux I__6023 (
            .O(N__28174),
            .I(N__28167));
    LocalMux I__6022 (
            .O(N__28171),
            .I(N__28164));
    InMux I__6021 (
            .O(N__28170),
            .I(N__28161));
    Span4Mux_v I__6020 (
            .O(N__28167),
            .I(N__28153));
    Span4Mux_h I__6019 (
            .O(N__28164),
            .I(N__28148));
    LocalMux I__6018 (
            .O(N__28161),
            .I(N__28148));
    InMux I__6017 (
            .O(N__28160),
            .I(N__28145));
    InMux I__6016 (
            .O(N__28159),
            .I(N__28140));
    InMux I__6015 (
            .O(N__28158),
            .I(N__28140));
    InMux I__6014 (
            .O(N__28157),
            .I(N__28135));
    InMux I__6013 (
            .O(N__28156),
            .I(N__28135));
    Odrv4 I__6012 (
            .O(N__28153),
            .I(\POWERLED.count_off_RNIG5N6N1Z0Z_11 ));
    Odrv4 I__6011 (
            .O(N__28148),
            .I(\POWERLED.count_off_RNIG5N6N1Z0Z_11 ));
    LocalMux I__6010 (
            .O(N__28145),
            .I(\POWERLED.count_off_RNIG5N6N1Z0Z_11 ));
    LocalMux I__6009 (
            .O(N__28140),
            .I(\POWERLED.count_off_RNIG5N6N1Z0Z_11 ));
    LocalMux I__6008 (
            .O(N__28135),
            .I(\POWERLED.count_off_RNIG5N6N1Z0Z_11 ));
    CascadeMux I__6007 (
            .O(N__28124),
            .I(N__28121));
    InMux I__6006 (
            .O(N__28121),
            .I(N__28117));
    InMux I__6005 (
            .O(N__28120),
            .I(N__28114));
    LocalMux I__6004 (
            .O(N__28117),
            .I(N__28111));
    LocalMux I__6003 (
            .O(N__28114),
            .I(N__28108));
    Span4Mux_h I__6002 (
            .O(N__28111),
            .I(N__28105));
    Odrv4 I__6001 (
            .O(N__28108),
            .I(\POWERLED.func_state_RNI_5Z0Z_1 ));
    Odrv4 I__6000 (
            .O(N__28105),
            .I(\POWERLED.func_state_RNI_5Z0Z_1 ));
    CascadeMux I__5999 (
            .O(N__28100),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_2_tz_0_cascade_ ));
    InMux I__5998 (
            .O(N__28097),
            .I(N__28094));
    LocalMux I__5997 (
            .O(N__28094),
            .I(N__28091));
    Odrv12 I__5996 (
            .O(N__28091),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_2 ));
    InMux I__5995 (
            .O(N__28088),
            .I(N__28084));
    InMux I__5994 (
            .O(N__28087),
            .I(N__28081));
    LocalMux I__5993 (
            .O(N__28084),
            .I(N__28076));
    LocalMux I__5992 (
            .O(N__28081),
            .I(N__28076));
    Odrv4 I__5991 (
            .O(N__28076),
            .I(\POWERLED.func_state_RNI_2Z0Z_0 ));
    CascadeMux I__5990 (
            .O(N__28073),
            .I(N__28069));
    InMux I__5989 (
            .O(N__28072),
            .I(N__28060));
    InMux I__5988 (
            .O(N__28069),
            .I(N__28060));
    InMux I__5987 (
            .O(N__28068),
            .I(N__28057));
    CascadeMux I__5986 (
            .O(N__28067),
            .I(N__28049));
    InMux I__5985 (
            .O(N__28066),
            .I(N__28045));
    InMux I__5984 (
            .O(N__28065),
            .I(N__28042));
    LocalMux I__5983 (
            .O(N__28060),
            .I(N__28038));
    LocalMux I__5982 (
            .O(N__28057),
            .I(N__28035));
    InMux I__5981 (
            .O(N__28056),
            .I(N__28032));
    InMux I__5980 (
            .O(N__28055),
            .I(N__28024));
    InMux I__5979 (
            .O(N__28054),
            .I(N__28021));
    InMux I__5978 (
            .O(N__28053),
            .I(N__28018));
    InMux I__5977 (
            .O(N__28052),
            .I(N__28015));
    InMux I__5976 (
            .O(N__28049),
            .I(N__28010));
    InMux I__5975 (
            .O(N__28048),
            .I(N__28010));
    LocalMux I__5974 (
            .O(N__28045),
            .I(N__28005));
    LocalMux I__5973 (
            .O(N__28042),
            .I(N__28005));
    CascadeMux I__5972 (
            .O(N__28041),
            .I(N__28002));
    Span4Mux_v I__5971 (
            .O(N__28038),
            .I(N__27996));
    Span4Mux_v I__5970 (
            .O(N__28035),
            .I(N__27996));
    LocalMux I__5969 (
            .O(N__28032),
            .I(N__27993));
    InMux I__5968 (
            .O(N__28031),
            .I(N__27990));
    InMux I__5967 (
            .O(N__28030),
            .I(N__27983));
    InMux I__5966 (
            .O(N__28029),
            .I(N__27983));
    InMux I__5965 (
            .O(N__28028),
            .I(N__27983));
    InMux I__5964 (
            .O(N__28027),
            .I(N__27980));
    LocalMux I__5963 (
            .O(N__28024),
            .I(N__27976));
    LocalMux I__5962 (
            .O(N__28021),
            .I(N__27973));
    LocalMux I__5961 (
            .O(N__28018),
            .I(N__27970));
    LocalMux I__5960 (
            .O(N__28015),
            .I(N__27965));
    LocalMux I__5959 (
            .O(N__28010),
            .I(N__27965));
    Span4Mux_v I__5958 (
            .O(N__28005),
            .I(N__27962));
    InMux I__5957 (
            .O(N__28002),
            .I(N__27957));
    InMux I__5956 (
            .O(N__28001),
            .I(N__27957));
    Span4Mux_v I__5955 (
            .O(N__27996),
            .I(N__27952));
    Span4Mux_v I__5954 (
            .O(N__27993),
            .I(N__27952));
    LocalMux I__5953 (
            .O(N__27990),
            .I(N__27949));
    LocalMux I__5952 (
            .O(N__27983),
            .I(N__27946));
    LocalMux I__5951 (
            .O(N__27980),
            .I(N__27943));
    InMux I__5950 (
            .O(N__27979),
            .I(N__27940));
    Span4Mux_v I__5949 (
            .O(N__27976),
            .I(N__27931));
    Span4Mux_s3_v I__5948 (
            .O(N__27973),
            .I(N__27931));
    Span4Mux_s3_v I__5947 (
            .O(N__27970),
            .I(N__27931));
    Span4Mux_v I__5946 (
            .O(N__27965),
            .I(N__27931));
    Span4Mux_h I__5945 (
            .O(N__27962),
            .I(N__27926));
    LocalMux I__5944 (
            .O(N__27957),
            .I(N__27926));
    Span4Mux_h I__5943 (
            .O(N__27952),
            .I(N__27919));
    Span4Mux_h I__5942 (
            .O(N__27949),
            .I(N__27919));
    Span4Mux_s3_v I__5941 (
            .O(N__27946),
            .I(N__27919));
    Span12Mux_s3_v I__5940 (
            .O(N__27943),
            .I(N__27914));
    LocalMux I__5939 (
            .O(N__27940),
            .I(N__27914));
    Span4Mux_h I__5938 (
            .O(N__27931),
            .I(N__27909));
    Span4Mux_v I__5937 (
            .O(N__27926),
            .I(N__27909));
    Odrv4 I__5936 (
            .O(N__27919),
            .I(gpio_fpga_soc_4));
    Odrv12 I__5935 (
            .O(N__27914),
            .I(gpio_fpga_soc_4));
    Odrv4 I__5934 (
            .O(N__27909),
            .I(gpio_fpga_soc_4));
    InMux I__5933 (
            .O(N__27902),
            .I(N__27899));
    LocalMux I__5932 (
            .O(N__27899),
            .I(N__27896));
    Span4Mux_h I__5931 (
            .O(N__27896),
            .I(N__27893));
    Odrv4 I__5930 (
            .O(N__27893),
            .I(\POWERLED.un1_func_state25_6_0_o_N_304_N ));
    InMux I__5929 (
            .O(N__27890),
            .I(N__27886));
    CascadeMux I__5928 (
            .O(N__27889),
            .I(N__27877));
    LocalMux I__5927 (
            .O(N__27886),
            .I(N__27873));
    InMux I__5926 (
            .O(N__27885),
            .I(N__27870));
    CascadeMux I__5925 (
            .O(N__27884),
            .I(N__27867));
    InMux I__5924 (
            .O(N__27883),
            .I(N__27860));
    InMux I__5923 (
            .O(N__27882),
            .I(N__27860));
    InMux I__5922 (
            .O(N__27881),
            .I(N__27860));
    CascadeMux I__5921 (
            .O(N__27880),
            .I(N__27856));
    InMux I__5920 (
            .O(N__27877),
            .I(N__27853));
    InMux I__5919 (
            .O(N__27876),
            .I(N__27850));
    Sp12to4 I__5918 (
            .O(N__27873),
            .I(N__27845));
    LocalMux I__5917 (
            .O(N__27870),
            .I(N__27845));
    InMux I__5916 (
            .O(N__27867),
            .I(N__27842));
    LocalMux I__5915 (
            .O(N__27860),
            .I(N__27839));
    InMux I__5914 (
            .O(N__27859),
            .I(N__27836));
    InMux I__5913 (
            .O(N__27856),
            .I(N__27832));
    LocalMux I__5912 (
            .O(N__27853),
            .I(N__27827));
    LocalMux I__5911 (
            .O(N__27850),
            .I(N__27827));
    Span12Mux_s11_v I__5910 (
            .O(N__27845),
            .I(N__27824));
    LocalMux I__5909 (
            .O(N__27842),
            .I(N__27819));
    Span4Mux_s3_h I__5908 (
            .O(N__27839),
            .I(N__27819));
    LocalMux I__5907 (
            .O(N__27836),
            .I(N__27816));
    InMux I__5906 (
            .O(N__27835),
            .I(N__27813));
    LocalMux I__5905 (
            .O(N__27832),
            .I(\POWERLED.un1_N_3_mux_0 ));
    Odrv4 I__5904 (
            .O(N__27827),
            .I(\POWERLED.un1_N_3_mux_0 ));
    Odrv12 I__5903 (
            .O(N__27824),
            .I(\POWERLED.un1_N_3_mux_0 ));
    Odrv4 I__5902 (
            .O(N__27819),
            .I(\POWERLED.un1_N_3_mux_0 ));
    Odrv12 I__5901 (
            .O(N__27816),
            .I(\POWERLED.un1_N_3_mux_0 ));
    LocalMux I__5900 (
            .O(N__27813),
            .I(\POWERLED.un1_N_3_mux_0 ));
    InMux I__5899 (
            .O(N__27800),
            .I(N__27791));
    CascadeMux I__5898 (
            .O(N__27799),
            .I(N__27788));
    InMux I__5897 (
            .O(N__27798),
            .I(N__27783));
    InMux I__5896 (
            .O(N__27797),
            .I(N__27783));
    InMux I__5895 (
            .O(N__27796),
            .I(N__27780));
    InMux I__5894 (
            .O(N__27795),
            .I(N__27772));
    InMux I__5893 (
            .O(N__27794),
            .I(N__27769));
    LocalMux I__5892 (
            .O(N__27791),
            .I(N__27764));
    InMux I__5891 (
            .O(N__27788),
            .I(N__27761));
    LocalMux I__5890 (
            .O(N__27783),
            .I(N__27756));
    LocalMux I__5889 (
            .O(N__27780),
            .I(N__27756));
    InMux I__5888 (
            .O(N__27779),
            .I(N__27749));
    InMux I__5887 (
            .O(N__27778),
            .I(N__27749));
    InMux I__5886 (
            .O(N__27777),
            .I(N__27749));
    InMux I__5885 (
            .O(N__27776),
            .I(N__27744));
    InMux I__5884 (
            .O(N__27775),
            .I(N__27744));
    LocalMux I__5883 (
            .O(N__27772),
            .I(N__27741));
    LocalMux I__5882 (
            .O(N__27769),
            .I(N__27729));
    InMux I__5881 (
            .O(N__27768),
            .I(N__27726));
    InMux I__5880 (
            .O(N__27767),
            .I(N__27723));
    Span4Mux_v I__5879 (
            .O(N__27764),
            .I(N__27720));
    LocalMux I__5878 (
            .O(N__27761),
            .I(N__27717));
    Span4Mux_v I__5877 (
            .O(N__27756),
            .I(N__27714));
    LocalMux I__5876 (
            .O(N__27749),
            .I(N__27709));
    LocalMux I__5875 (
            .O(N__27744),
            .I(N__27709));
    Span4Mux_v I__5874 (
            .O(N__27741),
            .I(N__27706));
    InMux I__5873 (
            .O(N__27740),
            .I(N__27703));
    InMux I__5872 (
            .O(N__27739),
            .I(N__27694));
    InMux I__5871 (
            .O(N__27738),
            .I(N__27694));
    InMux I__5870 (
            .O(N__27737),
            .I(N__27694));
    InMux I__5869 (
            .O(N__27736),
            .I(N__27694));
    InMux I__5868 (
            .O(N__27735),
            .I(N__27685));
    InMux I__5867 (
            .O(N__27734),
            .I(N__27685));
    InMux I__5866 (
            .O(N__27733),
            .I(N__27685));
    InMux I__5865 (
            .O(N__27732),
            .I(N__27685));
    Span4Mux_v I__5864 (
            .O(N__27729),
            .I(N__27678));
    LocalMux I__5863 (
            .O(N__27726),
            .I(N__27678));
    LocalMux I__5862 (
            .O(N__27723),
            .I(N__27678));
    Odrv4 I__5861 (
            .O(N__27720),
            .I(\POWERLED.func_state ));
    Odrv12 I__5860 (
            .O(N__27717),
            .I(\POWERLED.func_state ));
    Odrv4 I__5859 (
            .O(N__27714),
            .I(\POWERLED.func_state ));
    Odrv4 I__5858 (
            .O(N__27709),
            .I(\POWERLED.func_state ));
    Odrv4 I__5857 (
            .O(N__27706),
            .I(\POWERLED.func_state ));
    LocalMux I__5856 (
            .O(N__27703),
            .I(\POWERLED.func_state ));
    LocalMux I__5855 (
            .O(N__27694),
            .I(\POWERLED.func_state ));
    LocalMux I__5854 (
            .O(N__27685),
            .I(\POWERLED.func_state ));
    Odrv4 I__5853 (
            .O(N__27678),
            .I(\POWERLED.func_state ));
    InMux I__5852 (
            .O(N__27659),
            .I(N__27656));
    LocalMux I__5851 (
            .O(N__27656),
            .I(N__27653));
    Odrv4 I__5850 (
            .O(N__27653),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_2_0 ));
    CascadeMux I__5849 (
            .O(N__27650),
            .I(N__27647));
    InMux I__5848 (
            .O(N__27647),
            .I(N__27644));
    LocalMux I__5847 (
            .O(N__27644),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_3_0 ));
    InMux I__5846 (
            .O(N__27641),
            .I(N__27638));
    LocalMux I__5845 (
            .O(N__27638),
            .I(\POWERLED.count_off_1_2 ));
    CascadeMux I__5844 (
            .O(N__27635),
            .I(\POWERLED.count_off_1_2_cascade_ ));
    InMux I__5843 (
            .O(N__27632),
            .I(N__27626));
    InMux I__5842 (
            .O(N__27631),
            .I(N__27626));
    LocalMux I__5841 (
            .O(N__27626),
            .I(\POWERLED.count_offZ0Z_2 ));
    InMux I__5840 (
            .O(N__27623),
            .I(N__27620));
    LocalMux I__5839 (
            .O(N__27620),
            .I(\POWERLED.count_off_1_7 ));
    CascadeMux I__5838 (
            .O(N__27617),
            .I(\POWERLED.count_off_1_7_cascade_ ));
    InMux I__5837 (
            .O(N__27614),
            .I(N__27611));
    LocalMux I__5836 (
            .O(N__27611),
            .I(\POWERLED.un34_clk_100khz_3 ));
    InMux I__5835 (
            .O(N__27608),
            .I(N__27602));
    InMux I__5834 (
            .O(N__27607),
            .I(N__27602));
    LocalMux I__5833 (
            .O(N__27602),
            .I(\POWERLED.count_offZ0Z_7 ));
    InMux I__5832 (
            .O(N__27599),
            .I(N__27596));
    LocalMux I__5831 (
            .O(N__27596),
            .I(N__27593));
    Span4Mux_v I__5830 (
            .O(N__27593),
            .I(N__27590));
    Odrv4 I__5829 (
            .O(N__27590),
            .I(\POWERLED.count_off_1_11 ));
    CascadeMux I__5828 (
            .O(N__27587),
            .I(\POWERLED.count_off_1_11_cascade_ ));
    CascadeMux I__5827 (
            .O(N__27584),
            .I(N__27581));
    InMux I__5826 (
            .O(N__27581),
            .I(N__27578));
    LocalMux I__5825 (
            .O(N__27578),
            .I(N__27575));
    Span4Mux_v I__5824 (
            .O(N__27575),
            .I(N__27571));
    InMux I__5823 (
            .O(N__27574),
            .I(N__27568));
    Odrv4 I__5822 (
            .O(N__27571),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__5821 (
            .O(N__27568),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__5820 (
            .O(N__27563),
            .I(N__27560));
    LocalMux I__5819 (
            .O(N__27560),
            .I(\POWERLED.count_off_0_15 ));
    InMux I__5818 (
            .O(N__27557),
            .I(N__27554));
    LocalMux I__5817 (
            .O(N__27554),
            .I(\POWERLED.count_off_0_8 ));
    CascadeMux I__5816 (
            .O(N__27551),
            .I(\POWERLED.un34_clk_100khz_0_cascade_ ));
    InMux I__5815 (
            .O(N__27548),
            .I(N__27545));
    LocalMux I__5814 (
            .O(N__27545),
            .I(N__27542));
    Odrv12 I__5813 (
            .O(N__27542),
            .I(\POWERLED.un34_clk_100khz_12 ));
    InMux I__5812 (
            .O(N__27539),
            .I(N__27536));
    LocalMux I__5811 (
            .O(N__27536),
            .I(\POWERLED.un34_clk_100khz_1 ));
    InMux I__5810 (
            .O(N__27533),
            .I(N__27530));
    LocalMux I__5809 (
            .O(N__27530),
            .I(\POWERLED.count_off_1_6 ));
    CascadeMux I__5808 (
            .O(N__27527),
            .I(\POWERLED.count_off_1_6_cascade_ ));
    InMux I__5807 (
            .O(N__27524),
            .I(N__27520));
    InMux I__5806 (
            .O(N__27523),
            .I(N__27517));
    LocalMux I__5805 (
            .O(N__27520),
            .I(N__27514));
    LocalMux I__5804 (
            .O(N__27517),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    Odrv4 I__5803 (
            .O(N__27514),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__5802 (
            .O(N__27509),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    InMux I__5801 (
            .O(N__27506),
            .I(N__27502));
    InMux I__5800 (
            .O(N__27505),
            .I(N__27499));
    LocalMux I__5799 (
            .O(N__27502),
            .I(N__27496));
    LocalMux I__5798 (
            .O(N__27499),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    Odrv4 I__5797 (
            .O(N__27496),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    InMux I__5796 (
            .O(N__27491),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__5795 (
            .O(N__27488),
            .I(N__27484));
    InMux I__5794 (
            .O(N__27487),
            .I(N__27481));
    LocalMux I__5793 (
            .O(N__27484),
            .I(N__27478));
    LocalMux I__5792 (
            .O(N__27481),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    Odrv4 I__5791 (
            .O(N__27478),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__5790 (
            .O(N__27473),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    InMux I__5789 (
            .O(N__27470),
            .I(N__27465));
    InMux I__5788 (
            .O(N__27469),
            .I(N__27462));
    InMux I__5787 (
            .O(N__27468),
            .I(N__27457));
    LocalMux I__5786 (
            .O(N__27465),
            .I(N__27454));
    LocalMux I__5785 (
            .O(N__27462),
            .I(N__27450));
    InMux I__5784 (
            .O(N__27461),
            .I(N__27446));
    IoInMux I__5783 (
            .O(N__27460),
            .I(N__27442));
    LocalMux I__5782 (
            .O(N__27457),
            .I(N__27439));
    Span4Mux_s1_h I__5781 (
            .O(N__27454),
            .I(N__27436));
    InMux I__5780 (
            .O(N__27453),
            .I(N__27433));
    Span4Mux_v I__5779 (
            .O(N__27450),
            .I(N__27430));
    InMux I__5778 (
            .O(N__27449),
            .I(N__27427));
    LocalMux I__5777 (
            .O(N__27446),
            .I(N__27424));
    InMux I__5776 (
            .O(N__27445),
            .I(N__27421));
    LocalMux I__5775 (
            .O(N__27442),
            .I(N__27418));
    Span4Mux_v I__5774 (
            .O(N__27439),
            .I(N__27415));
    Span4Mux_h I__5773 (
            .O(N__27436),
            .I(N__27410));
    LocalMux I__5772 (
            .O(N__27433),
            .I(N__27410));
    Span4Mux_h I__5771 (
            .O(N__27430),
            .I(N__27405));
    LocalMux I__5770 (
            .O(N__27427),
            .I(N__27405));
    Span4Mux_v I__5769 (
            .O(N__27424),
            .I(N__27400));
    LocalMux I__5768 (
            .O(N__27421),
            .I(N__27400));
    Span4Mux_s3_h I__5767 (
            .O(N__27418),
            .I(N__27397));
    Span4Mux_v I__5766 (
            .O(N__27415),
            .I(N__27392));
    Span4Mux_v I__5765 (
            .O(N__27410),
            .I(N__27392));
    Span4Mux_v I__5764 (
            .O(N__27405),
            .I(N__27387));
    Span4Mux_h I__5763 (
            .O(N__27400),
            .I(N__27387));
    Odrv4 I__5762 (
            .O(N__27397),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5761 (
            .O(N__27392),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5760 (
            .O(N__27387),
            .I(CONSTANT_ONE_NET));
    InMux I__5759 (
            .O(N__27380),
            .I(bfn_9_15_0_));
    CascadeMux I__5758 (
            .O(N__27377),
            .I(N__27374));
    InMux I__5757 (
            .O(N__27374),
            .I(N__27370));
    InMux I__5756 (
            .O(N__27373),
            .I(N__27367));
    LocalMux I__5755 (
            .O(N__27370),
            .I(N__27364));
    LocalMux I__5754 (
            .O(N__27367),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    Odrv12 I__5753 (
            .O(N__27364),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    CascadeMux I__5752 (
            .O(N__27359),
            .I(N__27356));
    InMux I__5751 (
            .O(N__27356),
            .I(N__27353));
    LocalMux I__5750 (
            .O(N__27353),
            .I(\POWERLED.count_off_0_5 ));
    InMux I__5749 (
            .O(N__27350),
            .I(N__27346));
    InMux I__5748 (
            .O(N__27349),
            .I(N__27343));
    LocalMux I__5747 (
            .O(N__27346),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__5746 (
            .O(N__27343),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__5745 (
            .O(N__27338),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    InMux I__5744 (
            .O(N__27335),
            .I(N__27331));
    InMux I__5743 (
            .O(N__27334),
            .I(N__27328));
    LocalMux I__5742 (
            .O(N__27331),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__5741 (
            .O(N__27328),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    InMux I__5740 (
            .O(N__27323),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__5739 (
            .O(N__27320),
            .I(N__27316));
    InMux I__5738 (
            .O(N__27319),
            .I(N__27313));
    LocalMux I__5737 (
            .O(N__27316),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__5736 (
            .O(N__27313),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__5735 (
            .O(N__27308),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__5734 (
            .O(N__27305),
            .I(N__27301));
    InMux I__5733 (
            .O(N__27304),
            .I(N__27298));
    LocalMux I__5732 (
            .O(N__27301),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    LocalMux I__5731 (
            .O(N__27298),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__5730 (
            .O(N__27293),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    CascadeMux I__5729 (
            .O(N__27290),
            .I(N__27286));
    InMux I__5728 (
            .O(N__27289),
            .I(N__27283));
    InMux I__5727 (
            .O(N__27286),
            .I(N__27280));
    LocalMux I__5726 (
            .O(N__27283),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__5725 (
            .O(N__27280),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__5724 (
            .O(N__27275),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__5723 (
            .O(N__27272),
            .I(N__27268));
    InMux I__5722 (
            .O(N__27271),
            .I(N__27265));
    LocalMux I__5721 (
            .O(N__27268),
            .I(N__27262));
    LocalMux I__5720 (
            .O(N__27265),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    Odrv4 I__5719 (
            .O(N__27262),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__5718 (
            .O(N__27257),
            .I(bfn_9_14_0_));
    InMux I__5717 (
            .O(N__27254),
            .I(N__27250));
    InMux I__5716 (
            .O(N__27253),
            .I(N__27247));
    LocalMux I__5715 (
            .O(N__27250),
            .I(N__27244));
    LocalMux I__5714 (
            .O(N__27247),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    Odrv4 I__5713 (
            .O(N__27244),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__5712 (
            .O(N__27239),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    CascadeMux I__5711 (
            .O(N__27236),
            .I(N__27233));
    InMux I__5710 (
            .O(N__27233),
            .I(N__27229));
    InMux I__5709 (
            .O(N__27232),
            .I(N__27226));
    LocalMux I__5708 (
            .O(N__27229),
            .I(N__27223));
    LocalMux I__5707 (
            .O(N__27226),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    Odrv4 I__5706 (
            .O(N__27223),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__5705 (
            .O(N__27218),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    CascadeMux I__5704 (
            .O(N__27215),
            .I(N__27212));
    InMux I__5703 (
            .O(N__27212),
            .I(N__27208));
    InMux I__5702 (
            .O(N__27211),
            .I(N__27205));
    LocalMux I__5701 (
            .O(N__27208),
            .I(N__27202));
    LocalMux I__5700 (
            .O(N__27205),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    Odrv4 I__5699 (
            .O(N__27202),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__5698 (
            .O(N__27197),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    CascadeMux I__5697 (
            .O(N__27194),
            .I(N__27191));
    InMux I__5696 (
            .O(N__27191),
            .I(N__27188));
    LocalMux I__5695 (
            .O(N__27188),
            .I(N__27185));
    Odrv12 I__5694 (
            .O(N__27185),
            .I(\POWERLED.dutycycle_RNIZ0Z_1 ));
    InMux I__5693 (
            .O(N__27182),
            .I(N__27179));
    LocalMux I__5692 (
            .O(N__27179),
            .I(\VPP_VDDQ.un6_count_10 ));
    CascadeMux I__5691 (
            .O(N__27176),
            .I(\VPP_VDDQ.un6_count_8_cascade_ ));
    InMux I__5690 (
            .O(N__27173),
            .I(N__27170));
    LocalMux I__5689 (
            .O(N__27170),
            .I(\VPP_VDDQ.un6_count_11 ));
    InMux I__5688 (
            .O(N__27167),
            .I(N__27164));
    LocalMux I__5687 (
            .O(N__27164),
            .I(\VPP_VDDQ.un6_count_9 ));
    InMux I__5686 (
            .O(N__27161),
            .I(N__27157));
    InMux I__5685 (
            .O(N__27160),
            .I(N__27154));
    LocalMux I__5684 (
            .O(N__27157),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__5683 (
            .O(N__27154),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    InMux I__5682 (
            .O(N__27149),
            .I(N__27145));
    InMux I__5681 (
            .O(N__27148),
            .I(N__27142));
    LocalMux I__5680 (
            .O(N__27145),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__5679 (
            .O(N__27142),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__5678 (
            .O(N__27137),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__5677 (
            .O(N__27134),
            .I(N__27130));
    InMux I__5676 (
            .O(N__27133),
            .I(N__27127));
    LocalMux I__5675 (
            .O(N__27130),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__5674 (
            .O(N__27127),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    InMux I__5673 (
            .O(N__27122),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    InMux I__5672 (
            .O(N__27119),
            .I(N__27116));
    LocalMux I__5671 (
            .O(N__27116),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_0 ));
    InMux I__5670 (
            .O(N__27113),
            .I(N__27110));
    LocalMux I__5669 (
            .O(N__27110),
            .I(\POWERLED.un1_dutycycle_172_m3 ));
    InMux I__5668 (
            .O(N__27107),
            .I(N__27099));
    InMux I__5667 (
            .O(N__27106),
            .I(N__27094));
    InMux I__5666 (
            .O(N__27105),
            .I(N__27089));
    InMux I__5665 (
            .O(N__27104),
            .I(N__27086));
    InMux I__5664 (
            .O(N__27103),
            .I(N__27081));
    InMux I__5663 (
            .O(N__27102),
            .I(N__27081));
    LocalMux I__5662 (
            .O(N__27099),
            .I(N__27078));
    CascadeMux I__5661 (
            .O(N__27098),
            .I(N__27074));
    InMux I__5660 (
            .O(N__27097),
            .I(N__27071));
    LocalMux I__5659 (
            .O(N__27094),
            .I(N__27068));
    InMux I__5658 (
            .O(N__27093),
            .I(N__27065));
    InMux I__5657 (
            .O(N__27092),
            .I(N__27062));
    LocalMux I__5656 (
            .O(N__27089),
            .I(N__27055));
    LocalMux I__5655 (
            .O(N__27086),
            .I(N__27055));
    LocalMux I__5654 (
            .O(N__27081),
            .I(N__27055));
    Span4Mux_v I__5653 (
            .O(N__27078),
            .I(N__27049));
    InMux I__5652 (
            .O(N__27077),
            .I(N__27046));
    InMux I__5651 (
            .O(N__27074),
            .I(N__27043));
    LocalMux I__5650 (
            .O(N__27071),
            .I(N__27039));
    Span4Mux_v I__5649 (
            .O(N__27068),
            .I(N__27030));
    LocalMux I__5648 (
            .O(N__27065),
            .I(N__27030));
    LocalMux I__5647 (
            .O(N__27062),
            .I(N__27030));
    Span4Mux_v I__5646 (
            .O(N__27055),
            .I(N__27030));
    CascadeMux I__5645 (
            .O(N__27054),
            .I(N__27026));
    CascadeMux I__5644 (
            .O(N__27053),
            .I(N__27014));
    CascadeMux I__5643 (
            .O(N__27052),
            .I(N__27010));
    Span4Mux_v I__5642 (
            .O(N__27049),
            .I(N__27005));
    LocalMux I__5641 (
            .O(N__27046),
            .I(N__27005));
    LocalMux I__5640 (
            .O(N__27043),
            .I(N__27002));
    InMux I__5639 (
            .O(N__27042),
            .I(N__26999));
    Span4Mux_h I__5638 (
            .O(N__27039),
            .I(N__26994));
    Span4Mux_v I__5637 (
            .O(N__27030),
            .I(N__26994));
    InMux I__5636 (
            .O(N__27029),
            .I(N__26985));
    InMux I__5635 (
            .O(N__27026),
            .I(N__26985));
    InMux I__5634 (
            .O(N__27025),
            .I(N__26985));
    InMux I__5633 (
            .O(N__27024),
            .I(N__26985));
    InMux I__5632 (
            .O(N__27023),
            .I(N__26976));
    InMux I__5631 (
            .O(N__27022),
            .I(N__26976));
    InMux I__5630 (
            .O(N__27021),
            .I(N__26976));
    InMux I__5629 (
            .O(N__27020),
            .I(N__26976));
    InMux I__5628 (
            .O(N__27019),
            .I(N__26963));
    InMux I__5627 (
            .O(N__27018),
            .I(N__26963));
    InMux I__5626 (
            .O(N__27017),
            .I(N__26963));
    InMux I__5625 (
            .O(N__27014),
            .I(N__26963));
    InMux I__5624 (
            .O(N__27013),
            .I(N__26963));
    InMux I__5623 (
            .O(N__27010),
            .I(N__26963));
    Odrv4 I__5622 (
            .O(N__27005),
            .I(\POWERLED.N_2200_i ));
    Odrv4 I__5621 (
            .O(N__27002),
            .I(\POWERLED.N_2200_i ));
    LocalMux I__5620 (
            .O(N__26999),
            .I(\POWERLED.N_2200_i ));
    Odrv4 I__5619 (
            .O(N__26994),
            .I(\POWERLED.N_2200_i ));
    LocalMux I__5618 (
            .O(N__26985),
            .I(\POWERLED.N_2200_i ));
    LocalMux I__5617 (
            .O(N__26976),
            .I(\POWERLED.N_2200_i ));
    LocalMux I__5616 (
            .O(N__26963),
            .I(\POWERLED.N_2200_i ));
    InMux I__5615 (
            .O(N__26948),
            .I(N__26945));
    LocalMux I__5614 (
            .O(N__26945),
            .I(\POWERLED.un1_dutycycle_96_0_a3_1 ));
    CascadeMux I__5613 (
            .O(N__26942),
            .I(N__26934));
    CascadeMux I__5612 (
            .O(N__26941),
            .I(N__26929));
    InMux I__5611 (
            .O(N__26940),
            .I(N__26924));
    InMux I__5610 (
            .O(N__26939),
            .I(N__26924));
    InMux I__5609 (
            .O(N__26938),
            .I(N__26918));
    InMux I__5608 (
            .O(N__26937),
            .I(N__26913));
    InMux I__5607 (
            .O(N__26934),
            .I(N__26913));
    InMux I__5606 (
            .O(N__26933),
            .I(N__26910));
    InMux I__5605 (
            .O(N__26932),
            .I(N__26907));
    InMux I__5604 (
            .O(N__26929),
            .I(N__26904));
    LocalMux I__5603 (
            .O(N__26924),
            .I(N__26901));
    InMux I__5602 (
            .O(N__26923),
            .I(N__26894));
    InMux I__5601 (
            .O(N__26922),
            .I(N__26894));
    InMux I__5600 (
            .O(N__26921),
            .I(N__26894));
    LocalMux I__5599 (
            .O(N__26918),
            .I(N__26891));
    LocalMux I__5598 (
            .O(N__26913),
            .I(N__26888));
    LocalMux I__5597 (
            .O(N__26910),
            .I(N__26885));
    LocalMux I__5596 (
            .O(N__26907),
            .I(N__26879));
    LocalMux I__5595 (
            .O(N__26904),
            .I(N__26879));
    Span4Mux_h I__5594 (
            .O(N__26901),
            .I(N__26870));
    LocalMux I__5593 (
            .O(N__26894),
            .I(N__26870));
    Span4Mux_v I__5592 (
            .O(N__26891),
            .I(N__26870));
    Span4Mux_h I__5591 (
            .O(N__26888),
            .I(N__26870));
    Span4Mux_h I__5590 (
            .O(N__26885),
            .I(N__26867));
    InMux I__5589 (
            .O(N__26884),
            .I(N__26864));
    Span4Mux_v I__5588 (
            .O(N__26879),
            .I(N__26859));
    Span4Mux_v I__5587 (
            .O(N__26870),
            .I(N__26859));
    Odrv4 I__5586 (
            .O(N__26867),
            .I(\POWERLED.dutycycle ));
    LocalMux I__5585 (
            .O(N__26864),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__5584 (
            .O(N__26859),
            .I(\POWERLED.dutycycle ));
    InMux I__5583 (
            .O(N__26852),
            .I(N__26848));
    InMux I__5582 (
            .O(N__26851),
            .I(N__26845));
    LocalMux I__5581 (
            .O(N__26848),
            .I(\POWERLED.N_327 ));
    LocalMux I__5580 (
            .O(N__26845),
            .I(\POWERLED.N_327 ));
    InMux I__5579 (
            .O(N__26840),
            .I(N__26837));
    LocalMux I__5578 (
            .O(N__26837),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_0 ));
    InMux I__5577 (
            .O(N__26834),
            .I(N__26828));
    InMux I__5576 (
            .O(N__26833),
            .I(N__26823));
    InMux I__5575 (
            .O(N__26832),
            .I(N__26823));
    InMux I__5574 (
            .O(N__26831),
            .I(N__26820));
    LocalMux I__5573 (
            .O(N__26828),
            .I(N__26817));
    LocalMux I__5572 (
            .O(N__26823),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_5 ));
    LocalMux I__5571 (
            .O(N__26820),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_5 ));
    Odrv4 I__5570 (
            .O(N__26817),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_5 ));
    CascadeMux I__5569 (
            .O(N__26810),
            .I(\POWERLED.un1_dutycycle_53_axb_3_1_0_cascade_ ));
    CascadeMux I__5568 (
            .O(N__26807),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_1_cascade_ ));
    InMux I__5567 (
            .O(N__26804),
            .I(N__26801));
    LocalMux I__5566 (
            .O(N__26801),
            .I(N__26798));
    Odrv12 I__5565 (
            .O(N__26798),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_2 ));
    InMux I__5564 (
            .O(N__26795),
            .I(N__26792));
    LocalMux I__5563 (
            .O(N__26792),
            .I(N__26789));
    Span4Mux_v I__5562 (
            .O(N__26789),
            .I(N__26785));
    InMux I__5561 (
            .O(N__26788),
            .I(N__26782));
    Odrv4 I__5560 (
            .O(N__26785),
            .I(\POWERLED.N_342 ));
    LocalMux I__5559 (
            .O(N__26782),
            .I(\POWERLED.N_342 ));
    InMux I__5558 (
            .O(N__26777),
            .I(N__26774));
    LocalMux I__5557 (
            .O(N__26774),
            .I(N__26771));
    Span4Mux_v I__5556 (
            .O(N__26771),
            .I(N__26766));
    InMux I__5555 (
            .O(N__26770),
            .I(N__26763));
    InMux I__5554 (
            .O(N__26769),
            .I(N__26760));
    Span4Mux_h I__5553 (
            .O(N__26766),
            .I(N__26755));
    LocalMux I__5552 (
            .O(N__26763),
            .I(N__26755));
    LocalMux I__5551 (
            .O(N__26760),
            .I(\POWERLED.N_155 ));
    Odrv4 I__5550 (
            .O(N__26755),
            .I(\POWERLED.N_155 ));
    CascadeMux I__5549 (
            .O(N__26750),
            .I(N__26746));
    InMux I__5548 (
            .O(N__26749),
            .I(N__26743));
    InMux I__5547 (
            .O(N__26746),
            .I(N__26740));
    LocalMux I__5546 (
            .O(N__26743),
            .I(N__26736));
    LocalMux I__5545 (
            .O(N__26740),
            .I(N__26733));
    InMux I__5544 (
            .O(N__26739),
            .I(N__26730));
    Span4Mux_s3_h I__5543 (
            .O(N__26736),
            .I(N__26727));
    Span4Mux_v I__5542 (
            .O(N__26733),
            .I(N__26724));
    LocalMux I__5541 (
            .O(N__26730),
            .I(N__26721));
    Span4Mux_h I__5540 (
            .O(N__26727),
            .I(N__26718));
    Odrv4 I__5539 (
            .O(N__26724),
            .I(\POWERLED.N_336 ));
    Odrv4 I__5538 (
            .O(N__26721),
            .I(\POWERLED.N_336 ));
    Odrv4 I__5537 (
            .O(N__26718),
            .I(\POWERLED.N_336 ));
    InMux I__5536 (
            .O(N__26711),
            .I(N__26708));
    LocalMux I__5535 (
            .O(N__26708),
            .I(N__26704));
    InMux I__5534 (
            .O(N__26707),
            .I(N__26701));
    Odrv4 I__5533 (
            .O(N__26704),
            .I(\POWERLED.dutycycle_RNI_9Z0Z_0 ));
    LocalMux I__5532 (
            .O(N__26701),
            .I(\POWERLED.dutycycle_RNI_9Z0Z_0 ));
    CascadeMux I__5531 (
            .O(N__26696),
            .I(N__26689));
    InMux I__5530 (
            .O(N__26695),
            .I(N__26686));
    InMux I__5529 (
            .O(N__26694),
            .I(N__26683));
    CascadeMux I__5528 (
            .O(N__26693),
            .I(N__26678));
    CascadeMux I__5527 (
            .O(N__26692),
            .I(N__26672));
    InMux I__5526 (
            .O(N__26689),
            .I(N__26669));
    LocalMux I__5525 (
            .O(N__26686),
            .I(N__26666));
    LocalMux I__5524 (
            .O(N__26683),
            .I(N__26663));
    InMux I__5523 (
            .O(N__26682),
            .I(N__26660));
    InMux I__5522 (
            .O(N__26681),
            .I(N__26655));
    InMux I__5521 (
            .O(N__26678),
            .I(N__26655));
    InMux I__5520 (
            .O(N__26677),
            .I(N__26652));
    InMux I__5519 (
            .O(N__26676),
            .I(N__26647));
    InMux I__5518 (
            .O(N__26675),
            .I(N__26647));
    InMux I__5517 (
            .O(N__26672),
            .I(N__26644));
    LocalMux I__5516 (
            .O(N__26669),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv12 I__5515 (
            .O(N__26666),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv12 I__5514 (
            .O(N__26663),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__5513 (
            .O(N__26660),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__5512 (
            .O(N__26655),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__5511 (
            .O(N__26652),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__5510 (
            .O(N__26647),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__5509 (
            .O(N__26644),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    CascadeMux I__5508 (
            .O(N__26627),
            .I(N__26623));
    InMux I__5507 (
            .O(N__26626),
            .I(N__26619));
    InMux I__5506 (
            .O(N__26623),
            .I(N__26614));
    InMux I__5505 (
            .O(N__26622),
            .I(N__26614));
    LocalMux I__5504 (
            .O(N__26619),
            .I(N__26608));
    LocalMux I__5503 (
            .O(N__26614),
            .I(N__26608));
    InMux I__5502 (
            .O(N__26613),
            .I(N__26603));
    Span4Mux_v I__5501 (
            .O(N__26608),
            .I(N__26596));
    InMux I__5500 (
            .O(N__26607),
            .I(N__26591));
    InMux I__5499 (
            .O(N__26606),
            .I(N__26591));
    LocalMux I__5498 (
            .O(N__26603),
            .I(N__26588));
    InMux I__5497 (
            .O(N__26602),
            .I(N__26579));
    InMux I__5496 (
            .O(N__26601),
            .I(N__26579));
    InMux I__5495 (
            .O(N__26600),
            .I(N__26579));
    InMux I__5494 (
            .O(N__26599),
            .I(N__26579));
    Span4Mux_h I__5493 (
            .O(N__26596),
            .I(N__26569));
    LocalMux I__5492 (
            .O(N__26591),
            .I(N__26569));
    Span4Mux_h I__5491 (
            .O(N__26588),
            .I(N__26559));
    LocalMux I__5490 (
            .O(N__26579),
            .I(N__26559));
    InMux I__5489 (
            .O(N__26578),
            .I(N__26556));
    InMux I__5488 (
            .O(N__26577),
            .I(N__26551));
    InMux I__5487 (
            .O(N__26576),
            .I(N__26548));
    InMux I__5486 (
            .O(N__26575),
            .I(N__26543));
    InMux I__5485 (
            .O(N__26574),
            .I(N__26543));
    Span4Mux_h I__5484 (
            .O(N__26569),
            .I(N__26540));
    InMux I__5483 (
            .O(N__26568),
            .I(N__26529));
    InMux I__5482 (
            .O(N__26567),
            .I(N__26529));
    InMux I__5481 (
            .O(N__26566),
            .I(N__26529));
    InMux I__5480 (
            .O(N__26565),
            .I(N__26529));
    InMux I__5479 (
            .O(N__26564),
            .I(N__26529));
    Sp12to4 I__5478 (
            .O(N__26559),
            .I(N__26524));
    LocalMux I__5477 (
            .O(N__26556),
            .I(N__26524));
    InMux I__5476 (
            .O(N__26555),
            .I(N__26519));
    InMux I__5475 (
            .O(N__26554),
            .I(N__26519));
    LocalMux I__5474 (
            .O(N__26551),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__5473 (
            .O(N__26548),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__5472 (
            .O(N__26543),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__5471 (
            .O(N__26540),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__5470 (
            .O(N__26529),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv12 I__5469 (
            .O(N__26524),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__5468 (
            .O(N__26519),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    InMux I__5467 (
            .O(N__26504),
            .I(N__26501));
    LocalMux I__5466 (
            .O(N__26501),
            .I(N__26498));
    Span4Mux_h I__5465 (
            .O(N__26498),
            .I(N__26495));
    Odrv4 I__5464 (
            .O(N__26495),
            .I(\POWERLED.un1_i3_mux ));
    CascadeMux I__5463 (
            .O(N__26492),
            .I(N__26484));
    InMux I__5462 (
            .O(N__26491),
            .I(N__26479));
    InMux I__5461 (
            .O(N__26490),
            .I(N__26476));
    InMux I__5460 (
            .O(N__26489),
            .I(N__26472));
    InMux I__5459 (
            .O(N__26488),
            .I(N__26463));
    InMux I__5458 (
            .O(N__26487),
            .I(N__26463));
    InMux I__5457 (
            .O(N__26484),
            .I(N__26463));
    InMux I__5456 (
            .O(N__26483),
            .I(N__26463));
    CascadeMux I__5455 (
            .O(N__26482),
            .I(N__26459));
    LocalMux I__5454 (
            .O(N__26479),
            .I(N__26452));
    LocalMux I__5453 (
            .O(N__26476),
            .I(N__26449));
    InMux I__5452 (
            .O(N__26475),
            .I(N__26446));
    LocalMux I__5451 (
            .O(N__26472),
            .I(N__26441));
    LocalMux I__5450 (
            .O(N__26463),
            .I(N__26441));
    InMux I__5449 (
            .O(N__26462),
            .I(N__26438));
    InMux I__5448 (
            .O(N__26459),
            .I(N__26435));
    InMux I__5447 (
            .O(N__26458),
            .I(N__26426));
    InMux I__5446 (
            .O(N__26457),
            .I(N__26426));
    InMux I__5445 (
            .O(N__26456),
            .I(N__26426));
    InMux I__5444 (
            .O(N__26455),
            .I(N__26426));
    Span4Mux_v I__5443 (
            .O(N__26452),
            .I(N__26417));
    Span4Mux_h I__5442 (
            .O(N__26449),
            .I(N__26417));
    LocalMux I__5441 (
            .O(N__26446),
            .I(N__26417));
    Span4Mux_v I__5440 (
            .O(N__26441),
            .I(N__26417));
    LocalMux I__5439 (
            .O(N__26438),
            .I(N__26412));
    LocalMux I__5438 (
            .O(N__26435),
            .I(N__26412));
    LocalMux I__5437 (
            .O(N__26426),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__5436 (
            .O(N__26417),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__5435 (
            .O(N__26412),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    CascadeMux I__5434 (
            .O(N__26405),
            .I(N__26402));
    InMux I__5433 (
            .O(N__26402),
            .I(N__26398));
    CascadeMux I__5432 (
            .O(N__26401),
            .I(N__26384));
    LocalMux I__5431 (
            .O(N__26398),
            .I(N__26377));
    InMux I__5430 (
            .O(N__26397),
            .I(N__26372));
    InMux I__5429 (
            .O(N__26396),
            .I(N__26372));
    InMux I__5428 (
            .O(N__26395),
            .I(N__26367));
    InMux I__5427 (
            .O(N__26394),
            .I(N__26367));
    InMux I__5426 (
            .O(N__26393),
            .I(N__26364));
    InMux I__5425 (
            .O(N__26392),
            .I(N__26359));
    InMux I__5424 (
            .O(N__26391),
            .I(N__26359));
    InMux I__5423 (
            .O(N__26390),
            .I(N__26354));
    InMux I__5422 (
            .O(N__26389),
            .I(N__26347));
    InMux I__5421 (
            .O(N__26388),
            .I(N__26347));
    InMux I__5420 (
            .O(N__26387),
            .I(N__26347));
    InMux I__5419 (
            .O(N__26384),
            .I(N__26344));
    InMux I__5418 (
            .O(N__26383),
            .I(N__26335));
    InMux I__5417 (
            .O(N__26382),
            .I(N__26335));
    InMux I__5416 (
            .O(N__26381),
            .I(N__26335));
    InMux I__5415 (
            .O(N__26380),
            .I(N__26335));
    Span4Mux_h I__5414 (
            .O(N__26377),
            .I(N__26332));
    LocalMux I__5413 (
            .O(N__26372),
            .I(N__26325));
    LocalMux I__5412 (
            .O(N__26367),
            .I(N__26325));
    LocalMux I__5411 (
            .O(N__26364),
            .I(N__26325));
    LocalMux I__5410 (
            .O(N__26359),
            .I(N__26322));
    CascadeMux I__5409 (
            .O(N__26358),
            .I(N__26319));
    InMux I__5408 (
            .O(N__26357),
            .I(N__26316));
    LocalMux I__5407 (
            .O(N__26354),
            .I(N__26311));
    LocalMux I__5406 (
            .O(N__26347),
            .I(N__26311));
    LocalMux I__5405 (
            .O(N__26344),
            .I(N__26300));
    LocalMux I__5404 (
            .O(N__26335),
            .I(N__26300));
    Span4Mux_s1_v I__5403 (
            .O(N__26332),
            .I(N__26300));
    Span4Mux_h I__5402 (
            .O(N__26325),
            .I(N__26300));
    Span4Mux_h I__5401 (
            .O(N__26322),
            .I(N__26300));
    InMux I__5400 (
            .O(N__26319),
            .I(N__26297));
    LocalMux I__5399 (
            .O(N__26316),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__5398 (
            .O(N__26311),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__5397 (
            .O(N__26300),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__5396 (
            .O(N__26297),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    CascadeMux I__5395 (
            .O(N__26288),
            .I(N__26283));
    CascadeMux I__5394 (
            .O(N__26287),
            .I(N__26279));
    CascadeMux I__5393 (
            .O(N__26286),
            .I(N__26275));
    InMux I__5392 (
            .O(N__26283),
            .I(N__26270));
    InMux I__5391 (
            .O(N__26282),
            .I(N__26267));
    InMux I__5390 (
            .O(N__26279),
            .I(N__26260));
    InMux I__5389 (
            .O(N__26278),
            .I(N__26260));
    InMux I__5388 (
            .O(N__26275),
            .I(N__26253));
    InMux I__5387 (
            .O(N__26274),
            .I(N__26253));
    InMux I__5386 (
            .O(N__26273),
            .I(N__26253));
    LocalMux I__5385 (
            .O(N__26270),
            .I(N__26248));
    LocalMux I__5384 (
            .O(N__26267),
            .I(N__26248));
    InMux I__5383 (
            .O(N__26266),
            .I(N__26245));
    InMux I__5382 (
            .O(N__26265),
            .I(N__26242));
    LocalMux I__5381 (
            .O(N__26260),
            .I(N__26237));
    LocalMux I__5380 (
            .O(N__26253),
            .I(N__26234));
    Span4Mux_h I__5379 (
            .O(N__26248),
            .I(N__26229));
    LocalMux I__5378 (
            .O(N__26245),
            .I(N__26229));
    LocalMux I__5377 (
            .O(N__26242),
            .I(N__26226));
    CascadeMux I__5376 (
            .O(N__26241),
            .I(N__26223));
    InMux I__5375 (
            .O(N__26240),
            .I(N__26220));
    Span4Mux_h I__5374 (
            .O(N__26237),
            .I(N__26215));
    Span4Mux_h I__5373 (
            .O(N__26234),
            .I(N__26215));
    Span4Mux_h I__5372 (
            .O(N__26229),
            .I(N__26210));
    Span4Mux_v I__5371 (
            .O(N__26226),
            .I(N__26210));
    InMux I__5370 (
            .O(N__26223),
            .I(N__26207));
    LocalMux I__5369 (
            .O(N__26220),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__5368 (
            .O(N__26215),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__5367 (
            .O(N__26210),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__5366 (
            .O(N__26207),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    CascadeMux I__5365 (
            .O(N__26198),
            .I(N__26195));
    InMux I__5364 (
            .O(N__26195),
            .I(N__26185));
    InMux I__5363 (
            .O(N__26194),
            .I(N__26185));
    CascadeMux I__5362 (
            .O(N__26193),
            .I(N__26181));
    CascadeMux I__5361 (
            .O(N__26192),
            .I(N__26178));
    CascadeMux I__5360 (
            .O(N__26191),
            .I(N__26175));
    CascadeMux I__5359 (
            .O(N__26190),
            .I(N__26172));
    LocalMux I__5358 (
            .O(N__26185),
            .I(N__26167));
    CascadeMux I__5357 (
            .O(N__26184),
            .I(N__26162));
    InMux I__5356 (
            .O(N__26181),
            .I(N__26157));
    InMux I__5355 (
            .O(N__26178),
            .I(N__26157));
    InMux I__5354 (
            .O(N__26175),
            .I(N__26154));
    InMux I__5353 (
            .O(N__26172),
            .I(N__26150));
    InMux I__5352 (
            .O(N__26171),
            .I(N__26145));
    InMux I__5351 (
            .O(N__26170),
            .I(N__26145));
    Span4Mux_h I__5350 (
            .O(N__26167),
            .I(N__26142));
    InMux I__5349 (
            .O(N__26166),
            .I(N__26139));
    InMux I__5348 (
            .O(N__26165),
            .I(N__26136));
    InMux I__5347 (
            .O(N__26162),
            .I(N__26133));
    LocalMux I__5346 (
            .O(N__26157),
            .I(N__26128));
    LocalMux I__5345 (
            .O(N__26154),
            .I(N__26128));
    InMux I__5344 (
            .O(N__26153),
            .I(N__26125));
    LocalMux I__5343 (
            .O(N__26150),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5342 (
            .O(N__26145),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__5341 (
            .O(N__26142),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5340 (
            .O(N__26139),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5339 (
            .O(N__26136),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5338 (
            .O(N__26133),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__5337 (
            .O(N__26128),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5336 (
            .O(N__26125),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    InMux I__5335 (
            .O(N__26108),
            .I(N__26105));
    LocalMux I__5334 (
            .O(N__26105),
            .I(N__26102));
    Span4Mux_h I__5333 (
            .O(N__26102),
            .I(N__26099));
    Span4Mux_v I__5332 (
            .O(N__26099),
            .I(N__26094));
    InMux I__5331 (
            .O(N__26098),
            .I(N__26091));
    InMux I__5330 (
            .O(N__26097),
            .I(N__26088));
    Odrv4 I__5329 (
            .O(N__26094),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    LocalMux I__5328 (
            .O(N__26091),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    LocalMux I__5327 (
            .O(N__26088),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    CascadeMux I__5326 (
            .O(N__26081),
            .I(N__26078));
    InMux I__5325 (
            .O(N__26078),
            .I(N__26075));
    LocalMux I__5324 (
            .O(N__26075),
            .I(N__26072));
    Span4Mux_h I__5323 (
            .O(N__26072),
            .I(N__26069));
    Span4Mux_v I__5322 (
            .O(N__26069),
            .I(N__26066));
    Odrv4 I__5321 (
            .O(N__26066),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    CascadeMux I__5320 (
            .O(N__26063),
            .I(N__26060));
    InMux I__5319 (
            .O(N__26060),
            .I(N__26057));
    LocalMux I__5318 (
            .O(N__26057),
            .I(N__26054));
    Span4Mux_v I__5317 (
            .O(N__26054),
            .I(N__26050));
    InMux I__5316 (
            .O(N__26053),
            .I(N__26047));
    Odrv4 I__5315 (
            .O(N__26050),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_0 ));
    LocalMux I__5314 (
            .O(N__26047),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_0 ));
    CascadeMux I__5313 (
            .O(N__26042),
            .I(\POWERLED.un1_dutycycle_172_m4_bm_rn_0_cascade_ ));
    InMux I__5312 (
            .O(N__26039),
            .I(N__26036));
    LocalMux I__5311 (
            .O(N__26036),
            .I(\POWERLED.dutycycle_RNIMUFP1Z0Z_2 ));
    InMux I__5310 (
            .O(N__26033),
            .I(N__26023));
    InMux I__5309 (
            .O(N__26032),
            .I(N__26020));
    InMux I__5308 (
            .O(N__26031),
            .I(N__26017));
    CascadeMux I__5307 (
            .O(N__26030),
            .I(N__26013));
    CascadeMux I__5306 (
            .O(N__26029),
            .I(N__26010));
    CascadeMux I__5305 (
            .O(N__26028),
            .I(N__26007));
    CascadeMux I__5304 (
            .O(N__26027),
            .I(N__26004));
    InMux I__5303 (
            .O(N__26026),
            .I(N__25997));
    LocalMux I__5302 (
            .O(N__26023),
            .I(N__25992));
    LocalMux I__5301 (
            .O(N__26020),
            .I(N__25992));
    LocalMux I__5300 (
            .O(N__26017),
            .I(N__25989));
    InMux I__5299 (
            .O(N__26016),
            .I(N__25986));
    InMux I__5298 (
            .O(N__26013),
            .I(N__25973));
    InMux I__5297 (
            .O(N__26010),
            .I(N__25973));
    InMux I__5296 (
            .O(N__26007),
            .I(N__25973));
    InMux I__5295 (
            .O(N__26004),
            .I(N__25973));
    InMux I__5294 (
            .O(N__26003),
            .I(N__25973));
    InMux I__5293 (
            .O(N__26002),
            .I(N__25973));
    InMux I__5292 (
            .O(N__26001),
            .I(N__25970));
    InMux I__5291 (
            .O(N__26000),
            .I(N__25967));
    LocalMux I__5290 (
            .O(N__25997),
            .I(N__25964));
    Span4Mux_s3_v I__5289 (
            .O(N__25992),
            .I(N__25961));
    Span4Mux_v I__5288 (
            .O(N__25989),
            .I(N__25956));
    LocalMux I__5287 (
            .O(N__25986),
            .I(N__25956));
    LocalMux I__5286 (
            .O(N__25973),
            .I(N__25953));
    LocalMux I__5285 (
            .O(N__25970),
            .I(N__25950));
    LocalMux I__5284 (
            .O(N__25967),
            .I(N__25947));
    Span4Mux_s3_h I__5283 (
            .O(N__25964),
            .I(N__25944));
    Span4Mux_h I__5282 (
            .O(N__25961),
            .I(N__25941));
    Span4Mux_h I__5281 (
            .O(N__25956),
            .I(N__25938));
    Span4Mux_h I__5280 (
            .O(N__25953),
            .I(N__25933));
    Span4Mux_h I__5279 (
            .O(N__25950),
            .I(N__25933));
    Odrv4 I__5278 (
            .O(N__25947),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__5277 (
            .O(N__25944),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__5276 (
            .O(N__25941),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__5275 (
            .O(N__25938),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__5274 (
            .O(N__25933),
            .I(COUNTER_un4_counter_7_THRU_CO));
    IoInMux I__5273 (
            .O(N__25922),
            .I(N__25919));
    LocalMux I__5272 (
            .O(N__25919),
            .I(N__25916));
    IoSpan4Mux I__5271 (
            .O(N__25916),
            .I(N__25913));
    Span4Mux_s3_v I__5270 (
            .O(N__25913),
            .I(N__25910));
    Odrv4 I__5269 (
            .O(N__25910),
            .I(G_9));
    InMux I__5268 (
            .O(N__25907),
            .I(N__25904));
    LocalMux I__5267 (
            .O(N__25904),
            .I(\POWERLED.un1_dutycycle_172_m4_bm_sn ));
    InMux I__5266 (
            .O(N__25901),
            .I(N__25895));
    InMux I__5265 (
            .O(N__25900),
            .I(N__25895));
    LocalMux I__5264 (
            .O(N__25895),
            .I(N__25892));
    Span4Mux_h I__5263 (
            .O(N__25892),
            .I(N__25886));
    InMux I__5262 (
            .O(N__25891),
            .I(N__25883));
    InMux I__5261 (
            .O(N__25890),
            .I(N__25878));
    InMux I__5260 (
            .O(N__25889),
            .I(N__25878));
    Odrv4 I__5259 (
            .O(N__25886),
            .I(\POWERLED.N_20_i ));
    LocalMux I__5258 (
            .O(N__25883),
            .I(\POWERLED.N_20_i ));
    LocalMux I__5257 (
            .O(N__25878),
            .I(\POWERLED.N_20_i ));
    CascadeMux I__5256 (
            .O(N__25871),
            .I(N__25866));
    InMux I__5255 (
            .O(N__25870),
            .I(N__25862));
    InMux I__5254 (
            .O(N__25869),
            .I(N__25855));
    InMux I__5253 (
            .O(N__25866),
            .I(N__25855));
    InMux I__5252 (
            .O(N__25865),
            .I(N__25855));
    LocalMux I__5251 (
            .O(N__25862),
            .I(N__25851));
    LocalMux I__5250 (
            .O(N__25855),
            .I(N__25848));
    InMux I__5249 (
            .O(N__25854),
            .I(N__25843));
    Span4Mux_v I__5248 (
            .O(N__25851),
            .I(N__25838));
    Span4Mux_h I__5247 (
            .O(N__25848),
            .I(N__25838));
    InMux I__5246 (
            .O(N__25847),
            .I(N__25833));
    InMux I__5245 (
            .O(N__25846),
            .I(N__25833));
    LocalMux I__5244 (
            .O(N__25843),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    Odrv4 I__5243 (
            .O(N__25838),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    LocalMux I__5242 (
            .O(N__25833),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    CascadeMux I__5241 (
            .O(N__25826),
            .I(\POWERLED.un1_count_off_1_sqmuxa_2_0_cascade_ ));
    CascadeMux I__5240 (
            .O(N__25823),
            .I(N__25806));
    InMux I__5239 (
            .O(N__25822),
            .I(N__25802));
    CascadeMux I__5238 (
            .O(N__25821),
            .I(N__25798));
    CascadeMux I__5237 (
            .O(N__25820),
            .I(N__25794));
    InMux I__5236 (
            .O(N__25819),
            .I(N__25788));
    InMux I__5235 (
            .O(N__25818),
            .I(N__25788));
    InMux I__5234 (
            .O(N__25817),
            .I(N__25783));
    InMux I__5233 (
            .O(N__25816),
            .I(N__25783));
    InMux I__5232 (
            .O(N__25815),
            .I(N__25775));
    InMux I__5231 (
            .O(N__25814),
            .I(N__25775));
    InMux I__5230 (
            .O(N__25813),
            .I(N__25775));
    InMux I__5229 (
            .O(N__25812),
            .I(N__25768));
    InMux I__5228 (
            .O(N__25811),
            .I(N__25768));
    InMux I__5227 (
            .O(N__25810),
            .I(N__25768));
    InMux I__5226 (
            .O(N__25809),
            .I(N__25763));
    InMux I__5225 (
            .O(N__25806),
            .I(N__25760));
    InMux I__5224 (
            .O(N__25805),
            .I(N__25753));
    LocalMux I__5223 (
            .O(N__25802),
            .I(N__25750));
    InMux I__5222 (
            .O(N__25801),
            .I(N__25747));
    InMux I__5221 (
            .O(N__25798),
            .I(N__25742));
    InMux I__5220 (
            .O(N__25797),
            .I(N__25742));
    InMux I__5219 (
            .O(N__25794),
            .I(N__25739));
    CascadeMux I__5218 (
            .O(N__25793),
            .I(N__25735));
    LocalMux I__5217 (
            .O(N__25788),
            .I(N__25729));
    LocalMux I__5216 (
            .O(N__25783),
            .I(N__25724));
    InMux I__5215 (
            .O(N__25782),
            .I(N__25719));
    LocalMux I__5214 (
            .O(N__25775),
            .I(N__25712));
    LocalMux I__5213 (
            .O(N__25768),
            .I(N__25712));
    InMux I__5212 (
            .O(N__25767),
            .I(N__25707));
    InMux I__5211 (
            .O(N__25766),
            .I(N__25707));
    LocalMux I__5210 (
            .O(N__25763),
            .I(N__25702));
    LocalMux I__5209 (
            .O(N__25760),
            .I(N__25702));
    InMux I__5208 (
            .O(N__25759),
            .I(N__25699));
    InMux I__5207 (
            .O(N__25758),
            .I(N__25696));
    InMux I__5206 (
            .O(N__25757),
            .I(N__25691));
    InMux I__5205 (
            .O(N__25756),
            .I(N__25691));
    LocalMux I__5204 (
            .O(N__25753),
            .I(N__25680));
    Span4Mux_s1_v I__5203 (
            .O(N__25750),
            .I(N__25680));
    LocalMux I__5202 (
            .O(N__25747),
            .I(N__25680));
    LocalMux I__5201 (
            .O(N__25742),
            .I(N__25680));
    LocalMux I__5200 (
            .O(N__25739),
            .I(N__25680));
    InMux I__5199 (
            .O(N__25738),
            .I(N__25677));
    InMux I__5198 (
            .O(N__25735),
            .I(N__25668));
    InMux I__5197 (
            .O(N__25734),
            .I(N__25668));
    InMux I__5196 (
            .O(N__25733),
            .I(N__25668));
    InMux I__5195 (
            .O(N__25732),
            .I(N__25668));
    Span4Mux_v I__5194 (
            .O(N__25729),
            .I(N__25665));
    InMux I__5193 (
            .O(N__25728),
            .I(N__25660));
    InMux I__5192 (
            .O(N__25727),
            .I(N__25660));
    Span4Mux_v I__5191 (
            .O(N__25724),
            .I(N__25657));
    InMux I__5190 (
            .O(N__25723),
            .I(N__25652));
    InMux I__5189 (
            .O(N__25722),
            .I(N__25652));
    LocalMux I__5188 (
            .O(N__25719),
            .I(N__25649));
    InMux I__5187 (
            .O(N__25718),
            .I(N__25644));
    InMux I__5186 (
            .O(N__25717),
            .I(N__25644));
    Span4Mux_v I__5185 (
            .O(N__25712),
            .I(N__25637));
    LocalMux I__5184 (
            .O(N__25707),
            .I(N__25637));
    Span4Mux_v I__5183 (
            .O(N__25702),
            .I(N__25637));
    LocalMux I__5182 (
            .O(N__25699),
            .I(N__25628));
    LocalMux I__5181 (
            .O(N__25696),
            .I(N__25628));
    LocalMux I__5180 (
            .O(N__25691),
            .I(N__25628));
    Span4Mux_v I__5179 (
            .O(N__25680),
            .I(N__25628));
    LocalMux I__5178 (
            .O(N__25677),
            .I(N__25623));
    LocalMux I__5177 (
            .O(N__25668),
            .I(N__25623));
    Odrv4 I__5176 (
            .O(N__25665),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    LocalMux I__5175 (
            .O(N__25660),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    Odrv4 I__5174 (
            .O(N__25657),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    LocalMux I__5173 (
            .O(N__25652),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    Odrv4 I__5172 (
            .O(N__25649),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    LocalMux I__5171 (
            .O(N__25644),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    Odrv4 I__5170 (
            .O(N__25637),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    Odrv4 I__5169 (
            .O(N__25628),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    Odrv12 I__5168 (
            .O(N__25623),
            .I(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ));
    InMux I__5167 (
            .O(N__25604),
            .I(N__25598));
    InMux I__5166 (
            .O(N__25603),
            .I(N__25598));
    LocalMux I__5165 (
            .O(N__25598),
            .I(N__25591));
    InMux I__5164 (
            .O(N__25597),
            .I(N__25588));
    CascadeMux I__5163 (
            .O(N__25596),
            .I(N__25585));
    InMux I__5162 (
            .O(N__25595),
            .I(N__25573));
    InMux I__5161 (
            .O(N__25594),
            .I(N__25573));
    Span4Mux_h I__5160 (
            .O(N__25591),
            .I(N__25568));
    LocalMux I__5159 (
            .O(N__25588),
            .I(N__25568));
    InMux I__5158 (
            .O(N__25585),
            .I(N__25563));
    InMux I__5157 (
            .O(N__25584),
            .I(N__25563));
    InMux I__5156 (
            .O(N__25583),
            .I(N__25556));
    InMux I__5155 (
            .O(N__25582),
            .I(N__25556));
    InMux I__5154 (
            .O(N__25581),
            .I(N__25556));
    InMux I__5153 (
            .O(N__25580),
            .I(N__25553));
    InMux I__5152 (
            .O(N__25579),
            .I(N__25548));
    InMux I__5151 (
            .O(N__25578),
            .I(N__25548));
    LocalMux I__5150 (
            .O(N__25573),
            .I(N__25541));
    Span4Mux_v I__5149 (
            .O(N__25568),
            .I(N__25541));
    LocalMux I__5148 (
            .O(N__25563),
            .I(N__25541));
    LocalMux I__5147 (
            .O(N__25556),
            .I(N__25538));
    LocalMux I__5146 (
            .O(N__25553),
            .I(\POWERLED.N_2171_i ));
    LocalMux I__5145 (
            .O(N__25548),
            .I(\POWERLED.N_2171_i ));
    Odrv4 I__5144 (
            .O(N__25541),
            .I(\POWERLED.N_2171_i ));
    Odrv12 I__5143 (
            .O(N__25538),
            .I(\POWERLED.N_2171_i ));
    CascadeMux I__5142 (
            .O(N__25529),
            .I(\POWERLED.un1_dutycycle_172_m3_ns_1_cascade_ ));
    InMux I__5141 (
            .O(N__25526),
            .I(\POWERLED.un1_count_clk_2_cry_11 ));
    InMux I__5140 (
            .O(N__25523),
            .I(N__25519));
    InMux I__5139 (
            .O(N__25522),
            .I(N__25516));
    LocalMux I__5138 (
            .O(N__25519),
            .I(\POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ));
    LocalMux I__5137 (
            .O(N__25516),
            .I(\POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ));
    InMux I__5136 (
            .O(N__25511),
            .I(\POWERLED.un1_count_clk_2_cry_12 ));
    InMux I__5135 (
            .O(N__25508),
            .I(N__25504));
    InMux I__5134 (
            .O(N__25507),
            .I(N__25501));
    LocalMux I__5133 (
            .O(N__25504),
            .I(\POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ));
    LocalMux I__5132 (
            .O(N__25501),
            .I(\POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ));
    InMux I__5131 (
            .O(N__25496),
            .I(\POWERLED.un1_count_clk_2_cry_13 ));
    InMux I__5130 (
            .O(N__25493),
            .I(\POWERLED.un1_count_clk_2_cry_14 ));
    InMux I__5129 (
            .O(N__25490),
            .I(N__25486));
    InMux I__5128 (
            .O(N__25489),
            .I(N__25483));
    LocalMux I__5127 (
            .O(N__25486),
            .I(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ));
    LocalMux I__5126 (
            .O(N__25483),
            .I(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ));
    InMux I__5125 (
            .O(N__25478),
            .I(N__25475));
    LocalMux I__5124 (
            .O(N__25475),
            .I(\POWERLED.count_clk_0_15 ));
    InMux I__5123 (
            .O(N__25472),
            .I(N__25466));
    InMux I__5122 (
            .O(N__25471),
            .I(N__25466));
    LocalMux I__5121 (
            .O(N__25466),
            .I(N__25463));
    Odrv4 I__5120 (
            .O(N__25463),
            .I(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ));
    InMux I__5119 (
            .O(N__25460),
            .I(N__25457));
    LocalMux I__5118 (
            .O(N__25457),
            .I(\POWERLED.count_clk_0_7 ));
    InMux I__5117 (
            .O(N__25454),
            .I(N__25451));
    LocalMux I__5116 (
            .O(N__25451),
            .I(N__25448));
    Span4Mux_v I__5115 (
            .O(N__25448),
            .I(N__25444));
    InMux I__5114 (
            .O(N__25447),
            .I(N__25441));
    Odrv4 I__5113 (
            .O(N__25444),
            .I(\POWERLED.N_392 ));
    LocalMux I__5112 (
            .O(N__25441),
            .I(\POWERLED.N_392 ));
    CascadeMux I__5111 (
            .O(N__25436),
            .I(N__25433));
    InMux I__5110 (
            .O(N__25433),
            .I(N__25429));
    CascadeMux I__5109 (
            .O(N__25432),
            .I(N__25426));
    LocalMux I__5108 (
            .O(N__25429),
            .I(N__25423));
    InMux I__5107 (
            .O(N__25426),
            .I(N__25420));
    Span4Mux_h I__5106 (
            .O(N__25423),
            .I(N__25417));
    LocalMux I__5105 (
            .O(N__25420),
            .I(\POWERLED.mult1_un40_sum_i_5 ));
    Odrv4 I__5104 (
            .O(N__25417),
            .I(\POWERLED.mult1_un40_sum_i_5 ));
    InMux I__5103 (
            .O(N__25412),
            .I(N__25408));
    InMux I__5102 (
            .O(N__25411),
            .I(N__25405));
    LocalMux I__5101 (
            .O(N__25408),
            .I(N__25402));
    LocalMux I__5100 (
            .O(N__25405),
            .I(N__25399));
    Span4Mux_h I__5099 (
            .O(N__25402),
            .I(N__25396));
    Odrv4 I__5098 (
            .O(N__25399),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    Odrv4 I__5097 (
            .O(N__25396),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    InMux I__5096 (
            .O(N__25391),
            .I(N__25387));
    InMux I__5095 (
            .O(N__25390),
            .I(N__25384));
    LocalMux I__5094 (
            .O(N__25387),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    LocalMux I__5093 (
            .O(N__25384),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    InMux I__5092 (
            .O(N__25379),
            .I(\POWERLED.un1_count_clk_2_cry_2 ));
    InMux I__5091 (
            .O(N__25376),
            .I(N__25372));
    InMux I__5090 (
            .O(N__25375),
            .I(N__25369));
    LocalMux I__5089 (
            .O(N__25372),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    LocalMux I__5088 (
            .O(N__25369),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    InMux I__5087 (
            .O(N__25364),
            .I(\POWERLED.un1_count_clk_2_cry_3 ));
    InMux I__5086 (
            .O(N__25361),
            .I(N__25355));
    InMux I__5085 (
            .O(N__25360),
            .I(N__25355));
    LocalMux I__5084 (
            .O(N__25355),
            .I(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ));
    InMux I__5083 (
            .O(N__25352),
            .I(\POWERLED.un1_count_clk_2_cry_4 ));
    InMux I__5082 (
            .O(N__25349),
            .I(N__25343));
    InMux I__5081 (
            .O(N__25348),
            .I(N__25343));
    LocalMux I__5080 (
            .O(N__25343),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    InMux I__5079 (
            .O(N__25340),
            .I(\POWERLED.un1_count_clk_2_cry_5 ));
    InMux I__5078 (
            .O(N__25337),
            .I(\POWERLED.un1_count_clk_2_cry_6 ));
    InMux I__5077 (
            .O(N__25334),
            .I(N__25328));
    InMux I__5076 (
            .O(N__25333),
            .I(N__25328));
    LocalMux I__5075 (
            .O(N__25328),
            .I(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ));
    InMux I__5074 (
            .O(N__25325),
            .I(\POWERLED.un1_count_clk_2_cry_7_cZ0 ));
    InMux I__5073 (
            .O(N__25322),
            .I(N__25316));
    InMux I__5072 (
            .O(N__25321),
            .I(N__25316));
    LocalMux I__5071 (
            .O(N__25316),
            .I(N__25313));
    Odrv4 I__5070 (
            .O(N__25313),
            .I(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ));
    InMux I__5069 (
            .O(N__25310),
            .I(bfn_9_8_0_));
    InMux I__5068 (
            .O(N__25307),
            .I(\POWERLED.un1_count_clk_2_cry_9_cZ0 ));
    InMux I__5067 (
            .O(N__25304),
            .I(\POWERLED.un1_count_clk_2_cry_10_cZ0 ));
    InMux I__5066 (
            .O(N__25301),
            .I(N__25298));
    LocalMux I__5065 (
            .O(N__25298),
            .I(\POWERLED.count_clk_0_5 ));
    InMux I__5064 (
            .O(N__25295),
            .I(N__25292));
    LocalMux I__5063 (
            .O(N__25292),
            .I(\POWERLED.count_clk_0_6 ));
    InMux I__5062 (
            .O(N__25289),
            .I(N__25286));
    LocalMux I__5061 (
            .O(N__25286),
            .I(\POWERLED.count_clk_0_8 ));
    InMux I__5060 (
            .O(N__25283),
            .I(N__25280));
    LocalMux I__5059 (
            .O(N__25280),
            .I(\POWERLED.count_clk_0_9 ));
    CascadeMux I__5058 (
            .O(N__25277),
            .I(N__25273));
    InMux I__5057 (
            .O(N__25276),
            .I(N__25270));
    InMux I__5056 (
            .O(N__25273),
            .I(N__25267));
    LocalMux I__5055 (
            .O(N__25270),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    LocalMux I__5054 (
            .O(N__25267),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    InMux I__5053 (
            .O(N__25262),
            .I(\POWERLED.un1_count_clk_2_cry_1 ));
    InMux I__5052 (
            .O(N__25259),
            .I(N__25256));
    LocalMux I__5051 (
            .O(N__25256),
            .I(\POWERLED.un34_clk_100khz_5 ));
    InMux I__5050 (
            .O(N__25253),
            .I(N__25250));
    LocalMux I__5049 (
            .O(N__25250),
            .I(N__25244));
    InMux I__5048 (
            .O(N__25249),
            .I(N__25237));
    InMux I__5047 (
            .O(N__25248),
            .I(N__25237));
    InMux I__5046 (
            .O(N__25247),
            .I(N__25237));
    Span4Mux_h I__5045 (
            .O(N__25244),
            .I(N__25232));
    LocalMux I__5044 (
            .O(N__25237),
            .I(N__25232));
    Span4Mux_h I__5043 (
            .O(N__25232),
            .I(N__25229));
    Span4Mux_v I__5042 (
            .O(N__25229),
            .I(N__25226));
    Odrv4 I__5041 (
            .O(N__25226),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    CascadeMux I__5040 (
            .O(N__25223),
            .I(N__25220));
    InMux I__5039 (
            .O(N__25220),
            .I(N__25215));
    InMux I__5038 (
            .O(N__25219),
            .I(N__25208));
    InMux I__5037 (
            .O(N__25218),
            .I(N__25208));
    LocalMux I__5036 (
            .O(N__25215),
            .I(N__25205));
    InMux I__5035 (
            .O(N__25214),
            .I(N__25200));
    InMux I__5034 (
            .O(N__25213),
            .I(N__25200));
    LocalMux I__5033 (
            .O(N__25208),
            .I(N__25197));
    Odrv12 I__5032 (
            .O(N__25205),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__5031 (
            .O(N__25200),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__5030 (
            .O(N__25197),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    InMux I__5029 (
            .O(N__25190),
            .I(N__25187));
    LocalMux I__5028 (
            .O(N__25187),
            .I(N__25184));
    Span4Mux_h I__5027 (
            .O(N__25184),
            .I(N__25178));
    InMux I__5026 (
            .O(N__25183),
            .I(N__25175));
    InMux I__5025 (
            .O(N__25182),
            .I(N__25170));
    InMux I__5024 (
            .O(N__25181),
            .I(N__25170));
    Odrv4 I__5023 (
            .O(N__25178),
            .I(\POWERLED.count_RNIZ0Z_15 ));
    LocalMux I__5022 (
            .O(N__25175),
            .I(\POWERLED.count_RNIZ0Z_15 ));
    LocalMux I__5021 (
            .O(N__25170),
            .I(\POWERLED.count_RNIZ0Z_15 ));
    InMux I__5020 (
            .O(N__25163),
            .I(N__25160));
    LocalMux I__5019 (
            .O(N__25160),
            .I(N__25157));
    Span4Mux_h I__5018 (
            .O(N__25157),
            .I(N__25154));
    Odrv4 I__5017 (
            .O(N__25154),
            .I(\POWERLED.curr_state_1_0 ));
    CascadeMux I__5016 (
            .O(N__25151),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1_cascade_ ));
    InMux I__5015 (
            .O(N__25148),
            .I(N__25145));
    LocalMux I__5014 (
            .O(N__25145),
            .I(N__25142));
    Span4Mux_h I__5013 (
            .O(N__25142),
            .I(N__25137));
    InMux I__5012 (
            .O(N__25141),
            .I(N__25133));
    InMux I__5011 (
            .O(N__25140),
            .I(N__25130));
    Span4Mux_v I__5010 (
            .O(N__25137),
            .I(N__25127));
    InMux I__5009 (
            .O(N__25136),
            .I(N__25124));
    LocalMux I__5008 (
            .O(N__25133),
            .I(N__25121));
    LocalMux I__5007 (
            .O(N__25130),
            .I(N__25118));
    Odrv4 I__5006 (
            .O(N__25127),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__5005 (
            .O(N__25124),
            .I(\POWERLED.countZ0Z_1 ));
    Odrv4 I__5004 (
            .O(N__25121),
            .I(\POWERLED.countZ0Z_1 ));
    Odrv4 I__5003 (
            .O(N__25118),
            .I(\POWERLED.countZ0Z_1 ));
    InMux I__5002 (
            .O(N__25109),
            .I(N__25106));
    LocalMux I__5001 (
            .O(N__25106),
            .I(N__25103));
    Odrv12 I__5000 (
            .O(N__25103),
            .I(\POWERLED.count_0_1 ));
    InMux I__4999 (
            .O(N__25100),
            .I(N__25095));
    CascadeMux I__4998 (
            .O(N__25099),
            .I(N__25092));
    CascadeMux I__4997 (
            .O(N__25098),
            .I(N__25088));
    LocalMux I__4996 (
            .O(N__25095),
            .I(N__25085));
    InMux I__4995 (
            .O(N__25092),
            .I(N__25079));
    InMux I__4994 (
            .O(N__25091),
            .I(N__25079));
    InMux I__4993 (
            .O(N__25088),
            .I(N__25075));
    Span4Mux_s3_h I__4992 (
            .O(N__25085),
            .I(N__25072));
    InMux I__4991 (
            .O(N__25084),
            .I(N__25069));
    LocalMux I__4990 (
            .O(N__25079),
            .I(N__25066));
    InMux I__4989 (
            .O(N__25078),
            .I(N__25063));
    LocalMux I__4988 (
            .O(N__25075),
            .I(N__25060));
    Span4Mux_v I__4987 (
            .O(N__25072),
            .I(N__25051));
    LocalMux I__4986 (
            .O(N__25069),
            .I(N__25051));
    Span4Mux_h I__4985 (
            .O(N__25066),
            .I(N__25051));
    LocalMux I__4984 (
            .O(N__25063),
            .I(N__25051));
    Odrv4 I__4983 (
            .O(N__25060),
            .I(\POWERLED.countZ0Z_0 ));
    Odrv4 I__4982 (
            .O(N__25051),
            .I(\POWERLED.countZ0Z_0 ));
    InMux I__4981 (
            .O(N__25046),
            .I(N__25027));
    InMux I__4980 (
            .O(N__25045),
            .I(N__25024));
    InMux I__4979 (
            .O(N__25044),
            .I(N__25021));
    InMux I__4978 (
            .O(N__25043),
            .I(N__25014));
    InMux I__4977 (
            .O(N__25042),
            .I(N__25014));
    InMux I__4976 (
            .O(N__25041),
            .I(N__25014));
    InMux I__4975 (
            .O(N__25040),
            .I(N__25005));
    InMux I__4974 (
            .O(N__25039),
            .I(N__25005));
    InMux I__4973 (
            .O(N__25038),
            .I(N__25005));
    InMux I__4972 (
            .O(N__25037),
            .I(N__25005));
    InMux I__4971 (
            .O(N__25036),
            .I(N__24998));
    InMux I__4970 (
            .O(N__25035),
            .I(N__24998));
    InMux I__4969 (
            .O(N__25034),
            .I(N__24998));
    InMux I__4968 (
            .O(N__25033),
            .I(N__24989));
    InMux I__4967 (
            .O(N__25032),
            .I(N__24989));
    InMux I__4966 (
            .O(N__25031),
            .I(N__24989));
    InMux I__4965 (
            .O(N__25030),
            .I(N__24989));
    LocalMux I__4964 (
            .O(N__25027),
            .I(N__24986));
    LocalMux I__4963 (
            .O(N__25024),
            .I(N__24981));
    LocalMux I__4962 (
            .O(N__25021),
            .I(N__24981));
    LocalMux I__4961 (
            .O(N__25014),
            .I(N__24972));
    LocalMux I__4960 (
            .O(N__25005),
            .I(N__24972));
    LocalMux I__4959 (
            .O(N__24998),
            .I(N__24972));
    LocalMux I__4958 (
            .O(N__24989),
            .I(N__24972));
    Odrv4 I__4957 (
            .O(N__24986),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv12 I__4956 (
            .O(N__24981),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv4 I__4955 (
            .O(N__24972),
            .I(\POWERLED.count_0_sqmuxa_i ));
    InMux I__4954 (
            .O(N__24965),
            .I(N__24962));
    LocalMux I__4953 (
            .O(N__24962),
            .I(N__24959));
    Odrv12 I__4952 (
            .O(N__24959),
            .I(\POWERLED.count_0_0 ));
    CascadeMux I__4951 (
            .O(N__24956),
            .I(N__24947));
    CascadeMux I__4950 (
            .O(N__24955),
            .I(N__24943));
    InMux I__4949 (
            .O(N__24954),
            .I(N__24935));
    InMux I__4948 (
            .O(N__24953),
            .I(N__24935));
    InMux I__4947 (
            .O(N__24952),
            .I(N__24935));
    InMux I__4946 (
            .O(N__24951),
            .I(N__24930));
    InMux I__4945 (
            .O(N__24950),
            .I(N__24930));
    InMux I__4944 (
            .O(N__24947),
            .I(N__24923));
    InMux I__4943 (
            .O(N__24946),
            .I(N__24923));
    InMux I__4942 (
            .O(N__24943),
            .I(N__24923));
    InMux I__4941 (
            .O(N__24942),
            .I(N__24919));
    LocalMux I__4940 (
            .O(N__24935),
            .I(N__24916));
    LocalMux I__4939 (
            .O(N__24930),
            .I(N__24911));
    LocalMux I__4938 (
            .O(N__24923),
            .I(N__24911));
    InMux I__4937 (
            .O(N__24922),
            .I(N__24908));
    LocalMux I__4936 (
            .O(N__24919),
            .I(N__24903));
    Span4Mux_v I__4935 (
            .O(N__24916),
            .I(N__24900));
    Span4Mux_v I__4934 (
            .O(N__24911),
            .I(N__24895));
    LocalMux I__4933 (
            .O(N__24908),
            .I(N__24895));
    InMux I__4932 (
            .O(N__24907),
            .I(N__24890));
    InMux I__4931 (
            .O(N__24906),
            .I(N__24890));
    Span4Mux_v I__4930 (
            .O(N__24903),
            .I(N__24887));
    Span4Mux_v I__4929 (
            .O(N__24900),
            .I(N__24882));
    Span4Mux_v I__4928 (
            .O(N__24895),
            .I(N__24882));
    LocalMux I__4927 (
            .O(N__24890),
            .I(N__24879));
    Sp12to4 I__4926 (
            .O(N__24887),
            .I(N__24876));
    Span4Mux_h I__4925 (
            .O(N__24882),
            .I(N__24873));
    Span4Mux_h I__4924 (
            .O(N__24879),
            .I(N__24870));
    Span12Mux_s8_h I__4923 (
            .O(N__24876),
            .I(N__24867));
    Span4Mux_v I__4922 (
            .O(N__24873),
            .I(N__24862));
    Span4Mux_v I__4921 (
            .O(N__24870),
            .I(N__24862));
    Odrv12 I__4920 (
            .O(N__24867),
            .I(slp_s4n));
    Odrv4 I__4919 (
            .O(N__24862),
            .I(slp_s4n));
    InMux I__4918 (
            .O(N__24857),
            .I(N__24854));
    LocalMux I__4917 (
            .O(N__24854),
            .I(N__24850));
    InMux I__4916 (
            .O(N__24853),
            .I(N__24846));
    Span4Mux_h I__4915 (
            .O(N__24850),
            .I(N__24841));
    InMux I__4914 (
            .O(N__24849),
            .I(N__24838));
    LocalMux I__4913 (
            .O(N__24846),
            .I(N__24835));
    InMux I__4912 (
            .O(N__24845),
            .I(N__24832));
    InMux I__4911 (
            .O(N__24844),
            .I(N__24829));
    Span4Mux_v I__4910 (
            .O(N__24841),
            .I(N__24826));
    LocalMux I__4909 (
            .O(N__24838),
            .I(N__24821));
    Span4Mux_v I__4908 (
            .O(N__24835),
            .I(N__24821));
    LocalMux I__4907 (
            .O(N__24832),
            .I(N__24816));
    LocalMux I__4906 (
            .O(N__24829),
            .I(N__24816));
    Odrv4 I__4905 (
            .O(N__24826),
            .I(RSMRST_PWRGD_RSMRSTn_2_fast));
    Odrv4 I__4904 (
            .O(N__24821),
            .I(RSMRST_PWRGD_RSMRSTn_2_fast));
    Odrv12 I__4903 (
            .O(N__24816),
            .I(RSMRST_PWRGD_RSMRSTn_2_fast));
    InMux I__4902 (
            .O(N__24809),
            .I(N__24804));
    InMux I__4901 (
            .O(N__24808),
            .I(N__24801));
    InMux I__4900 (
            .O(N__24807),
            .I(N__24798));
    LocalMux I__4899 (
            .O(N__24804),
            .I(N__24791));
    LocalMux I__4898 (
            .O(N__24801),
            .I(N__24791));
    LocalMux I__4897 (
            .O(N__24798),
            .I(N__24791));
    Odrv4 I__4896 (
            .O(N__24791),
            .I(\POWERLED.N_150_i ));
    InMux I__4895 (
            .O(N__24788),
            .I(N__24785));
    LocalMux I__4894 (
            .O(N__24785),
            .I(N__24782));
    Span4Mux_h I__4893 (
            .O(N__24782),
            .I(N__24774));
    InMux I__4892 (
            .O(N__24781),
            .I(N__24771));
    InMux I__4891 (
            .O(N__24780),
            .I(N__24768));
    InMux I__4890 (
            .O(N__24779),
            .I(N__24765));
    InMux I__4889 (
            .O(N__24778),
            .I(N__24762));
    InMux I__4888 (
            .O(N__24777),
            .I(N__24759));
    Odrv4 I__4887 (
            .O(N__24774),
            .I(\POWERLED.N_154 ));
    LocalMux I__4886 (
            .O(N__24771),
            .I(\POWERLED.N_154 ));
    LocalMux I__4885 (
            .O(N__24768),
            .I(\POWERLED.N_154 ));
    LocalMux I__4884 (
            .O(N__24765),
            .I(\POWERLED.N_154 ));
    LocalMux I__4883 (
            .O(N__24762),
            .I(\POWERLED.N_154 ));
    LocalMux I__4882 (
            .O(N__24759),
            .I(\POWERLED.N_154 ));
    InMux I__4881 (
            .O(N__24746),
            .I(N__24743));
    LocalMux I__4880 (
            .O(N__24743),
            .I(\POWERLED.N_389 ));
    InMux I__4879 (
            .O(N__24740),
            .I(N__24737));
    LocalMux I__4878 (
            .O(N__24737),
            .I(\POWERLED.count_off_0_10 ));
    InMux I__4877 (
            .O(N__24734),
            .I(N__24728));
    InMux I__4876 (
            .O(N__24733),
            .I(N__24728));
    LocalMux I__4875 (
            .O(N__24728),
            .I(\POWERLED.count_off_1_9 ));
    InMux I__4874 (
            .O(N__24725),
            .I(N__24719));
    InMux I__4873 (
            .O(N__24724),
            .I(N__24719));
    LocalMux I__4872 (
            .O(N__24719),
            .I(\POWERLED.count_offZ0Z_9 ));
    CascadeMux I__4871 (
            .O(N__24716),
            .I(\POWERLED.count_offZ0Z_10_cascade_ ));
    CascadeMux I__4870 (
            .O(N__24713),
            .I(\POWERLED.un34_clk_100khz_4_cascade_ ));
    InMux I__4869 (
            .O(N__24710),
            .I(N__24706));
    InMux I__4868 (
            .O(N__24709),
            .I(N__24703));
    LocalMux I__4867 (
            .O(N__24706),
            .I(\HDA_STRAP.countZ0Z_13 ));
    LocalMux I__4866 (
            .O(N__24703),
            .I(\HDA_STRAP.countZ0Z_13 ));
    InMux I__4865 (
            .O(N__24698),
            .I(\HDA_STRAP.un1_count_1_cry_12 ));
    InMux I__4864 (
            .O(N__24695),
            .I(N__24691));
    InMux I__4863 (
            .O(N__24694),
            .I(N__24688));
    LocalMux I__4862 (
            .O(N__24691),
            .I(\HDA_STRAP.countZ0Z_14 ));
    LocalMux I__4861 (
            .O(N__24688),
            .I(\HDA_STRAP.countZ0Z_14 ));
    InMux I__4860 (
            .O(N__24683),
            .I(\HDA_STRAP.un1_count_1_cry_13 ));
    InMux I__4859 (
            .O(N__24680),
            .I(N__24676));
    InMux I__4858 (
            .O(N__24679),
            .I(N__24673));
    LocalMux I__4857 (
            .O(N__24676),
            .I(\HDA_STRAP.countZ0Z_15 ));
    LocalMux I__4856 (
            .O(N__24673),
            .I(\HDA_STRAP.countZ0Z_15 ));
    InMux I__4855 (
            .O(N__24668),
            .I(\HDA_STRAP.un1_count_1_cry_14 ));
    InMux I__4854 (
            .O(N__24665),
            .I(N__24661));
    InMux I__4853 (
            .O(N__24664),
            .I(N__24658));
    LocalMux I__4852 (
            .O(N__24661),
            .I(\HDA_STRAP.countZ0Z_16 ));
    LocalMux I__4851 (
            .O(N__24658),
            .I(\HDA_STRAP.countZ0Z_16 ));
    InMux I__4850 (
            .O(N__24653),
            .I(N__24650));
    LocalMux I__4849 (
            .O(N__24650),
            .I(\HDA_STRAP.count_RNO_0Z0Z_16 ));
    InMux I__4848 (
            .O(N__24647),
            .I(bfn_9_3_0_));
    InMux I__4847 (
            .O(N__24644),
            .I(N__24641));
    LocalMux I__4846 (
            .O(N__24641),
            .I(N__24638));
    Span4Mux_h I__4845 (
            .O(N__24638),
            .I(N__24634));
    InMux I__4844 (
            .O(N__24637),
            .I(N__24631));
    Odrv4 I__4843 (
            .O(N__24634),
            .I(\HDA_STRAP.countZ0Z_17 ));
    LocalMux I__4842 (
            .O(N__24631),
            .I(\HDA_STRAP.countZ0Z_17 ));
    InMux I__4841 (
            .O(N__24626),
            .I(\HDA_STRAP.un1_count_1_cry_16 ));
    InMux I__4840 (
            .O(N__24623),
            .I(N__24620));
    LocalMux I__4839 (
            .O(N__24620),
            .I(N__24617));
    Span4Mux_s2_v I__4838 (
            .O(N__24617),
            .I(N__24614));
    Odrv4 I__4837 (
            .O(N__24614),
            .I(\HDA_STRAP.count_RNO_0Z0Z_17 ));
    InMux I__4836 (
            .O(N__24611),
            .I(N__24608));
    LocalMux I__4835 (
            .O(N__24608),
            .I(N__24605));
    Odrv4 I__4834 (
            .O(N__24605),
            .I(\POWERLED.un1_func_state25_6_0_a2_1 ));
    CascadeMux I__4833 (
            .O(N__24602),
            .I(\POWERLED.un1_func_state25_6_0_o_N_305_N_cascade_ ));
    CascadeMux I__4832 (
            .O(N__24599),
            .I(\POWERLED.un1_func_state25_6_0_0_cascade_ ));
    CascadeMux I__4831 (
            .O(N__24596),
            .I(N__24593));
    InMux I__4830 (
            .O(N__24593),
            .I(N__24590));
    LocalMux I__4829 (
            .O(N__24590),
            .I(\POWERLED.un1_func_state25_6_0_1 ));
    InMux I__4828 (
            .O(N__24587),
            .I(\HDA_STRAP.un1_count_1_cry_3 ));
    InMux I__4827 (
            .O(N__24584),
            .I(N__24580));
    InMux I__4826 (
            .O(N__24583),
            .I(N__24577));
    LocalMux I__4825 (
            .O(N__24580),
            .I(\HDA_STRAP.countZ0Z_5 ));
    LocalMux I__4824 (
            .O(N__24577),
            .I(\HDA_STRAP.countZ0Z_5 ));
    InMux I__4823 (
            .O(N__24572),
            .I(\HDA_STRAP.un1_count_1_cry_4 ));
    InMux I__4822 (
            .O(N__24569),
            .I(N__24565));
    InMux I__4821 (
            .O(N__24568),
            .I(N__24562));
    LocalMux I__4820 (
            .O(N__24565),
            .I(\HDA_STRAP.countZ0Z_6 ));
    LocalMux I__4819 (
            .O(N__24562),
            .I(\HDA_STRAP.countZ0Z_6 ));
    CascadeMux I__4818 (
            .O(N__24557),
            .I(N__24554));
    InMux I__4817 (
            .O(N__24554),
            .I(N__24551));
    LocalMux I__4816 (
            .O(N__24551),
            .I(\HDA_STRAP.count_RNO_0Z0Z_6 ));
    InMux I__4815 (
            .O(N__24548),
            .I(\HDA_STRAP.un1_count_1_cry_5 ));
    CascadeMux I__4814 (
            .O(N__24545),
            .I(N__24542));
    InMux I__4813 (
            .O(N__24542),
            .I(N__24539));
    LocalMux I__4812 (
            .O(N__24539),
            .I(N__24535));
    InMux I__4811 (
            .O(N__24538),
            .I(N__24532));
    Odrv4 I__4810 (
            .O(N__24535),
            .I(\HDA_STRAP.countZ0Z_7 ));
    LocalMux I__4809 (
            .O(N__24532),
            .I(\HDA_STRAP.countZ0Z_7 ));
    InMux I__4808 (
            .O(N__24527),
            .I(\HDA_STRAP.un1_count_1_cry_6 ));
    CascadeMux I__4807 (
            .O(N__24524),
            .I(N__24521));
    InMux I__4806 (
            .O(N__24521),
            .I(N__24517));
    InMux I__4805 (
            .O(N__24520),
            .I(N__24514));
    LocalMux I__4804 (
            .O(N__24517),
            .I(\HDA_STRAP.countZ0Z_8 ));
    LocalMux I__4803 (
            .O(N__24514),
            .I(\HDA_STRAP.countZ0Z_8 ));
    InMux I__4802 (
            .O(N__24509),
            .I(N__24506));
    LocalMux I__4801 (
            .O(N__24506),
            .I(\HDA_STRAP.count_RNO_0Z0Z_8 ));
    InMux I__4800 (
            .O(N__24503),
            .I(bfn_9_2_0_));
    InMux I__4799 (
            .O(N__24500),
            .I(N__24496));
    InMux I__4798 (
            .O(N__24499),
            .I(N__24493));
    LocalMux I__4797 (
            .O(N__24496),
            .I(\HDA_STRAP.countZ0Z_9 ));
    LocalMux I__4796 (
            .O(N__24493),
            .I(\HDA_STRAP.countZ0Z_9 ));
    InMux I__4795 (
            .O(N__24488),
            .I(\HDA_STRAP.un1_count_1_cry_8 ));
    InMux I__4794 (
            .O(N__24485),
            .I(N__24481));
    InMux I__4793 (
            .O(N__24484),
            .I(N__24478));
    LocalMux I__4792 (
            .O(N__24481),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__4791 (
            .O(N__24478),
            .I(\HDA_STRAP.countZ0Z_10 ));
    CascadeMux I__4790 (
            .O(N__24473),
            .I(N__24470));
    InMux I__4789 (
            .O(N__24470),
            .I(N__24467));
    LocalMux I__4788 (
            .O(N__24467),
            .I(\HDA_STRAP.count_RNO_0Z0Z_10 ));
    InMux I__4787 (
            .O(N__24464),
            .I(\HDA_STRAP.un1_count_1_cry_9 ));
    InMux I__4786 (
            .O(N__24461),
            .I(N__24457));
    InMux I__4785 (
            .O(N__24460),
            .I(N__24454));
    LocalMux I__4784 (
            .O(N__24457),
            .I(\HDA_STRAP.countZ0Z_11 ));
    LocalMux I__4783 (
            .O(N__24454),
            .I(\HDA_STRAP.countZ0Z_11 ));
    InMux I__4782 (
            .O(N__24449),
            .I(N__24446));
    LocalMux I__4781 (
            .O(N__24446),
            .I(\HDA_STRAP.count_RNO_0Z0Z_11 ));
    InMux I__4780 (
            .O(N__24443),
            .I(\HDA_STRAP.un1_count_1_cry_10 ));
    InMux I__4779 (
            .O(N__24440),
            .I(N__24436));
    InMux I__4778 (
            .O(N__24439),
            .I(N__24433));
    LocalMux I__4777 (
            .O(N__24436),
            .I(\HDA_STRAP.countZ0Z_12 ));
    LocalMux I__4776 (
            .O(N__24433),
            .I(\HDA_STRAP.countZ0Z_12 ));
    InMux I__4775 (
            .O(N__24428),
            .I(\HDA_STRAP.un1_count_1_cry_11 ));
    CascadeMux I__4774 (
            .O(N__24425),
            .I(N__24417));
    CascadeMux I__4773 (
            .O(N__24424),
            .I(N__24410));
    CascadeMux I__4772 (
            .O(N__24423),
            .I(N__24407));
    InMux I__4771 (
            .O(N__24422),
            .I(N__24403));
    CascadeMux I__4770 (
            .O(N__24421),
            .I(N__24399));
    CascadeMux I__4769 (
            .O(N__24420),
            .I(N__24395));
    InMux I__4768 (
            .O(N__24417),
            .I(N__24389));
    InMux I__4767 (
            .O(N__24416),
            .I(N__24389));
    InMux I__4766 (
            .O(N__24415),
            .I(N__24383));
    InMux I__4765 (
            .O(N__24414),
            .I(N__24378));
    InMux I__4764 (
            .O(N__24413),
            .I(N__24378));
    InMux I__4763 (
            .O(N__24410),
            .I(N__24373));
    InMux I__4762 (
            .O(N__24407),
            .I(N__24373));
    CascadeMux I__4761 (
            .O(N__24406),
            .I(N__24370));
    LocalMux I__4760 (
            .O(N__24403),
            .I(N__24367));
    InMux I__4759 (
            .O(N__24402),
            .I(N__24358));
    InMux I__4758 (
            .O(N__24399),
            .I(N__24358));
    InMux I__4757 (
            .O(N__24398),
            .I(N__24358));
    InMux I__4756 (
            .O(N__24395),
            .I(N__24358));
    InMux I__4755 (
            .O(N__24394),
            .I(N__24353));
    LocalMux I__4754 (
            .O(N__24389),
            .I(N__24350));
    InMux I__4753 (
            .O(N__24388),
            .I(N__24345));
    InMux I__4752 (
            .O(N__24387),
            .I(N__24345));
    CascadeMux I__4751 (
            .O(N__24386),
            .I(N__24339));
    LocalMux I__4750 (
            .O(N__24383),
            .I(N__24334));
    LocalMux I__4749 (
            .O(N__24378),
            .I(N__24334));
    LocalMux I__4748 (
            .O(N__24373),
            .I(N__24331));
    InMux I__4747 (
            .O(N__24370),
            .I(N__24328));
    Span4Mux_v I__4746 (
            .O(N__24367),
            .I(N__24323));
    LocalMux I__4745 (
            .O(N__24358),
            .I(N__24323));
    InMux I__4744 (
            .O(N__24357),
            .I(N__24318));
    InMux I__4743 (
            .O(N__24356),
            .I(N__24318));
    LocalMux I__4742 (
            .O(N__24353),
            .I(N__24311));
    Span4Mux_h I__4741 (
            .O(N__24350),
            .I(N__24311));
    LocalMux I__4740 (
            .O(N__24345),
            .I(N__24311));
    InMux I__4739 (
            .O(N__24344),
            .I(N__24302));
    InMux I__4738 (
            .O(N__24343),
            .I(N__24302));
    InMux I__4737 (
            .O(N__24342),
            .I(N__24302));
    InMux I__4736 (
            .O(N__24339),
            .I(N__24302));
    Span4Mux_h I__4735 (
            .O(N__24334),
            .I(N__24295));
    Span4Mux_v I__4734 (
            .O(N__24331),
            .I(N__24295));
    LocalMux I__4733 (
            .O(N__24328),
            .I(N__24295));
    Odrv4 I__4732 (
            .O(N__24323),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__4731 (
            .O(N__24318),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__4730 (
            .O(N__24311),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__4729 (
            .O(N__24302),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__4728 (
            .O(N__24295),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    InMux I__4727 (
            .O(N__24284),
            .I(N__24276));
    InMux I__4726 (
            .O(N__24283),
            .I(N__24271));
    InMux I__4725 (
            .O(N__24282),
            .I(N__24271));
    InMux I__4724 (
            .O(N__24281),
            .I(N__24260));
    InMux I__4723 (
            .O(N__24280),
            .I(N__24255));
    InMux I__4722 (
            .O(N__24279),
            .I(N__24255));
    LocalMux I__4721 (
            .O(N__24276),
            .I(N__24250));
    LocalMux I__4720 (
            .O(N__24271),
            .I(N__24250));
    InMux I__4719 (
            .O(N__24270),
            .I(N__24241));
    InMux I__4718 (
            .O(N__24269),
            .I(N__24241));
    InMux I__4717 (
            .O(N__24268),
            .I(N__24241));
    InMux I__4716 (
            .O(N__24267),
            .I(N__24238));
    InMux I__4715 (
            .O(N__24266),
            .I(N__24235));
    CascadeMux I__4714 (
            .O(N__24265),
            .I(N__24232));
    InMux I__4713 (
            .O(N__24264),
            .I(N__24229));
    InMux I__4712 (
            .O(N__24263),
            .I(N__24226));
    LocalMux I__4711 (
            .O(N__24260),
            .I(N__24223));
    LocalMux I__4710 (
            .O(N__24255),
            .I(N__24218));
    Span4Mux_v I__4709 (
            .O(N__24250),
            .I(N__24218));
    InMux I__4708 (
            .O(N__24249),
            .I(N__24213));
    InMux I__4707 (
            .O(N__24248),
            .I(N__24213));
    LocalMux I__4706 (
            .O(N__24241),
            .I(N__24206));
    LocalMux I__4705 (
            .O(N__24238),
            .I(N__24206));
    LocalMux I__4704 (
            .O(N__24235),
            .I(N__24206));
    InMux I__4703 (
            .O(N__24232),
            .I(N__24203));
    LocalMux I__4702 (
            .O(N__24229),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__4701 (
            .O(N__24226),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__4700 (
            .O(N__24223),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__4699 (
            .O(N__24218),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__4698 (
            .O(N__24213),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__4697 (
            .O(N__24206),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__4696 (
            .O(N__24203),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    CascadeMux I__4695 (
            .O(N__24188),
            .I(\POWERLED.g0_i_a6_0_1_cascade_ ));
    InMux I__4694 (
            .O(N__24185),
            .I(N__24182));
    LocalMux I__4693 (
            .O(N__24182),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_12 ));
    InMux I__4692 (
            .O(N__24179),
            .I(N__24176));
    LocalMux I__4691 (
            .O(N__24176),
            .I(N__24172));
    InMux I__4690 (
            .O(N__24175),
            .I(N__24169));
    Span4Mux_s2_v I__4689 (
            .O(N__24172),
            .I(N__24164));
    LocalMux I__4688 (
            .O(N__24169),
            .I(N__24161));
    InMux I__4687 (
            .O(N__24168),
            .I(N__24153));
    InMux I__4686 (
            .O(N__24167),
            .I(N__24149));
    Span4Mux_h I__4685 (
            .O(N__24164),
            .I(N__24146));
    Span4Mux_h I__4684 (
            .O(N__24161),
            .I(N__24143));
    InMux I__4683 (
            .O(N__24160),
            .I(N__24136));
    InMux I__4682 (
            .O(N__24159),
            .I(N__24136));
    InMux I__4681 (
            .O(N__24158),
            .I(N__24136));
    InMux I__4680 (
            .O(N__24157),
            .I(N__24131));
    InMux I__4679 (
            .O(N__24156),
            .I(N__24131));
    LocalMux I__4678 (
            .O(N__24153),
            .I(N__24128));
    InMux I__4677 (
            .O(N__24152),
            .I(N__24125));
    LocalMux I__4676 (
            .O(N__24149),
            .I(N__24122));
    Odrv4 I__4675 (
            .O(N__24146),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__4674 (
            .O(N__24143),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__4673 (
            .O(N__24136),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__4672 (
            .O(N__24131),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv12 I__4671 (
            .O(N__24128),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__4670 (
            .O(N__24125),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__4669 (
            .O(N__24122),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    CascadeMux I__4668 (
            .O(N__24107),
            .I(N__24101));
    InMux I__4667 (
            .O(N__24106),
            .I(N__24094));
    InMux I__4666 (
            .O(N__24105),
            .I(N__24094));
    InMux I__4665 (
            .O(N__24104),
            .I(N__24091));
    InMux I__4664 (
            .O(N__24101),
            .I(N__24088));
    CascadeMux I__4663 (
            .O(N__24100),
            .I(N__24084));
    InMux I__4662 (
            .O(N__24099),
            .I(N__24077));
    LocalMux I__4661 (
            .O(N__24094),
            .I(N__24074));
    LocalMux I__4660 (
            .O(N__24091),
            .I(N__24069));
    LocalMux I__4659 (
            .O(N__24088),
            .I(N__24069));
    InMux I__4658 (
            .O(N__24087),
            .I(N__24066));
    InMux I__4657 (
            .O(N__24084),
            .I(N__24063));
    InMux I__4656 (
            .O(N__24083),
            .I(N__24056));
    InMux I__4655 (
            .O(N__24082),
            .I(N__24056));
    InMux I__4654 (
            .O(N__24081),
            .I(N__24056));
    InMux I__4653 (
            .O(N__24080),
            .I(N__24053));
    LocalMux I__4652 (
            .O(N__24077),
            .I(N__24050));
    Span4Mux_s3_v I__4651 (
            .O(N__24074),
            .I(N__24047));
    Span12Mux_s7_h I__4650 (
            .O(N__24069),
            .I(N__24036));
    LocalMux I__4649 (
            .O(N__24066),
            .I(N__24036));
    LocalMux I__4648 (
            .O(N__24063),
            .I(N__24036));
    LocalMux I__4647 (
            .O(N__24056),
            .I(N__24036));
    LocalMux I__4646 (
            .O(N__24053),
            .I(N__24036));
    Span4Mux_h I__4645 (
            .O(N__24050),
            .I(N__24033));
    Span4Mux_v I__4644 (
            .O(N__24047),
            .I(N__24030));
    Span12Mux_s5_v I__4643 (
            .O(N__24036),
            .I(N__24027));
    Odrv4 I__4642 (
            .O(N__24033),
            .I(\POWERLED.func_state_RNIC4OR2Z0Z_0 ));
    Odrv4 I__4641 (
            .O(N__24030),
            .I(\POWERLED.func_state_RNIC4OR2Z0Z_0 ));
    Odrv12 I__4640 (
            .O(N__24027),
            .I(\POWERLED.func_state_RNIC4OR2Z0Z_0 ));
    InMux I__4639 (
            .O(N__24020),
            .I(N__24014));
    InMux I__4638 (
            .O(N__24019),
            .I(N__24014));
    LocalMux I__4637 (
            .O(N__24014),
            .I(N__24005));
    InMux I__4636 (
            .O(N__24013),
            .I(N__24001));
    InMux I__4635 (
            .O(N__24012),
            .I(N__23996));
    InMux I__4634 (
            .O(N__24011),
            .I(N__23996));
    InMux I__4633 (
            .O(N__24010),
            .I(N__23989));
    InMux I__4632 (
            .O(N__24009),
            .I(N__23989));
    InMux I__4631 (
            .O(N__24008),
            .I(N__23989));
    Span4Mux_v I__4630 (
            .O(N__24005),
            .I(N__23986));
    InMux I__4629 (
            .O(N__24004),
            .I(N__23983));
    LocalMux I__4628 (
            .O(N__24001),
            .I(N__23976));
    LocalMux I__4627 (
            .O(N__23996),
            .I(N__23976));
    LocalMux I__4626 (
            .O(N__23989),
            .I(N__23976));
    Span4Mux_h I__4625 (
            .O(N__23986),
            .I(N__23971));
    LocalMux I__4624 (
            .O(N__23983),
            .I(N__23966));
    Span4Mux_v I__4623 (
            .O(N__23976),
            .I(N__23966));
    InMux I__4622 (
            .O(N__23975),
            .I(N__23961));
    InMux I__4621 (
            .O(N__23974),
            .I(N__23961));
    Odrv4 I__4620 (
            .O(N__23971),
            .I(\POWERLED.N_390 ));
    Odrv4 I__4619 (
            .O(N__23966),
            .I(\POWERLED.N_390 ));
    LocalMux I__4618 (
            .O(N__23961),
            .I(\POWERLED.N_390 ));
    InMux I__4617 (
            .O(N__23954),
            .I(N__23941));
    InMux I__4616 (
            .O(N__23953),
            .I(N__23938));
    InMux I__4615 (
            .O(N__23952),
            .I(N__23935));
    InMux I__4614 (
            .O(N__23951),
            .I(N__23932));
    InMux I__4613 (
            .O(N__23950),
            .I(N__23929));
    InMux I__4612 (
            .O(N__23949),
            .I(N__23926));
    InMux I__4611 (
            .O(N__23948),
            .I(N__23923));
    InMux I__4610 (
            .O(N__23947),
            .I(N__23916));
    InMux I__4609 (
            .O(N__23946),
            .I(N__23916));
    InMux I__4608 (
            .O(N__23945),
            .I(N__23916));
    InMux I__4607 (
            .O(N__23944),
            .I(N__23913));
    LocalMux I__4606 (
            .O(N__23941),
            .I(N__23910));
    LocalMux I__4605 (
            .O(N__23938),
            .I(N__23905));
    LocalMux I__4604 (
            .O(N__23935),
            .I(N__23905));
    LocalMux I__4603 (
            .O(N__23932),
            .I(N__23900));
    LocalMux I__4602 (
            .O(N__23929),
            .I(N__23897));
    LocalMux I__4601 (
            .O(N__23926),
            .I(N__23894));
    LocalMux I__4600 (
            .O(N__23923),
            .I(N__23888));
    LocalMux I__4599 (
            .O(N__23916),
            .I(N__23885));
    LocalMux I__4598 (
            .O(N__23913),
            .I(N__23879));
    Span4Mux_v I__4597 (
            .O(N__23910),
            .I(N__23874));
    Span4Mux_v I__4596 (
            .O(N__23905),
            .I(N__23874));
    InMux I__4595 (
            .O(N__23904),
            .I(N__23871));
    InMux I__4594 (
            .O(N__23903),
            .I(N__23868));
    Span4Mux_h I__4593 (
            .O(N__23900),
            .I(N__23863));
    Span4Mux_s2_v I__4592 (
            .O(N__23897),
            .I(N__23863));
    Span4Mux_v I__4591 (
            .O(N__23894),
            .I(N__23860));
    InMux I__4590 (
            .O(N__23893),
            .I(N__23857));
    InMux I__4589 (
            .O(N__23892),
            .I(N__23852));
    InMux I__4588 (
            .O(N__23891),
            .I(N__23852));
    Span4Mux_h I__4587 (
            .O(N__23888),
            .I(N__23847));
    Span4Mux_v I__4586 (
            .O(N__23885),
            .I(N__23847));
    InMux I__4585 (
            .O(N__23884),
            .I(N__23840));
    InMux I__4584 (
            .O(N__23883),
            .I(N__23840));
    InMux I__4583 (
            .O(N__23882),
            .I(N__23840));
    Span4Mux_v I__4582 (
            .O(N__23879),
            .I(N__23829));
    Span4Mux_v I__4581 (
            .O(N__23874),
            .I(N__23829));
    LocalMux I__4580 (
            .O(N__23871),
            .I(N__23829));
    LocalMux I__4579 (
            .O(N__23868),
            .I(N__23829));
    Span4Mux_v I__4578 (
            .O(N__23863),
            .I(N__23829));
    Odrv4 I__4577 (
            .O(N__23860),
            .I(\POWERLED.N_209 ));
    LocalMux I__4576 (
            .O(N__23857),
            .I(\POWERLED.N_209 ));
    LocalMux I__4575 (
            .O(N__23852),
            .I(\POWERLED.N_209 ));
    Odrv4 I__4574 (
            .O(N__23847),
            .I(\POWERLED.N_209 ));
    LocalMux I__4573 (
            .O(N__23840),
            .I(\POWERLED.N_209 ));
    Odrv4 I__4572 (
            .O(N__23829),
            .I(\POWERLED.N_209 ));
    CascadeMux I__4571 (
            .O(N__23816),
            .I(\POWERLED.N_145_N_cascade_ ));
    InMux I__4570 (
            .O(N__23813),
            .I(N__23801));
    InMux I__4569 (
            .O(N__23812),
            .I(N__23798));
    InMux I__4568 (
            .O(N__23811),
            .I(N__23793));
    InMux I__4567 (
            .O(N__23810),
            .I(N__23793));
    InMux I__4566 (
            .O(N__23809),
            .I(N__23790));
    InMux I__4565 (
            .O(N__23808),
            .I(N__23784));
    InMux I__4564 (
            .O(N__23807),
            .I(N__23784));
    IoInMux I__4563 (
            .O(N__23806),
            .I(N__23781));
    InMux I__4562 (
            .O(N__23805),
            .I(N__23772));
    InMux I__4561 (
            .O(N__23804),
            .I(N__23772));
    LocalMux I__4560 (
            .O(N__23801),
            .I(N__23765));
    LocalMux I__4559 (
            .O(N__23798),
            .I(N__23765));
    LocalMux I__4558 (
            .O(N__23793),
            .I(N__23765));
    LocalMux I__4557 (
            .O(N__23790),
            .I(N__23762));
    CascadeMux I__4556 (
            .O(N__23789),
            .I(N__23759));
    LocalMux I__4555 (
            .O(N__23784),
            .I(N__23752));
    LocalMux I__4554 (
            .O(N__23781),
            .I(N__23752));
    InMux I__4553 (
            .O(N__23780),
            .I(N__23743));
    InMux I__4552 (
            .O(N__23779),
            .I(N__23743));
    InMux I__4551 (
            .O(N__23778),
            .I(N__23743));
    InMux I__4550 (
            .O(N__23777),
            .I(N__23743));
    LocalMux I__4549 (
            .O(N__23772),
            .I(N__23734));
    Span4Mux_s3_v I__4548 (
            .O(N__23765),
            .I(N__23729));
    Span4Mux_s3_v I__4547 (
            .O(N__23762),
            .I(N__23729));
    InMux I__4546 (
            .O(N__23759),
            .I(N__23722));
    InMux I__4545 (
            .O(N__23758),
            .I(N__23722));
    InMux I__4544 (
            .O(N__23757),
            .I(N__23722));
    Span4Mux_s3_h I__4543 (
            .O(N__23752),
            .I(N__23717));
    LocalMux I__4542 (
            .O(N__23743),
            .I(N__23717));
    InMux I__4541 (
            .O(N__23742),
            .I(N__23712));
    InMux I__4540 (
            .O(N__23741),
            .I(N__23712));
    InMux I__4539 (
            .O(N__23740),
            .I(N__23707));
    InMux I__4538 (
            .O(N__23739),
            .I(N__23707));
    CascadeMux I__4537 (
            .O(N__23738),
            .I(N__23704));
    InMux I__4536 (
            .O(N__23737),
            .I(N__23700));
    Span4Mux_v I__4535 (
            .O(N__23734),
            .I(N__23696));
    Span4Mux_v I__4534 (
            .O(N__23729),
            .I(N__23688));
    LocalMux I__4533 (
            .O(N__23722),
            .I(N__23688));
    Span4Mux_h I__4532 (
            .O(N__23717),
            .I(N__23688));
    LocalMux I__4531 (
            .O(N__23712),
            .I(N__23683));
    LocalMux I__4530 (
            .O(N__23707),
            .I(N__23683));
    InMux I__4529 (
            .O(N__23704),
            .I(N__23678));
    InMux I__4528 (
            .O(N__23703),
            .I(N__23678));
    LocalMux I__4527 (
            .O(N__23700),
            .I(N__23675));
    CascadeMux I__4526 (
            .O(N__23699),
            .I(N__23672));
    Span4Mux_v I__4525 (
            .O(N__23696),
            .I(N__23669));
    InMux I__4524 (
            .O(N__23695),
            .I(N__23666));
    Span4Mux_v I__4523 (
            .O(N__23688),
            .I(N__23663));
    Sp12to4 I__4522 (
            .O(N__23683),
            .I(N__23656));
    LocalMux I__4521 (
            .O(N__23678),
            .I(N__23656));
    Span12Mux_s3_v I__4520 (
            .O(N__23675),
            .I(N__23656));
    InMux I__4519 (
            .O(N__23672),
            .I(N__23653));
    Odrv4 I__4518 (
            .O(N__23669),
            .I(G_154));
    LocalMux I__4517 (
            .O(N__23666),
            .I(G_154));
    Odrv4 I__4516 (
            .O(N__23663),
            .I(G_154));
    Odrv12 I__4515 (
            .O(N__23656),
            .I(G_154));
    LocalMux I__4514 (
            .O(N__23653),
            .I(G_154));
    InMux I__4513 (
            .O(N__23642),
            .I(N__23639));
    LocalMux I__4512 (
            .O(N__23639),
            .I(N__23636));
    Span4Mux_h I__4511 (
            .O(N__23636),
            .I(N__23632));
    InMux I__4510 (
            .O(N__23635),
            .I(N__23629));
    Odrv4 I__4509 (
            .O(N__23632),
            .I(\POWERLED.dutycycle_en_9 ));
    LocalMux I__4508 (
            .O(N__23629),
            .I(\POWERLED.dutycycle_en_9 ));
    CascadeMux I__4507 (
            .O(N__23624),
            .I(N__23621));
    InMux I__4506 (
            .O(N__23621),
            .I(N__23617));
    InMux I__4505 (
            .O(N__23620),
            .I(N__23614));
    LocalMux I__4504 (
            .O(N__23617),
            .I(\HDA_STRAP.countZ0Z_0 ));
    LocalMux I__4503 (
            .O(N__23614),
            .I(\HDA_STRAP.countZ0Z_0 ));
    CascadeMux I__4502 (
            .O(N__23609),
            .I(N__23605));
    InMux I__4501 (
            .O(N__23608),
            .I(N__23602));
    InMux I__4500 (
            .O(N__23605),
            .I(N__23599));
    LocalMux I__4499 (
            .O(N__23602),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_1 ));
    LocalMux I__4498 (
            .O(N__23599),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_1 ));
    InMux I__4497 (
            .O(N__23594),
            .I(N__23591));
    LocalMux I__4496 (
            .O(N__23591),
            .I(\HDA_STRAP.count_RNO_0Z0Z_0 ));
    InMux I__4495 (
            .O(N__23588),
            .I(N__23584));
    InMux I__4494 (
            .O(N__23587),
            .I(N__23581));
    LocalMux I__4493 (
            .O(N__23584),
            .I(\HDA_STRAP.countZ0Z_1 ));
    LocalMux I__4492 (
            .O(N__23581),
            .I(\HDA_STRAP.countZ0Z_1 ));
    InMux I__4491 (
            .O(N__23576),
            .I(\HDA_STRAP.un1_count_1_cry_0 ));
    CascadeMux I__4490 (
            .O(N__23573),
            .I(N__23570));
    InMux I__4489 (
            .O(N__23570),
            .I(N__23566));
    InMux I__4488 (
            .O(N__23569),
            .I(N__23563));
    LocalMux I__4487 (
            .O(N__23566),
            .I(\HDA_STRAP.countZ0Z_2 ));
    LocalMux I__4486 (
            .O(N__23563),
            .I(\HDA_STRAP.countZ0Z_2 ));
    InMux I__4485 (
            .O(N__23558),
            .I(\HDA_STRAP.un1_count_1_cry_1 ));
    InMux I__4484 (
            .O(N__23555),
            .I(N__23551));
    InMux I__4483 (
            .O(N__23554),
            .I(N__23548));
    LocalMux I__4482 (
            .O(N__23551),
            .I(\HDA_STRAP.countZ0Z_3 ));
    LocalMux I__4481 (
            .O(N__23548),
            .I(\HDA_STRAP.countZ0Z_3 ));
    InMux I__4480 (
            .O(N__23543),
            .I(\HDA_STRAP.un1_count_1_cry_2 ));
    InMux I__4479 (
            .O(N__23540),
            .I(N__23536));
    InMux I__4478 (
            .O(N__23539),
            .I(N__23533));
    LocalMux I__4477 (
            .O(N__23536),
            .I(\HDA_STRAP.countZ0Z_4 ));
    LocalMux I__4476 (
            .O(N__23533),
            .I(\HDA_STRAP.countZ0Z_4 ));
    CascadeMux I__4475 (
            .O(N__23528),
            .I(\POWERLED.count_clk_RNIBVNSZ0Z_4_cascade_ ));
    CascadeMux I__4474 (
            .O(N__23525),
            .I(N__23522));
    InMux I__4473 (
            .O(N__23522),
            .I(N__23516));
    InMux I__4472 (
            .O(N__23521),
            .I(N__23516));
    LocalMux I__4471 (
            .O(N__23516),
            .I(\POWERLED.dutycycle_eena_2 ));
    InMux I__4470 (
            .O(N__23513),
            .I(N__23509));
    CascadeMux I__4469 (
            .O(N__23512),
            .I(N__23506));
    LocalMux I__4468 (
            .O(N__23509),
            .I(N__23503));
    InMux I__4467 (
            .O(N__23506),
            .I(N__23500));
    Span4Mux_v I__4466 (
            .O(N__23503),
            .I(N__23497));
    LocalMux I__4465 (
            .O(N__23500),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    Odrv4 I__4464 (
            .O(N__23497),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    InMux I__4463 (
            .O(N__23492),
            .I(N__23489));
    LocalMux I__4462 (
            .O(N__23489),
            .I(N__23485));
    CascadeMux I__4461 (
            .O(N__23488),
            .I(N__23482));
    Span4Mux_h I__4460 (
            .O(N__23485),
            .I(N__23479));
    InMux I__4459 (
            .O(N__23482),
            .I(N__23476));
    Odrv4 I__4458 (
            .O(N__23479),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ));
    LocalMux I__4457 (
            .O(N__23476),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ));
    InMux I__4456 (
            .O(N__23471),
            .I(N__23462));
    InMux I__4455 (
            .O(N__23470),
            .I(N__23457));
    InMux I__4454 (
            .O(N__23469),
            .I(N__23457));
    InMux I__4453 (
            .O(N__23468),
            .I(N__23454));
    InMux I__4452 (
            .O(N__23467),
            .I(N__23450));
    CascadeMux I__4451 (
            .O(N__23466),
            .I(N__23446));
    CascadeMux I__4450 (
            .O(N__23465),
            .I(N__23443));
    LocalMux I__4449 (
            .O(N__23462),
            .I(N__23435));
    LocalMux I__4448 (
            .O(N__23457),
            .I(N__23435));
    LocalMux I__4447 (
            .O(N__23454),
            .I(N__23435));
    CascadeMux I__4446 (
            .O(N__23453),
            .I(N__23430));
    LocalMux I__4445 (
            .O(N__23450),
            .I(N__23427));
    InMux I__4444 (
            .O(N__23449),
            .I(N__23422));
    InMux I__4443 (
            .O(N__23446),
            .I(N__23422));
    InMux I__4442 (
            .O(N__23443),
            .I(N__23417));
    InMux I__4441 (
            .O(N__23442),
            .I(N__23417));
    Span4Mux_h I__4440 (
            .O(N__23435),
            .I(N__23414));
    InMux I__4439 (
            .O(N__23434),
            .I(N__23409));
    InMux I__4438 (
            .O(N__23433),
            .I(N__23409));
    InMux I__4437 (
            .O(N__23430),
            .I(N__23406));
    Odrv4 I__4436 (
            .O(N__23427),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4435 (
            .O(N__23422),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4434 (
            .O(N__23417),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__4433 (
            .O(N__23414),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4432 (
            .O(N__23409),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4431 (
            .O(N__23406),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    CascadeMux I__4430 (
            .O(N__23393),
            .I(\POWERLED.dutycycleZ0Z_7_cascade_ ));
    InMux I__4429 (
            .O(N__23390),
            .I(N__23387));
    LocalMux I__4428 (
            .O(N__23387),
            .I(\POWERLED.un1_dutycycle_53_50_3 ));
    InMux I__4427 (
            .O(N__23384),
            .I(N__23381));
    LocalMux I__4426 (
            .O(N__23381),
            .I(N__23375));
    InMux I__4425 (
            .O(N__23380),
            .I(N__23372));
    InMux I__4424 (
            .O(N__23379),
            .I(N__23368));
    CascadeMux I__4423 (
            .O(N__23378),
            .I(N__23363));
    Span4Mux_h I__4422 (
            .O(N__23375),
            .I(N__23358));
    LocalMux I__4421 (
            .O(N__23372),
            .I(N__23358));
    InMux I__4420 (
            .O(N__23371),
            .I(N__23355));
    LocalMux I__4419 (
            .O(N__23368),
            .I(N__23352));
    InMux I__4418 (
            .O(N__23367),
            .I(N__23349));
    InMux I__4417 (
            .O(N__23366),
            .I(N__23344));
    InMux I__4416 (
            .O(N__23363),
            .I(N__23344));
    Odrv4 I__4415 (
            .O(N__23358),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__4414 (
            .O(N__23355),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    Odrv12 I__4413 (
            .O(N__23352),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__4412 (
            .O(N__23349),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__4411 (
            .O(N__23344),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    CascadeMux I__4410 (
            .O(N__23333),
            .I(\POWERLED.un1_dutycycle_53_51_0_cascade_ ));
    InMux I__4409 (
            .O(N__23330),
            .I(N__23327));
    LocalMux I__4408 (
            .O(N__23327),
            .I(N__23324));
    Span4Mux_h I__4407 (
            .O(N__23324),
            .I(N__23321));
    Odrv4 I__4406 (
            .O(N__23321),
            .I(\POWERLED.un1_dutycycle_53_50_4 ));
    InMux I__4405 (
            .O(N__23318),
            .I(N__23315));
    LocalMux I__4404 (
            .O(N__23315),
            .I(N__23312));
    Span4Mux_h I__4403 (
            .O(N__23312),
            .I(N__23309));
    Odrv4 I__4402 (
            .O(N__23309),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_15 ));
    CascadeMux I__4401 (
            .O(N__23306),
            .I(N__23303));
    InMux I__4400 (
            .O(N__23303),
            .I(N__23300));
    LocalMux I__4399 (
            .O(N__23300),
            .I(N__23294));
    InMux I__4398 (
            .O(N__23299),
            .I(N__23289));
    InMux I__4397 (
            .O(N__23298),
            .I(N__23289));
    CascadeMux I__4396 (
            .O(N__23297),
            .I(N__23286));
    Span4Mux_s3_v I__4395 (
            .O(N__23294),
            .I(N__23283));
    LocalMux I__4394 (
            .O(N__23289),
            .I(N__23280));
    InMux I__4393 (
            .O(N__23286),
            .I(N__23277));
    Span4Mux_v I__4392 (
            .O(N__23283),
            .I(N__23274));
    Span4Mux_v I__4391 (
            .O(N__23280),
            .I(N__23269));
    LocalMux I__4390 (
            .O(N__23277),
            .I(N__23269));
    Odrv4 I__4389 (
            .O(N__23274),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_1 ));
    Odrv4 I__4388 (
            .O(N__23269),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_1 ));
    InMux I__4387 (
            .O(N__23264),
            .I(N__23261));
    LocalMux I__4386 (
            .O(N__23261),
            .I(N__23251));
    InMux I__4385 (
            .O(N__23260),
            .I(N__23246));
    InMux I__4384 (
            .O(N__23259),
            .I(N__23237));
    InMux I__4383 (
            .O(N__23258),
            .I(N__23237));
    InMux I__4382 (
            .O(N__23257),
            .I(N__23237));
    InMux I__4381 (
            .O(N__23256),
            .I(N__23232));
    InMux I__4380 (
            .O(N__23255),
            .I(N__23232));
    CascadeMux I__4379 (
            .O(N__23254),
            .I(N__23225));
    Span4Mux_v I__4378 (
            .O(N__23251),
            .I(N__23222));
    InMux I__4377 (
            .O(N__23250),
            .I(N__23217));
    InMux I__4376 (
            .O(N__23249),
            .I(N__23217));
    LocalMux I__4375 (
            .O(N__23246),
            .I(N__23214));
    InMux I__4374 (
            .O(N__23245),
            .I(N__23209));
    InMux I__4373 (
            .O(N__23244),
            .I(N__23209));
    LocalMux I__4372 (
            .O(N__23237),
            .I(N__23204));
    LocalMux I__4371 (
            .O(N__23232),
            .I(N__23204));
    InMux I__4370 (
            .O(N__23231),
            .I(N__23201));
    InMux I__4369 (
            .O(N__23230),
            .I(N__23194));
    InMux I__4368 (
            .O(N__23229),
            .I(N__23194));
    InMux I__4367 (
            .O(N__23228),
            .I(N__23194));
    InMux I__4366 (
            .O(N__23225),
            .I(N__23191));
    Odrv4 I__4365 (
            .O(N__23222),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__4364 (
            .O(N__23217),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__4363 (
            .O(N__23214),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__4362 (
            .O(N__23209),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__4361 (
            .O(N__23204),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__4360 (
            .O(N__23201),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__4359 (
            .O(N__23194),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__4358 (
            .O(N__23191),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    InMux I__4357 (
            .O(N__23174),
            .I(N__23171));
    LocalMux I__4356 (
            .O(N__23171),
            .I(\POWERLED.un1_clk_100khz_30_and_i_o2_0_0_1 ));
    InMux I__4355 (
            .O(N__23168),
            .I(N__23165));
    LocalMux I__4354 (
            .O(N__23165),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_7 ));
    CascadeMux I__4353 (
            .O(N__23162),
            .I(N__23159));
    InMux I__4352 (
            .O(N__23159),
            .I(N__23156));
    LocalMux I__4351 (
            .O(N__23156),
            .I(\POWERLED.N_8_1 ));
    CascadeMux I__4350 (
            .O(N__23153),
            .I(N__23150));
    InMux I__4349 (
            .O(N__23150),
            .I(N__23147));
    LocalMux I__4348 (
            .O(N__23147),
            .I(N__23144));
    Span4Mux_h I__4347 (
            .O(N__23144),
            .I(N__23141));
    Odrv4 I__4346 (
            .O(N__23141),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3 ));
    CascadeMux I__4345 (
            .O(N__23138),
            .I(N__23135));
    InMux I__4344 (
            .O(N__23135),
            .I(N__23121));
    InMux I__4343 (
            .O(N__23134),
            .I(N__23121));
    InMux I__4342 (
            .O(N__23133),
            .I(N__23121));
    InMux I__4341 (
            .O(N__23132),
            .I(N__23112));
    InMux I__4340 (
            .O(N__23131),
            .I(N__23112));
    InMux I__4339 (
            .O(N__23130),
            .I(N__23112));
    CascadeMux I__4338 (
            .O(N__23129),
            .I(N__23109));
    CascadeMux I__4337 (
            .O(N__23128),
            .I(N__23101));
    LocalMux I__4336 (
            .O(N__23121),
            .I(N__23096));
    InMux I__4335 (
            .O(N__23120),
            .I(N__23091));
    InMux I__4334 (
            .O(N__23119),
            .I(N__23091));
    LocalMux I__4333 (
            .O(N__23112),
            .I(N__23088));
    InMux I__4332 (
            .O(N__23109),
            .I(N__23085));
    InMux I__4331 (
            .O(N__23108),
            .I(N__23082));
    InMux I__4330 (
            .O(N__23107),
            .I(N__23073));
    InMux I__4329 (
            .O(N__23106),
            .I(N__23073));
    InMux I__4328 (
            .O(N__23105),
            .I(N__23073));
    InMux I__4327 (
            .O(N__23104),
            .I(N__23073));
    InMux I__4326 (
            .O(N__23101),
            .I(N__23066));
    InMux I__4325 (
            .O(N__23100),
            .I(N__23066));
    InMux I__4324 (
            .O(N__23099),
            .I(N__23066));
    Span4Mux_h I__4323 (
            .O(N__23096),
            .I(N__23057));
    LocalMux I__4322 (
            .O(N__23091),
            .I(N__23057));
    Span4Mux_h I__4321 (
            .O(N__23088),
            .I(N__23057));
    LocalMux I__4320 (
            .O(N__23085),
            .I(N__23057));
    LocalMux I__4319 (
            .O(N__23082),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__4318 (
            .O(N__23073),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__4317 (
            .O(N__23066),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__4316 (
            .O(N__23057),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    CascadeMux I__4315 (
            .O(N__23048),
            .I(\POWERLED.dutycycleZ0Z_9_cascade_ ));
    InMux I__4314 (
            .O(N__23045),
            .I(N__23041));
    CascadeMux I__4313 (
            .O(N__23044),
            .I(N__23037));
    LocalMux I__4312 (
            .O(N__23041),
            .I(N__23031));
    InMux I__4311 (
            .O(N__23040),
            .I(N__23028));
    InMux I__4310 (
            .O(N__23037),
            .I(N__23023));
    InMux I__4309 (
            .O(N__23036),
            .I(N__23023));
    InMux I__4308 (
            .O(N__23035),
            .I(N__23017));
    InMux I__4307 (
            .O(N__23034),
            .I(N__23014));
    Span4Mux_h I__4306 (
            .O(N__23031),
            .I(N__23009));
    LocalMux I__4305 (
            .O(N__23028),
            .I(N__23009));
    LocalMux I__4304 (
            .O(N__23023),
            .I(N__23006));
    InMux I__4303 (
            .O(N__23022),
            .I(N__23001));
    InMux I__4302 (
            .O(N__23021),
            .I(N__23001));
    CascadeMux I__4301 (
            .O(N__23020),
            .I(N__22998));
    LocalMux I__4300 (
            .O(N__23017),
            .I(N__22993));
    LocalMux I__4299 (
            .O(N__23014),
            .I(N__22993));
    Span4Mux_v I__4298 (
            .O(N__23009),
            .I(N__22986));
    Span4Mux_h I__4297 (
            .O(N__23006),
            .I(N__22986));
    LocalMux I__4296 (
            .O(N__23001),
            .I(N__22986));
    InMux I__4295 (
            .O(N__22998),
            .I(N__22983));
    Span4Mux_v I__4294 (
            .O(N__22993),
            .I(N__22980));
    Sp12to4 I__4293 (
            .O(N__22986),
            .I(N__22975));
    LocalMux I__4292 (
            .O(N__22983),
            .I(N__22975));
    Odrv4 I__4291 (
            .O(N__22980),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv12 I__4290 (
            .O(N__22975),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    InMux I__4289 (
            .O(N__22970),
            .I(N__22966));
    InMux I__4288 (
            .O(N__22969),
            .I(N__22963));
    LocalMux I__4287 (
            .O(N__22966),
            .I(N__22960));
    LocalMux I__4286 (
            .O(N__22963),
            .I(N__22957));
    Span4Mux_h I__4285 (
            .O(N__22960),
            .I(N__22954));
    Odrv4 I__4284 (
            .O(N__22957),
            .I(\POWERLED.dutycycle_RNI_11Z0Z_7 ));
    Odrv4 I__4283 (
            .O(N__22954),
            .I(\POWERLED.dutycycle_RNI_11Z0Z_7 ));
    InMux I__4282 (
            .O(N__22949),
            .I(N__22946));
    LocalMux I__4281 (
            .O(N__22946),
            .I(\POWERLED.un1_dutycycle_53_50_a0_1 ));
    CascadeMux I__4280 (
            .O(N__22943),
            .I(\POWERLED.un1_dutycycle_53_2_1_cascade_ ));
    InMux I__4279 (
            .O(N__22940),
            .I(N__22934));
    InMux I__4278 (
            .O(N__22939),
            .I(N__22934));
    LocalMux I__4277 (
            .O(N__22934),
            .I(N__22931));
    Span4Mux_h I__4276 (
            .O(N__22931),
            .I(N__22928));
    Odrv4 I__4275 (
            .O(N__22928),
            .I(\POWERLED.dutycycle_RNIZ0Z_8 ));
    InMux I__4274 (
            .O(N__22925),
            .I(N__22919));
    InMux I__4273 (
            .O(N__22924),
            .I(N__22919));
    LocalMux I__4272 (
            .O(N__22919),
            .I(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ));
    InMux I__4271 (
            .O(N__22916),
            .I(N__22910));
    InMux I__4270 (
            .O(N__22915),
            .I(N__22910));
    LocalMux I__4269 (
            .O(N__22910),
            .I(\POWERLED.dutycycleZ1Z_11 ));
    SRMux I__4268 (
            .O(N__22907),
            .I(N__22897));
    SRMux I__4267 (
            .O(N__22906),
            .I(N__22894));
    SRMux I__4266 (
            .O(N__22905),
            .I(N__22891));
    SRMux I__4265 (
            .O(N__22904),
            .I(N__22888));
    SRMux I__4264 (
            .O(N__22903),
            .I(N__22885));
    SRMux I__4263 (
            .O(N__22902),
            .I(N__22881));
    SRMux I__4262 (
            .O(N__22901),
            .I(N__22875));
    SRMux I__4261 (
            .O(N__22900),
            .I(N__22872));
    LocalMux I__4260 (
            .O(N__22897),
            .I(N__22869));
    LocalMux I__4259 (
            .O(N__22894),
            .I(N__22865));
    LocalMux I__4258 (
            .O(N__22891),
            .I(N__22862));
    LocalMux I__4257 (
            .O(N__22888),
            .I(N__22859));
    LocalMux I__4256 (
            .O(N__22885),
            .I(N__22856));
    SRMux I__4255 (
            .O(N__22884),
            .I(N__22853));
    LocalMux I__4254 (
            .O(N__22881),
            .I(N__22850));
    SRMux I__4253 (
            .O(N__22880),
            .I(N__22847));
    SRMux I__4252 (
            .O(N__22879),
            .I(N__22844));
    SRMux I__4251 (
            .O(N__22878),
            .I(N__22841));
    LocalMux I__4250 (
            .O(N__22875),
            .I(N__22838));
    LocalMux I__4249 (
            .O(N__22872),
            .I(N__22835));
    Span4Mux_s2_v I__4248 (
            .O(N__22869),
            .I(N__22832));
    SRMux I__4247 (
            .O(N__22868),
            .I(N__22829));
    Span4Mux_h I__4246 (
            .O(N__22865),
            .I(N__22824));
    Span4Mux_h I__4245 (
            .O(N__22862),
            .I(N__22824));
    Span4Mux_v I__4244 (
            .O(N__22859),
            .I(N__22821));
    Span4Mux_h I__4243 (
            .O(N__22856),
            .I(N__22818));
    LocalMux I__4242 (
            .O(N__22853),
            .I(N__22813));
    Span4Mux_h I__4241 (
            .O(N__22850),
            .I(N__22813));
    LocalMux I__4240 (
            .O(N__22847),
            .I(N__22810));
    LocalMux I__4239 (
            .O(N__22844),
            .I(N__22807));
    LocalMux I__4238 (
            .O(N__22841),
            .I(N__22804));
    Span4Mux_h I__4237 (
            .O(N__22838),
            .I(N__22801));
    Span4Mux_h I__4236 (
            .O(N__22835),
            .I(N__22798));
    Sp12to4 I__4235 (
            .O(N__22832),
            .I(N__22793));
    LocalMux I__4234 (
            .O(N__22829),
            .I(N__22793));
    Span4Mux_h I__4233 (
            .O(N__22824),
            .I(N__22790));
    Span4Mux_h I__4232 (
            .O(N__22821),
            .I(N__22783));
    Span4Mux_h I__4231 (
            .O(N__22818),
            .I(N__22783));
    Span4Mux_v I__4230 (
            .O(N__22813),
            .I(N__22783));
    Span4Mux_h I__4229 (
            .O(N__22810),
            .I(N__22778));
    Span4Mux_h I__4228 (
            .O(N__22807),
            .I(N__22778));
    Span4Mux_v I__4227 (
            .O(N__22804),
            .I(N__22775));
    Span4Mux_v I__4226 (
            .O(N__22801),
            .I(N__22770));
    Span4Mux_h I__4225 (
            .O(N__22798),
            .I(N__22770));
    Span12Mux_s10_v I__4224 (
            .O(N__22793),
            .I(N__22767));
    Span4Mux_v I__4223 (
            .O(N__22790),
            .I(N__22764));
    Sp12to4 I__4222 (
            .O(N__22783),
            .I(N__22761));
    Span4Mux_v I__4221 (
            .O(N__22778),
            .I(N__22758));
    Odrv4 I__4220 (
            .O(N__22775),
            .I(\POWERLED.N_209_iZ0 ));
    Odrv4 I__4219 (
            .O(N__22770),
            .I(\POWERLED.N_209_iZ0 ));
    Odrv12 I__4218 (
            .O(N__22767),
            .I(\POWERLED.N_209_iZ0 ));
    Odrv4 I__4217 (
            .O(N__22764),
            .I(\POWERLED.N_209_iZ0 ));
    Odrv12 I__4216 (
            .O(N__22761),
            .I(\POWERLED.N_209_iZ0 ));
    Odrv4 I__4215 (
            .O(N__22758),
            .I(\POWERLED.N_209_iZ0 ));
    CascadeMux I__4214 (
            .O(N__22745),
            .I(N__22742));
    InMux I__4213 (
            .O(N__22742),
            .I(N__22738));
    InMux I__4212 (
            .O(N__22741),
            .I(N__22735));
    LocalMux I__4211 (
            .O(N__22738),
            .I(\POWERLED.un1_dutycycle_53_31_a7_0 ));
    LocalMux I__4210 (
            .O(N__22735),
            .I(\POWERLED.un1_dutycycle_53_31_a7_0 ));
    CascadeMux I__4209 (
            .O(N__22730),
            .I(\POWERLED.N_144_N_cascade_ ));
    CascadeMux I__4208 (
            .O(N__22727),
            .I(N__22724));
    InMux I__4207 (
            .O(N__22724),
            .I(N__22721));
    LocalMux I__4206 (
            .O(N__22721),
            .I(N__22717));
    InMux I__4205 (
            .O(N__22720),
            .I(N__22714));
    Odrv4 I__4204 (
            .O(N__22717),
            .I(\POWERLED.dutycycle_en_7 ));
    LocalMux I__4203 (
            .O(N__22714),
            .I(\POWERLED.dutycycle_en_7 ));
    CascadeMux I__4202 (
            .O(N__22709),
            .I(N__22705));
    InMux I__4201 (
            .O(N__22708),
            .I(N__22701));
    InMux I__4200 (
            .O(N__22705),
            .I(N__22696));
    InMux I__4199 (
            .O(N__22704),
            .I(N__22696));
    LocalMux I__4198 (
            .O(N__22701),
            .I(N__22691));
    LocalMux I__4197 (
            .O(N__22696),
            .I(N__22691));
    Odrv4 I__4196 (
            .O(N__22691),
            .I(\POWERLED.dutycycle_eena_3_0_1 ));
    InMux I__4195 (
            .O(N__22688),
            .I(N__22679));
    InMux I__4194 (
            .O(N__22687),
            .I(N__22679));
    InMux I__4193 (
            .O(N__22686),
            .I(N__22679));
    LocalMux I__4192 (
            .O(N__22679),
            .I(N__22676));
    Odrv4 I__4191 (
            .O(N__22676),
            .I(\POWERLED.dutycycle_eena_3_d_0 ));
    InMux I__4190 (
            .O(N__22673),
            .I(N__22669));
    InMux I__4189 (
            .O(N__22672),
            .I(N__22666));
    LocalMux I__4188 (
            .O(N__22669),
            .I(N__22663));
    LocalMux I__4187 (
            .O(N__22666),
            .I(N__22660));
    Span4Mux_s1_v I__4186 (
            .O(N__22663),
            .I(N__22655));
    Span4Mux_h I__4185 (
            .O(N__22660),
            .I(N__22655));
    Odrv4 I__4184 (
            .O(N__22655),
            .I(\POWERLED.dutycycle_en_3 ));
    CascadeMux I__4183 (
            .O(N__22652),
            .I(\POWERLED.un1_dutycycle_53_10_1_0_1_cascade_ ));
    InMux I__4182 (
            .O(N__22649),
            .I(N__22646));
    LocalMux I__4181 (
            .O(N__22646),
            .I(N__22643));
    Odrv12 I__4180 (
            .O(N__22643),
            .I(\POWERLED.un1_dutycycle_53_10_1_0 ));
    InMux I__4179 (
            .O(N__22640),
            .I(N__22637));
    LocalMux I__4178 (
            .O(N__22637),
            .I(N__22634));
    Odrv12 I__4177 (
            .O(N__22634),
            .I(\POWERLED.un2_count_clk_17_0_a2_4 ));
    InMux I__4176 (
            .O(N__22631),
            .I(N__22625));
    InMux I__4175 (
            .O(N__22630),
            .I(N__22625));
    LocalMux I__4174 (
            .O(N__22625),
            .I(N__22622));
    Odrv4 I__4173 (
            .O(N__22622),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    CascadeMux I__4172 (
            .O(N__22619),
            .I(N__22615));
    InMux I__4171 (
            .O(N__22618),
            .I(N__22610));
    InMux I__4170 (
            .O(N__22615),
            .I(N__22610));
    LocalMux I__4169 (
            .O(N__22610),
            .I(\POWERLED.dutycycle_RNI4VJH7Z0Z_4 ));
    CascadeMux I__4168 (
            .O(N__22607),
            .I(N__22604));
    InMux I__4167 (
            .O(N__22604),
            .I(N__22598));
    InMux I__4166 (
            .O(N__22603),
            .I(N__22598));
    LocalMux I__4165 (
            .O(N__22598),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    InMux I__4164 (
            .O(N__22595),
            .I(N__22591));
    InMux I__4163 (
            .O(N__22594),
            .I(N__22588));
    LocalMux I__4162 (
            .O(N__22591),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ));
    LocalMux I__4161 (
            .O(N__22588),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ));
    CascadeMux I__4160 (
            .O(N__22583),
            .I(N__22579));
    CascadeMux I__4159 (
            .O(N__22582),
            .I(N__22576));
    InMux I__4158 (
            .O(N__22579),
            .I(N__22573));
    InMux I__4157 (
            .O(N__22576),
            .I(N__22570));
    LocalMux I__4156 (
            .O(N__22573),
            .I(N__22567));
    LocalMux I__4155 (
            .O(N__22570),
            .I(\POWERLED.dutycycleZ1Z_3 ));
    Odrv4 I__4154 (
            .O(N__22567),
            .I(\POWERLED.dutycycleZ1Z_3 ));
    CascadeMux I__4153 (
            .O(N__22562),
            .I(\POWERLED.dutycycleZ0Z_8_cascade_ ));
    CascadeMux I__4152 (
            .O(N__22559),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_3_cascade_ ));
    InMux I__4151 (
            .O(N__22556),
            .I(N__22550));
    InMux I__4150 (
            .O(N__22555),
            .I(N__22550));
    LocalMux I__4149 (
            .O(N__22550),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_0 ));
    InMux I__4148 (
            .O(N__22547),
            .I(N__22544));
    LocalMux I__4147 (
            .O(N__22544),
            .I(N__22540));
    CascadeMux I__4146 (
            .O(N__22543),
            .I(N__22537));
    Span4Mux_h I__4145 (
            .O(N__22540),
            .I(N__22534));
    InMux I__4144 (
            .O(N__22537),
            .I(N__22531));
    Span4Mux_s3_h I__4143 (
            .O(N__22534),
            .I(N__22528));
    LocalMux I__4142 (
            .O(N__22531),
            .I(N__22525));
    Odrv4 I__4141 (
            .O(N__22528),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_3 ));
    Odrv4 I__4140 (
            .O(N__22525),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_3 ));
    InMux I__4139 (
            .O(N__22520),
            .I(N__22514));
    InMux I__4138 (
            .O(N__22519),
            .I(N__22514));
    LocalMux I__4137 (
            .O(N__22514),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_3 ));
    InMux I__4136 (
            .O(N__22511),
            .I(N__22508));
    LocalMux I__4135 (
            .O(N__22508),
            .I(\POWERLED.un1_dutycycle_53_13_2 ));
    InMux I__4134 (
            .O(N__22505),
            .I(N__22502));
    LocalMux I__4133 (
            .O(N__22502),
            .I(\POWERLED.un1_dutycycle_53_31_4_1 ));
    InMux I__4132 (
            .O(N__22499),
            .I(N__22493));
    InMux I__4131 (
            .O(N__22498),
            .I(N__22493));
    LocalMux I__4130 (
            .O(N__22493),
            .I(\POWERLED.dutycycle_en_8 ));
    CascadeMux I__4129 (
            .O(N__22490),
            .I(N__22486));
    InMux I__4128 (
            .O(N__22489),
            .I(N__22481));
    InMux I__4127 (
            .O(N__22486),
            .I(N__22476));
    InMux I__4126 (
            .O(N__22485),
            .I(N__22476));
    InMux I__4125 (
            .O(N__22484),
            .I(N__22469));
    LocalMux I__4124 (
            .O(N__22481),
            .I(N__22466));
    LocalMux I__4123 (
            .O(N__22476),
            .I(N__22461));
    InMux I__4122 (
            .O(N__22475),
            .I(N__22456));
    InMux I__4121 (
            .O(N__22474),
            .I(N__22456));
    InMux I__4120 (
            .O(N__22473),
            .I(N__22451));
    InMux I__4119 (
            .O(N__22472),
            .I(N__22451));
    LocalMux I__4118 (
            .O(N__22469),
            .I(N__22448));
    Span4Mux_v I__4117 (
            .O(N__22466),
            .I(N__22445));
    InMux I__4116 (
            .O(N__22465),
            .I(N__22440));
    InMux I__4115 (
            .O(N__22464),
            .I(N__22440));
    Span4Mux_h I__4114 (
            .O(N__22461),
            .I(N__22437));
    LocalMux I__4113 (
            .O(N__22456),
            .I(N__22432));
    LocalMux I__4112 (
            .O(N__22451),
            .I(N__22432));
    Span4Mux_v I__4111 (
            .O(N__22448),
            .I(N__22429));
    Sp12to4 I__4110 (
            .O(N__22445),
            .I(N__22424));
    LocalMux I__4109 (
            .O(N__22440),
            .I(N__22424));
    Sp12to4 I__4108 (
            .O(N__22437),
            .I(N__22419));
    Span12Mux_s10_h I__4107 (
            .O(N__22432),
            .I(N__22419));
    Span4Mux_h I__4106 (
            .O(N__22429),
            .I(N__22416));
    Span12Mux_s10_h I__4105 (
            .O(N__22424),
            .I(N__22413));
    Odrv12 I__4104 (
            .O(N__22419),
            .I(slp_s3n));
    Odrv4 I__4103 (
            .O(N__22416),
            .I(slp_s3n));
    Odrv12 I__4102 (
            .O(N__22413),
            .I(slp_s3n));
    IoInMux I__4101 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__4100 (
            .O(N__22403),
            .I(N__22400));
    IoSpan4Mux I__4099 (
            .O(N__22400),
            .I(N__22396));
    InMux I__4098 (
            .O(N__22399),
            .I(N__22393));
    Span4Mux_s0_v I__4097 (
            .O(N__22396),
            .I(N__22388));
    LocalMux I__4096 (
            .O(N__22393),
            .I(N__22381));
    InMux I__4095 (
            .O(N__22392),
            .I(N__22376));
    InMux I__4094 (
            .O(N__22391),
            .I(N__22376));
    Span4Mux_v I__4093 (
            .O(N__22388),
            .I(N__22373));
    InMux I__4092 (
            .O(N__22387),
            .I(N__22370));
    InMux I__4091 (
            .O(N__22386),
            .I(N__22367));
    InMux I__4090 (
            .O(N__22385),
            .I(N__22362));
    InMux I__4089 (
            .O(N__22384),
            .I(N__22362));
    Span4Mux_v I__4088 (
            .O(N__22381),
            .I(N__22359));
    LocalMux I__4087 (
            .O(N__22376),
            .I(N__22356));
    Span4Mux_v I__4086 (
            .O(N__22373),
            .I(N__22351));
    LocalMux I__4085 (
            .O(N__22370),
            .I(N__22351));
    LocalMux I__4084 (
            .O(N__22367),
            .I(N__22346));
    LocalMux I__4083 (
            .O(N__22362),
            .I(N__22346));
    Span4Mux_h I__4082 (
            .O(N__22359),
            .I(N__22341));
    Span4Mux_h I__4081 (
            .O(N__22356),
            .I(N__22341));
    Odrv4 I__4080 (
            .O(N__22351),
            .I(rsmrstn));
    Odrv12 I__4079 (
            .O(N__22346),
            .I(rsmrstn));
    Odrv4 I__4078 (
            .O(N__22341),
            .I(rsmrstn));
    InMux I__4077 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__4076 (
            .O(N__22331),
            .I(\POWERLED.N_222 ));
    InMux I__4075 (
            .O(N__22328),
            .I(N__22325));
    LocalMux I__4074 (
            .O(N__22325),
            .I(\POWERLED.un1_dutycycle_172_sm3 ));
    InMux I__4073 (
            .O(N__22322),
            .I(N__22319));
    LocalMux I__4072 (
            .O(N__22319),
            .I(\POWERLED.un1_clk_100khz_52_and_i_m2_1 ));
    CascadeMux I__4071 (
            .O(N__22316),
            .I(\POWERLED.un1_dutycycle_172_m4_cascade_ ));
    InMux I__4070 (
            .O(N__22313),
            .I(N__22310));
    LocalMux I__4069 (
            .O(N__22310),
            .I(N__22307));
    Odrv12 I__4068 (
            .O(N__22307),
            .I(\POWERLED.un1_clk_100khz_52_and_i_0Z0Z_0 ));
    CascadeMux I__4067 (
            .O(N__22304),
            .I(\POWERLED.N_225_cascade_ ));
    CascadeMux I__4066 (
            .O(N__22301),
            .I(\POWERLED.dutycycle_eena_14_cascade_ ));
    InMux I__4065 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__4064 (
            .O(N__22295),
            .I(N__22292));
    Span4Mux_h I__4063 (
            .O(N__22292),
            .I(N__22289));
    Odrv4 I__4062 (
            .O(N__22289),
            .I(\POWERLED.dutycycle_eena_14 ));
    InMux I__4061 (
            .O(N__22286),
            .I(N__22280));
    InMux I__4060 (
            .O(N__22285),
            .I(N__22280));
    LocalMux I__4059 (
            .O(N__22280),
            .I(N__22277));
    Span4Mux_v I__4058 (
            .O(N__22277),
            .I(N__22274));
    Odrv4 I__4057 (
            .O(N__22274),
            .I(\POWERLED.dutycycle_set_1 ));
    InMux I__4056 (
            .O(N__22271),
            .I(N__22265));
    InMux I__4055 (
            .O(N__22270),
            .I(N__22265));
    LocalMux I__4054 (
            .O(N__22265),
            .I(\POWERLED.dutycycle_0_5 ));
    InMux I__4053 (
            .O(N__22262),
            .I(N__22259));
    LocalMux I__4052 (
            .O(N__22259),
            .I(\POWERLED.count_clk_0_3 ));
    InMux I__4051 (
            .O(N__22256),
            .I(N__22253));
    LocalMux I__4050 (
            .O(N__22253),
            .I(\POWERLED.count_clk_0_4 ));
    CascadeMux I__4049 (
            .O(N__22250),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_5_cascade_ ));
    CascadeMux I__4048 (
            .O(N__22247),
            .I(N__22239));
    InMux I__4047 (
            .O(N__22246),
            .I(N__22234));
    InMux I__4046 (
            .O(N__22245),
            .I(N__22234));
    InMux I__4045 (
            .O(N__22244),
            .I(N__22231));
    InMux I__4044 (
            .O(N__22243),
            .I(N__22223));
    InMux I__4043 (
            .O(N__22242),
            .I(N__22223));
    InMux I__4042 (
            .O(N__22239),
            .I(N__22223));
    LocalMux I__4041 (
            .O(N__22234),
            .I(N__22216));
    LocalMux I__4040 (
            .O(N__22231),
            .I(N__22216));
    InMux I__4039 (
            .O(N__22230),
            .I(N__22213));
    LocalMux I__4038 (
            .O(N__22223),
            .I(N__22210));
    InMux I__4037 (
            .O(N__22222),
            .I(N__22207));
    InMux I__4036 (
            .O(N__22221),
            .I(N__22204));
    Span4Mux_v I__4035 (
            .O(N__22216),
            .I(N__22201));
    LocalMux I__4034 (
            .O(N__22213),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__4033 (
            .O(N__22210),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__4032 (
            .O(N__22207),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__4031 (
            .O(N__22204),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__4030 (
            .O(N__22201),
            .I(\POWERLED.func_stateZ0Z_0 ));
    InMux I__4029 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__4028 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_v I__4027 (
            .O(N__22184),
            .I(N__22180));
    InMux I__4026 (
            .O(N__22183),
            .I(N__22177));
    Odrv4 I__4025 (
            .O(N__22180),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_0 ));
    LocalMux I__4024 (
            .O(N__22177),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_0 ));
    CascadeMux I__4023 (
            .O(N__22172),
            .I(N__22166));
    InMux I__4022 (
            .O(N__22171),
            .I(N__22161));
    InMux I__4021 (
            .O(N__22170),
            .I(N__22161));
    CascadeMux I__4020 (
            .O(N__22169),
            .I(N__22158));
    InMux I__4019 (
            .O(N__22166),
            .I(N__22155));
    LocalMux I__4018 (
            .O(N__22161),
            .I(N__22152));
    InMux I__4017 (
            .O(N__22158),
            .I(N__22149));
    LocalMux I__4016 (
            .O(N__22155),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_0 ));
    Odrv12 I__4015 (
            .O(N__22152),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_0 ));
    LocalMux I__4014 (
            .O(N__22149),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_0 ));
    CascadeMux I__4013 (
            .O(N__22142),
            .I(N__22137));
    InMux I__4012 (
            .O(N__22141),
            .I(N__22133));
    InMux I__4011 (
            .O(N__22140),
            .I(N__22128));
    InMux I__4010 (
            .O(N__22137),
            .I(N__22123));
    InMux I__4009 (
            .O(N__22136),
            .I(N__22123));
    LocalMux I__4008 (
            .O(N__22133),
            .I(N__22119));
    InMux I__4007 (
            .O(N__22132),
            .I(N__22114));
    InMux I__4006 (
            .O(N__22131),
            .I(N__22114));
    LocalMux I__4005 (
            .O(N__22128),
            .I(N__22111));
    LocalMux I__4004 (
            .O(N__22123),
            .I(N__22108));
    InMux I__4003 (
            .O(N__22122),
            .I(N__22105));
    Span4Mux_v I__4002 (
            .O(N__22119),
            .I(N__22100));
    LocalMux I__4001 (
            .O(N__22114),
            .I(N__22100));
    Span4Mux_h I__4000 (
            .O(N__22111),
            .I(N__22097));
    Span4Mux_v I__3999 (
            .O(N__22108),
            .I(N__22092));
    LocalMux I__3998 (
            .O(N__22105),
            .I(N__22092));
    Span4Mux_v I__3997 (
            .O(N__22100),
            .I(N__22089));
    Span4Mux_v I__3996 (
            .O(N__22097),
            .I(N__22086));
    Span4Mux_v I__3995 (
            .O(N__22092),
            .I(N__22083));
    Odrv4 I__3994 (
            .O(N__22089),
            .I(\POWERLED.N_337 ));
    Odrv4 I__3993 (
            .O(N__22086),
            .I(\POWERLED.N_337 ));
    Odrv4 I__3992 (
            .O(N__22083),
            .I(\POWERLED.N_337 ));
    InMux I__3991 (
            .O(N__22076),
            .I(N__22073));
    LocalMux I__3990 (
            .O(N__22073),
            .I(N__22069));
    InMux I__3989 (
            .O(N__22072),
            .I(N__22065));
    Span4Mux_h I__3988 (
            .O(N__22069),
            .I(N__22062));
    InMux I__3987 (
            .O(N__22068),
            .I(N__22059));
    LocalMux I__3986 (
            .O(N__22065),
            .I(SUSWARN_N_fast));
    Odrv4 I__3985 (
            .O(N__22062),
            .I(SUSWARN_N_fast));
    LocalMux I__3984 (
            .O(N__22059),
            .I(SUSWARN_N_fast));
    CascadeMux I__3983 (
            .O(N__22052),
            .I(\POWERLED.N_390_cascade_ ));
    CascadeMux I__3982 (
            .O(N__22049),
            .I(N__22045));
    InMux I__3981 (
            .O(N__22048),
            .I(N__22042));
    InMux I__3980 (
            .O(N__22045),
            .I(N__22037));
    LocalMux I__3979 (
            .O(N__22042),
            .I(N__22034));
    InMux I__3978 (
            .O(N__22041),
            .I(N__22031));
    CascadeMux I__3977 (
            .O(N__22040),
            .I(N__22026));
    LocalMux I__3976 (
            .O(N__22037),
            .I(N__22023));
    Sp12to4 I__3975 (
            .O(N__22034),
            .I(N__22018));
    LocalMux I__3974 (
            .O(N__22031),
            .I(N__22018));
    InMux I__3973 (
            .O(N__22030),
            .I(N__22015));
    InMux I__3972 (
            .O(N__22029),
            .I(N__22010));
    InMux I__3971 (
            .O(N__22026),
            .I(N__22010));
    Odrv4 I__3970 (
            .O(N__22023),
            .I(SUSWARN_N_rep1));
    Odrv12 I__3969 (
            .O(N__22018),
            .I(SUSWARN_N_rep1));
    LocalMux I__3968 (
            .O(N__22015),
            .I(SUSWARN_N_rep1));
    LocalMux I__3967 (
            .O(N__22010),
            .I(SUSWARN_N_rep1));
    CascadeMux I__3966 (
            .O(N__22001),
            .I(\POWERLED.dutycycle_eena_3_0_0_sx_cascade_ ));
    InMux I__3965 (
            .O(N__21998),
            .I(N__21995));
    LocalMux I__3964 (
            .O(N__21995),
            .I(N__21991));
    InMux I__3963 (
            .O(N__21994),
            .I(N__21987));
    Span4Mux_v I__3962 (
            .O(N__21991),
            .I(N__21984));
    InMux I__3961 (
            .O(N__21990),
            .I(N__21981));
    LocalMux I__3960 (
            .O(N__21987),
            .I(N__21978));
    Span4Mux_h I__3959 (
            .O(N__21984),
            .I(N__21973));
    LocalMux I__3958 (
            .O(N__21981),
            .I(N__21973));
    Span4Mux_h I__3957 (
            .O(N__21978),
            .I(N__21970));
    Odrv4 I__3956 (
            .O(N__21973),
            .I(\POWERLED.countZ0Z_12 ));
    Odrv4 I__3955 (
            .O(N__21970),
            .I(\POWERLED.countZ0Z_12 ));
    CascadeMux I__3954 (
            .O(N__21965),
            .I(N__21962));
    InMux I__3953 (
            .O(N__21962),
            .I(N__21956));
    InMux I__3952 (
            .O(N__21961),
            .I(N__21956));
    LocalMux I__3951 (
            .O(N__21956),
            .I(N__21953));
    Odrv4 I__3950 (
            .O(N__21953),
            .I(\POWERLED.un1_count_cry_11_c_RNISEHZ0Z7 ));
    InMux I__3949 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__3948 (
            .O(N__21947),
            .I(\POWERLED.count_0_12 ));
    InMux I__3947 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__3946 (
            .O(N__21941),
            .I(\POWERLED.count_clk_0_2 ));
    InMux I__3945 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__3944 (
            .O(N__21935),
            .I(\POWERLED.count_clk_0_13 ));
    InMux I__3943 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__3942 (
            .O(N__21929),
            .I(N__21926));
    Odrv4 I__3941 (
            .O(N__21926),
            .I(\POWERLED.count_clk_0_14 ));
    CascadeMux I__3940 (
            .O(N__21923),
            .I(\POWERLED.un1_clk_100khz_48_and_i_o2_2_0_cascade_ ));
    InMux I__3939 (
            .O(N__21920),
            .I(N__21917));
    LocalMux I__3938 (
            .O(N__21917),
            .I(\POWERLED.un1_clk_100khz_48_and_i_o2_3_0 ));
    InMux I__3937 (
            .O(N__21914),
            .I(N__21910));
    InMux I__3936 (
            .O(N__21913),
            .I(N__21907));
    LocalMux I__3935 (
            .O(N__21910),
            .I(\POWERLED.N_197 ));
    LocalMux I__3934 (
            .O(N__21907),
            .I(\POWERLED.N_197 ));
    CascadeMux I__3933 (
            .O(N__21902),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ));
    InMux I__3932 (
            .O(N__21899),
            .I(N__21896));
    LocalMux I__3931 (
            .O(N__21896),
            .I(N__21893));
    Span4Mux_h I__3930 (
            .O(N__21893),
            .I(N__21888));
    CascadeMux I__3929 (
            .O(N__21892),
            .I(N__21885));
    CascadeMux I__3928 (
            .O(N__21891),
            .I(N__21882));
    Span4Mux_v I__3927 (
            .O(N__21888),
            .I(N__21877));
    InMux I__3926 (
            .O(N__21885),
            .I(N__21874));
    InMux I__3925 (
            .O(N__21882),
            .I(N__21871));
    InMux I__3924 (
            .O(N__21881),
            .I(N__21868));
    InMux I__3923 (
            .O(N__21880),
            .I(N__21865));
    Span4Mux_v I__3922 (
            .O(N__21877),
            .I(N__21862));
    LocalMux I__3921 (
            .O(N__21874),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__3920 (
            .O(N__21871),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__3919 (
            .O(N__21868),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__3918 (
            .O(N__21865),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    Odrv4 I__3917 (
            .O(N__21862),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    CascadeMux I__3916 (
            .O(N__21851),
            .I(N__21848));
    InMux I__3915 (
            .O(N__21848),
            .I(N__21845));
    LocalMux I__3914 (
            .O(N__21845),
            .I(N__21842));
    Span4Mux_v I__3913 (
            .O(N__21842),
            .I(N__21839));
    Span4Mux_h I__3912 (
            .O(N__21839),
            .I(N__21836));
    Odrv4 I__3911 (
            .O(N__21836),
            .I(\POWERLED.un85_clk_100khz_10 ));
    InMux I__3910 (
            .O(N__21833),
            .I(N__21830));
    LocalMux I__3909 (
            .O(N__21830),
            .I(\POWERLED.un1_func_state25_6_0_o_N_287_N ));
    InMux I__3908 (
            .O(N__21827),
            .I(N__21824));
    LocalMux I__3907 (
            .O(N__21824),
            .I(\POWERLED.func_state_RNI_1Z0Z_0 ));
    CascadeMux I__3906 (
            .O(N__21821),
            .I(\POWERLED.func_state_RNI_1Z0Z_0_cascade_ ));
    CascadeMux I__3905 (
            .O(N__21818),
            .I(N__21815));
    InMux I__3904 (
            .O(N__21815),
            .I(N__21812));
    LocalMux I__3903 (
            .O(N__21812),
            .I(N__21807));
    InMux I__3902 (
            .O(N__21811),
            .I(N__21804));
    InMux I__3901 (
            .O(N__21810),
            .I(N__21801));
    Odrv12 I__3900 (
            .O(N__21807),
            .I(\POWERLED.func_state_RNIBK1UZ0Z_0 ));
    LocalMux I__3899 (
            .O(N__21804),
            .I(\POWERLED.func_state_RNIBK1UZ0Z_0 ));
    LocalMux I__3898 (
            .O(N__21801),
            .I(\POWERLED.func_state_RNIBK1UZ0Z_0 ));
    CascadeMux I__3897 (
            .O(N__21794),
            .I(N__21790));
    CascadeMux I__3896 (
            .O(N__21793),
            .I(N__21787));
    InMux I__3895 (
            .O(N__21790),
            .I(N__21783));
    InMux I__3894 (
            .O(N__21787),
            .I(N__21780));
    CascadeMux I__3893 (
            .O(N__21786),
            .I(N__21777));
    LocalMux I__3892 (
            .O(N__21783),
            .I(N__21772));
    LocalMux I__3891 (
            .O(N__21780),
            .I(N__21769));
    InMux I__3890 (
            .O(N__21777),
            .I(N__21764));
    InMux I__3889 (
            .O(N__21776),
            .I(N__21764));
    InMux I__3888 (
            .O(N__21775),
            .I(N__21760));
    Span4Mux_v I__3887 (
            .O(N__21772),
            .I(N__21755));
    Span4Mux_v I__3886 (
            .O(N__21769),
            .I(N__21755));
    LocalMux I__3885 (
            .O(N__21764),
            .I(N__21752));
    InMux I__3884 (
            .O(N__21763),
            .I(N__21748));
    LocalMux I__3883 (
            .O(N__21760),
            .I(N__21745));
    Span4Mux_h I__3882 (
            .O(N__21755),
            .I(N__21740));
    Span4Mux_v I__3881 (
            .O(N__21752),
            .I(N__21740));
    InMux I__3880 (
            .O(N__21751),
            .I(N__21737));
    LocalMux I__3879 (
            .O(N__21748),
            .I(\POWERLED.N_326_0 ));
    Odrv12 I__3878 (
            .O(N__21745),
            .I(\POWERLED.N_326_0 ));
    Odrv4 I__3877 (
            .O(N__21740),
            .I(\POWERLED.N_326_0 ));
    LocalMux I__3876 (
            .O(N__21737),
            .I(\POWERLED.N_326_0 ));
    InMux I__3875 (
            .O(N__21728),
            .I(N__21725));
    LocalMux I__3874 (
            .O(N__21725),
            .I(N__21722));
    Span4Mux_h I__3873 (
            .O(N__21722),
            .I(N__21718));
    InMux I__3872 (
            .O(N__21721),
            .I(N__21715));
    Span4Mux_h I__3871 (
            .O(N__21718),
            .I(N__21712));
    LocalMux I__3870 (
            .O(N__21715),
            .I(\POWERLED.func_stateZ1Z_0 ));
    Odrv4 I__3869 (
            .O(N__21712),
            .I(\POWERLED.func_stateZ1Z_0 ));
    InMux I__3868 (
            .O(N__21707),
            .I(N__21704));
    LocalMux I__3867 (
            .O(N__21704),
            .I(N__21701));
    Span4Mux_v I__3866 (
            .O(N__21701),
            .I(N__21698));
    Span4Mux_h I__3865 (
            .O(N__21698),
            .I(N__21695));
    Span4Mux_h I__3864 (
            .O(N__21695),
            .I(N__21691));
    InMux I__3863 (
            .O(N__21694),
            .I(N__21688));
    Odrv4 I__3862 (
            .O(N__21691),
            .I(\POWERLED.func_state_RNIB74H7Z0Z_1 ));
    LocalMux I__3861 (
            .O(N__21688),
            .I(\POWERLED.func_state_RNIB74H7Z0Z_1 ));
    InMux I__3860 (
            .O(N__21683),
            .I(N__21680));
    LocalMux I__3859 (
            .O(N__21680),
            .I(N__21677));
    Odrv12 I__3858 (
            .O(N__21677),
            .I(\POWERLED.func_state_RNI6RANZ0Z_1 ));
    CascadeMux I__3857 (
            .O(N__21674),
            .I(\POWERLED.func_stateZ0Z_0_cascade_ ));
    InMux I__3856 (
            .O(N__21671),
            .I(N__21668));
    LocalMux I__3855 (
            .O(N__21668),
            .I(N__21665));
    Span4Mux_v I__3854 (
            .O(N__21665),
            .I(N__21662));
    Odrv4 I__3853 (
            .O(N__21662),
            .I(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ));
    CascadeMux I__3852 (
            .O(N__21659),
            .I(\POWERLED.N_275_cascade_ ));
    CascadeMux I__3851 (
            .O(N__21656),
            .I(\POWERLED.count_off_RNIZ0Z_11_cascade_ ));
    InMux I__3850 (
            .O(N__21653),
            .I(N__21650));
    LocalMux I__3849 (
            .O(N__21650),
            .I(\POWERLED.N_310 ));
    CascadeMux I__3848 (
            .O(N__21647),
            .I(\POWERLED.N_314_cascade_ ));
    CascadeMux I__3847 (
            .O(N__21644),
            .I(N__21641));
    InMux I__3846 (
            .O(N__21641),
            .I(N__21636));
    InMux I__3845 (
            .O(N__21640),
            .I(N__21631));
    InMux I__3844 (
            .O(N__21639),
            .I(N__21631));
    LocalMux I__3843 (
            .O(N__21636),
            .I(N__21624));
    LocalMux I__3842 (
            .O(N__21631),
            .I(N__21624));
    InMux I__3841 (
            .O(N__21630),
            .I(N__21621));
    InMux I__3840 (
            .O(N__21629),
            .I(N__21618));
    Odrv4 I__3839 (
            .O(N__21624),
            .I(\POWERLED.count_off_RNIZ0Z_11 ));
    LocalMux I__3838 (
            .O(N__21621),
            .I(\POWERLED.count_off_RNIZ0Z_11 ));
    LocalMux I__3837 (
            .O(N__21618),
            .I(\POWERLED.count_off_RNIZ0Z_11 ));
    CascadeMux I__3836 (
            .O(N__21611),
            .I(\POWERLED.func_state_1_ss0_i_0_o2_1_cascade_ ));
    InMux I__3835 (
            .O(N__21608),
            .I(N__21605));
    LocalMux I__3834 (
            .O(N__21605),
            .I(\POWERLED.func_state_RNIHDGK3_0Z0Z_1 ));
    InMux I__3833 (
            .O(N__21602),
            .I(N__21599));
    LocalMux I__3832 (
            .O(N__21599),
            .I(N__21595));
    InMux I__3831 (
            .O(N__21598),
            .I(N__21592));
    Odrv4 I__3830 (
            .O(N__21595),
            .I(\POWERLED.N_67 ));
    LocalMux I__3829 (
            .O(N__21592),
            .I(\POWERLED.N_67 ));
    InMux I__3828 (
            .O(N__21587),
            .I(N__21584));
    LocalMux I__3827 (
            .O(N__21584),
            .I(\POWERLED.func_state_1_m0_0 ));
    CascadeMux I__3826 (
            .O(N__21581),
            .I(\POWERLED.func_state_RNIHDGK3_0Z0Z_1_cascade_ ));
    CascadeMux I__3825 (
            .O(N__21578),
            .I(N__21566));
    InMux I__3824 (
            .O(N__21577),
            .I(N__21548));
    InMux I__3823 (
            .O(N__21576),
            .I(N__21548));
    InMux I__3822 (
            .O(N__21575),
            .I(N__21548));
    InMux I__3821 (
            .O(N__21574),
            .I(N__21548));
    InMux I__3820 (
            .O(N__21573),
            .I(N__21548));
    InMux I__3819 (
            .O(N__21572),
            .I(N__21548));
    InMux I__3818 (
            .O(N__21571),
            .I(N__21548));
    InMux I__3817 (
            .O(N__21570),
            .I(N__21537));
    InMux I__3816 (
            .O(N__21569),
            .I(N__21537));
    InMux I__3815 (
            .O(N__21566),
            .I(N__21537));
    InMux I__3814 (
            .O(N__21565),
            .I(N__21537));
    InMux I__3813 (
            .O(N__21564),
            .I(N__21537));
    InMux I__3812 (
            .O(N__21563),
            .I(N__21534));
    LocalMux I__3811 (
            .O(N__21548),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__3810 (
            .O(N__21537),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__3809 (
            .O(N__21534),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    CascadeMux I__3808 (
            .O(N__21527),
            .I(N__21519));
    CascadeMux I__3807 (
            .O(N__21526),
            .I(N__21515));
    CascadeMux I__3806 (
            .O(N__21525),
            .I(N__21512));
    CascadeMux I__3805 (
            .O(N__21524),
            .I(N__21509));
    CascadeMux I__3804 (
            .O(N__21523),
            .I(N__21500));
    InMux I__3803 (
            .O(N__21522),
            .I(N__21496));
    InMux I__3802 (
            .O(N__21519),
            .I(N__21493));
    InMux I__3801 (
            .O(N__21518),
            .I(N__21480));
    InMux I__3800 (
            .O(N__21515),
            .I(N__21480));
    InMux I__3799 (
            .O(N__21512),
            .I(N__21480));
    InMux I__3798 (
            .O(N__21509),
            .I(N__21480));
    InMux I__3797 (
            .O(N__21508),
            .I(N__21480));
    InMux I__3796 (
            .O(N__21507),
            .I(N__21480));
    InMux I__3795 (
            .O(N__21506),
            .I(N__21473));
    InMux I__3794 (
            .O(N__21505),
            .I(N__21473));
    InMux I__3793 (
            .O(N__21504),
            .I(N__21473));
    InMux I__3792 (
            .O(N__21503),
            .I(N__21466));
    InMux I__3791 (
            .O(N__21500),
            .I(N__21466));
    InMux I__3790 (
            .O(N__21499),
            .I(N__21466));
    LocalMux I__3789 (
            .O(N__21496),
            .I(N__21463));
    LocalMux I__3788 (
            .O(N__21493),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__3787 (
            .O(N__21480),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__3786 (
            .O(N__21473),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__3785 (
            .O(N__21466),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    Odrv4 I__3784 (
            .O(N__21463),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    InMux I__3783 (
            .O(N__21452),
            .I(N__21428));
    InMux I__3782 (
            .O(N__21451),
            .I(N__21428));
    InMux I__3781 (
            .O(N__21450),
            .I(N__21428));
    InMux I__3780 (
            .O(N__21449),
            .I(N__21428));
    InMux I__3779 (
            .O(N__21448),
            .I(N__21428));
    InMux I__3778 (
            .O(N__21447),
            .I(N__21428));
    InMux I__3777 (
            .O(N__21446),
            .I(N__21428));
    InMux I__3776 (
            .O(N__21445),
            .I(N__21421));
    InMux I__3775 (
            .O(N__21444),
            .I(N__21421));
    InMux I__3774 (
            .O(N__21443),
            .I(N__21421));
    LocalMux I__3773 (
            .O(N__21428),
            .I(\HDA_STRAP.un4_count ));
    LocalMux I__3772 (
            .O(N__21421),
            .I(\HDA_STRAP.un4_count ));
    InMux I__3771 (
            .O(N__21416),
            .I(N__21413));
    LocalMux I__3770 (
            .O(N__21413),
            .I(\POWERLED.func_state_1_m2s2_i_0 ));
    CascadeMux I__3769 (
            .O(N__21410),
            .I(\POWERLED.func_state_1_m2s2_i_1_cascade_ ));
    InMux I__3768 (
            .O(N__21407),
            .I(N__21404));
    LocalMux I__3767 (
            .O(N__21404),
            .I(N__21401));
    Span4Mux_s3_v I__3766 (
            .O(N__21401),
            .I(N__21398));
    Odrv4 I__3765 (
            .O(N__21398),
            .I(\POWERLED.func_state_1_m0_0_1_0 ));
    CascadeMux I__3764 (
            .O(N__21395),
            .I(\HDA_STRAP.un4_count_9_cascade_ ));
    InMux I__3763 (
            .O(N__21392),
            .I(N__21389));
    LocalMux I__3762 (
            .O(N__21389),
            .I(\HDA_STRAP.un4_count_13 ));
    InMux I__3761 (
            .O(N__21386),
            .I(N__21383));
    LocalMux I__3760 (
            .O(N__21383),
            .I(\HDA_STRAP.un4_count_11 ));
    InMux I__3759 (
            .O(N__21380),
            .I(N__21377));
    LocalMux I__3758 (
            .O(N__21377),
            .I(\HDA_STRAP.un4_count_10 ));
    CascadeMux I__3757 (
            .O(N__21374),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_0_0_cascade_ ));
    CascadeMux I__3756 (
            .O(N__21371),
            .I(N__21368));
    InMux I__3755 (
            .O(N__21368),
            .I(N__21365));
    LocalMux I__3754 (
            .O(N__21365),
            .I(\POWERLED.dutycycle_RNIEB706Z0Z_7 ));
    InMux I__3753 (
            .O(N__21362),
            .I(N__21356));
    InMux I__3752 (
            .O(N__21361),
            .I(N__21356));
    LocalMux I__3751 (
            .O(N__21356),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    CascadeMux I__3750 (
            .O(N__21353),
            .I(\POWERLED.dutycycle_RNIEB706Z0Z_7_cascade_ ));
    InMux I__3749 (
            .O(N__21350),
            .I(N__21344));
    InMux I__3748 (
            .O(N__21349),
            .I(N__21344));
    LocalMux I__3747 (
            .O(N__21344),
            .I(N__21341));
    Odrv4 I__3746 (
            .O(N__21341),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ));
    CascadeMux I__3745 (
            .O(N__21338),
            .I(\POWERLED.dutycycleZ1Z_6_cascade_ ));
    InMux I__3744 (
            .O(N__21335),
            .I(N__21332));
    LocalMux I__3743 (
            .O(N__21332),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_d_0 ));
    CascadeMux I__3742 (
            .O(N__21329),
            .I(\POWERLED.N_143_N_cascade_ ));
    CascadeMux I__3741 (
            .O(N__21326),
            .I(N__21322));
    InMux I__3740 (
            .O(N__21325),
            .I(N__21317));
    InMux I__3739 (
            .O(N__21322),
            .I(N__21317));
    LocalMux I__3738 (
            .O(N__21317),
            .I(N__21314));
    Span4Mux_h I__3737 (
            .O(N__21314),
            .I(N__21311));
    Odrv4 I__3736 (
            .O(N__21311),
            .I(\POWERLED.dutycycle_en_4 ));
    InMux I__3735 (
            .O(N__21308),
            .I(N__21305));
    LocalMux I__3734 (
            .O(N__21305),
            .I(N__21301));
    InMux I__3733 (
            .O(N__21304),
            .I(N__21298));
    Span4Mux_s1_v I__3732 (
            .O(N__21301),
            .I(N__21293));
    LocalMux I__3731 (
            .O(N__21298),
            .I(N__21293));
    Odrv4 I__3730 (
            .O(N__21293),
            .I(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ));
    CascadeMux I__3729 (
            .O(N__21290),
            .I(N__21287));
    InMux I__3728 (
            .O(N__21287),
            .I(N__21283));
    InMux I__3727 (
            .O(N__21286),
            .I(N__21280));
    LocalMux I__3726 (
            .O(N__21283),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    LocalMux I__3725 (
            .O(N__21280),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    CascadeMux I__3724 (
            .O(N__21275),
            .I(N__21272));
    InMux I__3723 (
            .O(N__21272),
            .I(N__21269));
    LocalMux I__3722 (
            .O(N__21269),
            .I(\HDA_STRAP.un4_count_12 ));
    CascadeMux I__3721 (
            .O(N__21266),
            .I(\POWERLED.g0_i_1_cascade_ ));
    InMux I__3720 (
            .O(N__21263),
            .I(N__21260));
    LocalMux I__3719 (
            .O(N__21260),
            .I(\POWERLED.g0_i_0 ));
    InMux I__3718 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__3717 (
            .O(N__21254),
            .I(N__21251));
    Span4Mux_v I__3716 (
            .O(N__21251),
            .I(N__21248));
    Odrv4 I__3715 (
            .O(N__21248),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_13 ));
    InMux I__3714 (
            .O(N__21245),
            .I(N__21239));
    InMux I__3713 (
            .O(N__21244),
            .I(N__21239));
    LocalMux I__3712 (
            .O(N__21239),
            .I(N__21236));
    Odrv4 I__3711 (
            .O(N__21236),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    CascadeMux I__3710 (
            .O(N__21233),
            .I(N__21229));
    InMux I__3709 (
            .O(N__21232),
            .I(N__21224));
    InMux I__3708 (
            .O(N__21229),
            .I(N__21224));
    LocalMux I__3707 (
            .O(N__21224),
            .I(\POWERLED.dutycycle_rst_1 ));
    CascadeMux I__3706 (
            .O(N__21221),
            .I(\POWERLED.dutycycleZ0Z_4_cascade_ ));
    CascadeMux I__3705 (
            .O(N__21218),
            .I(\POWERLED.g0_1_cascade_ ));
    CascadeMux I__3704 (
            .O(N__21215),
            .I(N__21212));
    InMux I__3703 (
            .O(N__21212),
            .I(N__21206));
    InMux I__3702 (
            .O(N__21211),
            .I(N__21206));
    LocalMux I__3701 (
            .O(N__21206),
            .I(N__21201));
    InMux I__3700 (
            .O(N__21205),
            .I(N__21196));
    CascadeMux I__3699 (
            .O(N__21204),
            .I(N__21193));
    Span4Mux_h I__3698 (
            .O(N__21201),
            .I(N__21190));
    CascadeMux I__3697 (
            .O(N__21200),
            .I(N__21186));
    CascadeMux I__3696 (
            .O(N__21199),
            .I(N__21183));
    LocalMux I__3695 (
            .O(N__21196),
            .I(N__21179));
    InMux I__3694 (
            .O(N__21193),
            .I(N__21176));
    Span4Mux_v I__3693 (
            .O(N__21190),
            .I(N__21173));
    InMux I__3692 (
            .O(N__21189),
            .I(N__21168));
    InMux I__3691 (
            .O(N__21186),
            .I(N__21168));
    InMux I__3690 (
            .O(N__21183),
            .I(N__21163));
    InMux I__3689 (
            .O(N__21182),
            .I(N__21163));
    Span4Mux_s3_v I__3688 (
            .O(N__21179),
            .I(N__21158));
    LocalMux I__3687 (
            .O(N__21176),
            .I(N__21158));
    Odrv4 I__3686 (
            .O(N__21173),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3685 (
            .O(N__21168),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3684 (
            .O(N__21163),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__3683 (
            .O(N__21158),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    CascadeMux I__3682 (
            .O(N__21149),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_12_cascade_ ));
    CascadeMux I__3681 (
            .O(N__21146),
            .I(N__21143));
    InMux I__3680 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__3679 (
            .O(N__21140),
            .I(N__21137));
    Span4Mux_h I__3678 (
            .O(N__21137),
            .I(N__21134));
    Odrv4 I__3677 (
            .O(N__21134),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_14 ));
    InMux I__3676 (
            .O(N__21131),
            .I(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ));
    InMux I__3675 (
            .O(N__21128),
            .I(bfn_7_13_0_));
    InMux I__3674 (
            .O(N__21125),
            .I(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ));
    InMux I__3673 (
            .O(N__21122),
            .I(N__21116));
    InMux I__3672 (
            .O(N__21121),
            .I(N__21116));
    LocalMux I__3671 (
            .O(N__21116),
            .I(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ));
    InMux I__3670 (
            .O(N__21113),
            .I(\POWERLED.un1_dutycycle_94_cry_9 ));
    InMux I__3669 (
            .O(N__21110),
            .I(\POWERLED.un1_dutycycle_94_cry_10 ));
    InMux I__3668 (
            .O(N__21107),
            .I(\POWERLED.un1_dutycycle_94_cry_11 ));
    InMux I__3667 (
            .O(N__21104),
            .I(N__21098));
    InMux I__3666 (
            .O(N__21103),
            .I(N__21098));
    LocalMux I__3665 (
            .O(N__21098),
            .I(N__21095));
    Odrv12 I__3664 (
            .O(N__21095),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ));
    InMux I__3663 (
            .O(N__21092),
            .I(\POWERLED.un1_dutycycle_94_cry_12 ));
    CascadeMux I__3662 (
            .O(N__21089),
            .I(N__21085));
    InMux I__3661 (
            .O(N__21088),
            .I(N__21080));
    InMux I__3660 (
            .O(N__21085),
            .I(N__21080));
    LocalMux I__3659 (
            .O(N__21080),
            .I(N__21077));
    Odrv4 I__3658 (
            .O(N__21077),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ));
    InMux I__3657 (
            .O(N__21074),
            .I(\POWERLED.un1_dutycycle_94_cry_13 ));
    InMux I__3656 (
            .O(N__21071),
            .I(\POWERLED.un1_dutycycle_94_cry_14 ));
    InMux I__3655 (
            .O(N__21068),
            .I(N__21065));
    LocalMux I__3654 (
            .O(N__21065),
            .I(N__21062));
    Span4Mux_h I__3653 (
            .O(N__21062),
            .I(N__21058));
    InMux I__3652 (
            .O(N__21061),
            .I(N__21055));
    Odrv4 I__3651 (
            .O(N__21058),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ));
    LocalMux I__3650 (
            .O(N__21055),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ));
    CascadeMux I__3649 (
            .O(N__21050),
            .I(\POWERLED.un1_dutycycle_53_13_4_cascade_ ));
    InMux I__3648 (
            .O(N__21047),
            .I(N__21044));
    LocalMux I__3647 (
            .O(N__21044),
            .I(N__21041));
    Span4Mux_v I__3646 (
            .O(N__21041),
            .I(N__21038));
    Odrv4 I__3645 (
            .O(N__21038),
            .I(\POWERLED.un1_dutycycle_53_13_3 ));
    CascadeMux I__3644 (
            .O(N__21035),
            .I(N__21032));
    InMux I__3643 (
            .O(N__21032),
            .I(N__21029));
    LocalMux I__3642 (
            .O(N__21029),
            .I(N__21026));
    Span4Mux_h I__3641 (
            .O(N__21026),
            .I(N__21023));
    Odrv4 I__3640 (
            .O(N__21023),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_11 ));
    InMux I__3639 (
            .O(N__21020),
            .I(N__21014));
    InMux I__3638 (
            .O(N__21019),
            .I(N__21014));
    LocalMux I__3637 (
            .O(N__21014),
            .I(\POWERLED.g0_0_1 ));
    InMux I__3636 (
            .O(N__21011),
            .I(N__21008));
    LocalMux I__3635 (
            .O(N__21008),
            .I(N__21005));
    Odrv12 I__3634 (
            .O(N__21005),
            .I(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ));
    InMux I__3633 (
            .O(N__21002),
            .I(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ));
    InMux I__3632 (
            .O(N__20999),
            .I(N__20996));
    LocalMux I__3631 (
            .O(N__20996),
            .I(N__20993));
    Odrv12 I__3630 (
            .O(N__20993),
            .I(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ));
    InMux I__3629 (
            .O(N__20990),
            .I(\POWERLED.un1_dutycycle_94_cry_1 ));
    InMux I__3628 (
            .O(N__20987),
            .I(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ));
    InMux I__3627 (
            .O(N__20984),
            .I(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ));
    InMux I__3626 (
            .O(N__20981),
            .I(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ));
    InMux I__3625 (
            .O(N__20978),
            .I(N__20975));
    LocalMux I__3624 (
            .O(N__20975),
            .I(N__20972));
    Odrv4 I__3623 (
            .O(N__20972),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ));
    InMux I__3622 (
            .O(N__20969),
            .I(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ));
    CascadeMux I__3621 (
            .O(N__20966),
            .I(\POWERLED.d_i3_mux_cascade_ ));
    InMux I__3620 (
            .O(N__20963),
            .I(N__20960));
    LocalMux I__3619 (
            .O(N__20960),
            .I(N__20957));
    Span4Mux_h I__3618 (
            .O(N__20957),
            .I(N__20954));
    Odrv4 I__3617 (
            .O(N__20954),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_5 ));
    CascadeMux I__3616 (
            .O(N__20951),
            .I(N__20948));
    InMux I__3615 (
            .O(N__20948),
            .I(N__20945));
    LocalMux I__3614 (
            .O(N__20945),
            .I(N__20942));
    Odrv12 I__3613 (
            .O(N__20942),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_0 ));
    CascadeMux I__3612 (
            .O(N__20939),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3_cascade_ ));
    CascadeMux I__3611 (
            .O(N__20936),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_9_cascade_ ));
    CascadeMux I__3610 (
            .O(N__20933),
            .I(N__20930));
    InMux I__3609 (
            .O(N__20930),
            .I(N__20927));
    LocalMux I__3608 (
            .O(N__20927),
            .I(N__20924));
    Odrv4 I__3607 (
            .O(N__20924),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_7 ));
    InMux I__3606 (
            .O(N__20921),
            .I(N__20918));
    LocalMux I__3605 (
            .O(N__20918),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    InMux I__3604 (
            .O(N__20915),
            .I(N__20912));
    LocalMux I__3603 (
            .O(N__20912),
            .I(N__20909));
    Odrv4 I__3602 (
            .O(N__20909),
            .I(\POWERLED.dutycycle_RNIZ0Z_5 ));
    CascadeMux I__3601 (
            .O(N__20906),
            .I(N__20903));
    InMux I__3600 (
            .O(N__20903),
            .I(N__20900));
    LocalMux I__3599 (
            .O(N__20900),
            .I(N__20897));
    Span4Mux_v I__3598 (
            .O(N__20897),
            .I(N__20894));
    Odrv4 I__3597 (
            .O(N__20894),
            .I(\POWERLED.un1_dutycycle_53_13_4_1 ));
    CascadeMux I__3596 (
            .O(N__20891),
            .I(\POWERLED.func_state_RNIBVNS_1Z0Z_0_cascade_ ));
    InMux I__3595 (
            .O(N__20888),
            .I(N__20885));
    LocalMux I__3594 (
            .O(N__20885),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_ns_1 ));
    CascadeMux I__3593 (
            .O(N__20882),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ));
    InMux I__3592 (
            .O(N__20879),
            .I(N__20873));
    InMux I__3591 (
            .O(N__20878),
            .I(N__20873));
    LocalMux I__3590 (
            .O(N__20873),
            .I(\POWERLED.N_171 ));
    InMux I__3589 (
            .O(N__20870),
            .I(N__20867));
    LocalMux I__3588 (
            .O(N__20867),
            .I(\POWERLED.N_283 ));
    CascadeMux I__3587 (
            .O(N__20864),
            .I(N__20861));
    InMux I__3586 (
            .O(N__20861),
            .I(N__20858));
    LocalMux I__3585 (
            .O(N__20858),
            .I(N__20855));
    Span4Mux_v I__3584 (
            .O(N__20855),
            .I(N__20852));
    Odrv4 I__3583 (
            .O(N__20852),
            .I(\POWERLED.N_275_0 ));
    CascadeMux I__3582 (
            .O(N__20849),
            .I(N__20846));
    InMux I__3581 (
            .O(N__20846),
            .I(N__20843));
    LocalMux I__3580 (
            .O(N__20843),
            .I(\POWERLED.dutycycle_set_0_0 ));
    InMux I__3579 (
            .O(N__20840),
            .I(N__20834));
    InMux I__3578 (
            .O(N__20839),
            .I(N__20834));
    LocalMux I__3577 (
            .O(N__20834),
            .I(\POWERLED.dutycycle_eena_13_0 ));
    CascadeMux I__3576 (
            .O(N__20831),
            .I(\POWERLED.dutycycle_set_0_0_cascade_ ));
    InMux I__3575 (
            .O(N__20828),
            .I(N__20822));
    InMux I__3574 (
            .O(N__20827),
            .I(N__20822));
    LocalMux I__3573 (
            .O(N__20822),
            .I(\POWERLED.dutycycle_0_6 ));
    CascadeMux I__3572 (
            .O(N__20819),
            .I(\POWERLED.dutycycleZ0Z_6_cascade_ ));
    CascadeMux I__3571 (
            .O(N__20816),
            .I(N__20813));
    InMux I__3570 (
            .O(N__20813),
            .I(N__20810));
    LocalMux I__3569 (
            .O(N__20810),
            .I(N__20807));
    Sp12to4 I__3568 (
            .O(N__20807),
            .I(N__20804));
    Span12Mux_s9_v I__3567 (
            .O(N__20804),
            .I(N__20800));
    InMux I__3566 (
            .O(N__20803),
            .I(N__20797));
    Odrv12 I__3565 (
            .O(N__20800),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_0 ));
    LocalMux I__3564 (
            .O(N__20797),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_0 ));
    CascadeMux I__3563 (
            .O(N__20792),
            .I(\POWERLED.dutycycle_en_10_cascade_ ));
    InMux I__3562 (
            .O(N__20789),
            .I(N__20783));
    InMux I__3561 (
            .O(N__20788),
            .I(N__20783));
    LocalMux I__3560 (
            .O(N__20783),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    InMux I__3559 (
            .O(N__20780),
            .I(N__20777));
    LocalMux I__3558 (
            .O(N__20777),
            .I(N__20774));
    Odrv4 I__3557 (
            .O(N__20774),
            .I(\POWERLED.un1_func_state25_4_i_a2_1 ));
    CascadeMux I__3556 (
            .O(N__20771),
            .I(\POWERLED.N_301_cascade_ ));
    InMux I__3555 (
            .O(N__20768),
            .I(N__20765));
    LocalMux I__3554 (
            .O(N__20765),
            .I(N__20762));
    Span4Mux_v I__3553 (
            .O(N__20762),
            .I(N__20758));
    InMux I__3552 (
            .O(N__20761),
            .I(N__20755));
    Odrv4 I__3551 (
            .O(N__20758),
            .I(\POWERLED.N_341 ));
    LocalMux I__3550 (
            .O(N__20755),
            .I(\POWERLED.N_341 ));
    CascadeMux I__3549 (
            .O(N__20750),
            .I(\POWERLED.count_clk_en_1_0_cascade_ ));
    CascadeMux I__3548 (
            .O(N__20747),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_0_cascade_ ));
    CascadeMux I__3547 (
            .O(N__20744),
            .I(\POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_cascade_ ));
    InMux I__3546 (
            .O(N__20741),
            .I(N__20738));
    LocalMux I__3545 (
            .O(N__20738),
            .I(N__20735));
    Span4Mux_v I__3544 (
            .O(N__20735),
            .I(N__20732));
    Span4Mux_h I__3543 (
            .O(N__20732),
            .I(N__20727));
    InMux I__3542 (
            .O(N__20731),
            .I(N__20724));
    InMux I__3541 (
            .O(N__20730),
            .I(N__20721));
    Odrv4 I__3540 (
            .O(N__20727),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__3539 (
            .O(N__20724),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__3538 (
            .O(N__20721),
            .I(\POWERLED.countZ0Z_5 ));
    CascadeMux I__3537 (
            .O(N__20714),
            .I(N__20711));
    InMux I__3536 (
            .O(N__20711),
            .I(N__20705));
    InMux I__3535 (
            .O(N__20710),
            .I(N__20705));
    LocalMux I__3534 (
            .O(N__20705),
            .I(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ));
    InMux I__3533 (
            .O(N__20702),
            .I(N__20699));
    LocalMux I__3532 (
            .O(N__20699),
            .I(\POWERLED.count_0_5 ));
    InMux I__3531 (
            .O(N__20696),
            .I(N__20693));
    LocalMux I__3530 (
            .O(N__20693),
            .I(N__20690));
    Span4Mux_v I__3529 (
            .O(N__20690),
            .I(N__20687));
    Span4Mux_h I__3528 (
            .O(N__20687),
            .I(N__20682));
    InMux I__3527 (
            .O(N__20686),
            .I(N__20679));
    InMux I__3526 (
            .O(N__20685),
            .I(N__20676));
    Odrv4 I__3525 (
            .O(N__20682),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__3524 (
            .O(N__20679),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__3523 (
            .O(N__20676),
            .I(\POWERLED.countZ0Z_14 ));
    CascadeMux I__3522 (
            .O(N__20669),
            .I(N__20666));
    InMux I__3521 (
            .O(N__20666),
            .I(N__20660));
    InMux I__3520 (
            .O(N__20665),
            .I(N__20660));
    LocalMux I__3519 (
            .O(N__20660),
            .I(\POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ));
    InMux I__3518 (
            .O(N__20657),
            .I(N__20654));
    LocalMux I__3517 (
            .O(N__20654),
            .I(\POWERLED.count_0_14 ));
    InMux I__3516 (
            .O(N__20651),
            .I(N__20648));
    LocalMux I__3515 (
            .O(N__20648),
            .I(N__20645));
    Span4Mux_v I__3514 (
            .O(N__20645),
            .I(N__20642));
    Span4Mux_h I__3513 (
            .O(N__20642),
            .I(N__20637));
    InMux I__3512 (
            .O(N__20641),
            .I(N__20634));
    InMux I__3511 (
            .O(N__20640),
            .I(N__20631));
    Odrv4 I__3510 (
            .O(N__20637),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__3509 (
            .O(N__20634),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__3508 (
            .O(N__20631),
            .I(\POWERLED.countZ0Z_6 ));
    CascadeMux I__3507 (
            .O(N__20624),
            .I(N__20621));
    InMux I__3506 (
            .O(N__20621),
            .I(N__20615));
    InMux I__3505 (
            .O(N__20620),
            .I(N__20615));
    LocalMux I__3504 (
            .O(N__20615),
            .I(\POWERLED.un1_count_cry_5_c_RNIFAZ0Z49 ));
    InMux I__3503 (
            .O(N__20612),
            .I(N__20609));
    LocalMux I__3502 (
            .O(N__20609),
            .I(\POWERLED.count_0_6 ));
    CascadeMux I__3501 (
            .O(N__20606),
            .I(\POWERLED.dutycycleZ0Z_11_cascade_ ));
    CascadeMux I__3500 (
            .O(N__20603),
            .I(\POWERLED.N_148_N_cascade_ ));
    CascadeMux I__3499 (
            .O(N__20600),
            .I(N__20597));
    InMux I__3498 (
            .O(N__20597),
            .I(N__20594));
    LocalMux I__3497 (
            .O(N__20594),
            .I(\POWERLED.dutycycle_en_10 ));
    InMux I__3496 (
            .O(N__20591),
            .I(N__20588));
    LocalMux I__3495 (
            .O(N__20588),
            .I(\POWERLED.dutycycle_1_0_0 ));
    InMux I__3494 (
            .O(N__20585),
            .I(N__20581));
    InMux I__3493 (
            .O(N__20584),
            .I(N__20578));
    LocalMux I__3492 (
            .O(N__20581),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    LocalMux I__3491 (
            .O(N__20578),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    CascadeMux I__3490 (
            .O(N__20573),
            .I(\POWERLED.dutycycle_1_0_0_cascade_ ));
    InMux I__3489 (
            .O(N__20570),
            .I(N__20564));
    InMux I__3488 (
            .O(N__20569),
            .I(N__20564));
    LocalMux I__3487 (
            .O(N__20564),
            .I(N__20561));
    Span4Mux_h I__3486 (
            .O(N__20561),
            .I(N__20558));
    Odrv4 I__3485 (
            .O(N__20558),
            .I(\POWERLED.dutycycle_eena ));
    CascadeMux I__3484 (
            .O(N__20555),
            .I(N__20552));
    InMux I__3483 (
            .O(N__20552),
            .I(N__20549));
    LocalMux I__3482 (
            .O(N__20549),
            .I(N__20546));
    Span4Mux_h I__3481 (
            .O(N__20546),
            .I(N__20542));
    InMux I__3480 (
            .O(N__20545),
            .I(N__20539));
    Span4Mux_h I__3479 (
            .O(N__20542),
            .I(N__20536));
    LocalMux I__3478 (
            .O(N__20539),
            .I(\POWERLED.func_stateZ0Z_1 ));
    Odrv4 I__3477 (
            .O(N__20536),
            .I(\POWERLED.func_stateZ0Z_1 ));
    InMux I__3476 (
            .O(N__20531),
            .I(N__20528));
    LocalMux I__3475 (
            .O(N__20528),
            .I(N__20525));
    Span12Mux_s6_h I__3474 (
            .O(N__20525),
            .I(N__20521));
    InMux I__3473 (
            .O(N__20524),
            .I(N__20518));
    Odrv12 I__3472 (
            .O(N__20521),
            .I(\POWERLED.func_state_RNIG5G37Z0Z_1 ));
    LocalMux I__3471 (
            .O(N__20518),
            .I(\POWERLED.func_state_RNIG5G37Z0Z_1 ));
    CascadeMux I__3470 (
            .O(N__20513),
            .I(\POWERLED.func_state_cascade_ ));
    CascadeMux I__3469 (
            .O(N__20510),
            .I(N__20507));
    InMux I__3468 (
            .O(N__20507),
            .I(N__20504));
    LocalMux I__3467 (
            .O(N__20504),
            .I(N__20500));
    InMux I__3466 (
            .O(N__20503),
            .I(N__20497));
    Span4Mux_v I__3465 (
            .O(N__20500),
            .I(N__20494));
    LocalMux I__3464 (
            .O(N__20497),
            .I(N__20491));
    Odrv4 I__3463 (
            .O(N__20494),
            .I(\POWERLED.dutycycle_1_0_1 ));
    Odrv4 I__3462 (
            .O(N__20491),
            .I(\POWERLED.dutycycle_1_0_1 ));
    InMux I__3461 (
            .O(N__20486),
            .I(N__20483));
    LocalMux I__3460 (
            .O(N__20483),
            .I(N__20480));
    Span4Mux_v I__3459 (
            .O(N__20480),
            .I(N__20477));
    Span4Mux_h I__3458 (
            .O(N__20477),
            .I(N__20472));
    InMux I__3457 (
            .O(N__20476),
            .I(N__20469));
    InMux I__3456 (
            .O(N__20475),
            .I(N__20466));
    Odrv4 I__3455 (
            .O(N__20472),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__3454 (
            .O(N__20469),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__3453 (
            .O(N__20466),
            .I(\POWERLED.countZ0Z_13 ));
    CascadeMux I__3452 (
            .O(N__20459),
            .I(N__20456));
    InMux I__3451 (
            .O(N__20456),
            .I(N__20450));
    InMux I__3450 (
            .O(N__20455),
            .I(N__20450));
    LocalMux I__3449 (
            .O(N__20450),
            .I(\POWERLED.un1_count_cry_12_c_RNITGIZ0Z7 ));
    InMux I__3448 (
            .O(N__20447),
            .I(N__20444));
    LocalMux I__3447 (
            .O(N__20444),
            .I(\POWERLED.count_0_13 ));
    InMux I__3446 (
            .O(N__20441),
            .I(N__20438));
    LocalMux I__3445 (
            .O(N__20438),
            .I(N__20435));
    Sp12to4 I__3444 (
            .O(N__20435),
            .I(N__20432));
    Odrv12 I__3443 (
            .O(N__20432),
            .I(\POWERLED.func_state_RNIMQ0FZ0Z_1 ));
    InMux I__3442 (
            .O(N__20429),
            .I(N__20426));
    LocalMux I__3441 (
            .O(N__20426),
            .I(\POWERLED.N_309 ));
    CascadeMux I__3440 (
            .O(N__20423),
            .I(\POWERLED.func_state_1_m0_1_cascade_ ));
    CascadeMux I__3439 (
            .O(N__20420),
            .I(\POWERLED.count_RNI_0_1_cascade_ ));
    CascadeMux I__3438 (
            .O(N__20417),
            .I(\POWERLED.dutycycle_1_0_iv_i_a3_1_0_2_cascade_ ));
    InMux I__3437 (
            .O(N__20414),
            .I(N__20408));
    InMux I__3436 (
            .O(N__20413),
            .I(N__20408));
    LocalMux I__3435 (
            .O(N__20408),
            .I(N__20405));
    Span4Mux_v I__3434 (
            .O(N__20405),
            .I(N__20402));
    Odrv4 I__3433 (
            .O(N__20402),
            .I(\POWERLED.N_64 ));
    CascadeMux I__3432 (
            .O(N__20399),
            .I(\POWERLED.g0_0_a3_1_cascade_ ));
    InMux I__3431 (
            .O(N__20396),
            .I(N__20393));
    LocalMux I__3430 (
            .O(N__20393),
            .I(N__20390));
    Span4Mux_v I__3429 (
            .O(N__20390),
            .I(N__20387));
    Odrv4 I__3428 (
            .O(N__20387),
            .I(\POWERLED.g0_3_1 ));
    InMux I__3427 (
            .O(N__20384),
            .I(N__20381));
    LocalMux I__3426 (
            .O(N__20381),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_2 ));
    CascadeMux I__3425 (
            .O(N__20378),
            .I(\HDA_STRAP.N_14_cascade_ ));
    InMux I__3424 (
            .O(N__20375),
            .I(N__20369));
    InMux I__3423 (
            .O(N__20374),
            .I(N__20369));
    LocalMux I__3422 (
            .O(N__20369),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    IoInMux I__3421 (
            .O(N__20366),
            .I(N__20363));
    LocalMux I__3420 (
            .O(N__20363),
            .I(N__20360));
    IoSpan4Mux I__3419 (
            .O(N__20360),
            .I(N__20357));
    Span4Mux_s2_h I__3418 (
            .O(N__20357),
            .I(N__20354));
    Span4Mux_h I__3417 (
            .O(N__20354),
            .I(N__20351));
    Odrv4 I__3416 (
            .O(N__20351),
            .I(hda_sdo_atp));
    InMux I__3415 (
            .O(N__20348),
            .I(N__20345));
    LocalMux I__3414 (
            .O(N__20345),
            .I(N__20342));
    Span4Mux_h I__3413 (
            .O(N__20342),
            .I(N__20339));
    Odrv4 I__3412 (
            .O(N__20339),
            .I(gpio_fpga_soc_1));
    CascadeMux I__3411 (
            .O(N__20336),
            .I(\HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_ ));
    InMux I__3410 (
            .O(N__20333),
            .I(N__20327));
    InMux I__3409 (
            .O(N__20332),
            .I(N__20327));
    LocalMux I__3408 (
            .O(N__20327),
            .I(N__20323));
    InMux I__3407 (
            .O(N__20326),
            .I(N__20320));
    Odrv12 I__3406 (
            .O(N__20323),
            .I(PCH_PWRGD_delayed_vccin_ok));
    LocalMux I__3405 (
            .O(N__20320),
            .I(PCH_PWRGD_delayed_vccin_ok));
    InMux I__3404 (
            .O(N__20315),
            .I(N__20312));
    LocalMux I__3403 (
            .O(N__20312),
            .I(\HDA_STRAP.curr_state_RNO_0Z0Z_0 ));
    InMux I__3402 (
            .O(N__20309),
            .I(N__20306));
    LocalMux I__3401 (
            .O(N__20306),
            .I(\HDA_STRAP.N_5_0 ));
    CascadeMux I__3400 (
            .O(N__20303),
            .I(\POWERLED.N_341_cascade_ ));
    CascadeMux I__3399 (
            .O(N__20300),
            .I(\POWERLED.dutycycle_RNI_11Z0Z_7_cascade_ ));
    CascadeMux I__3398 (
            .O(N__20297),
            .I(N__20294));
    InMux I__3397 (
            .O(N__20294),
            .I(N__20291));
    LocalMux I__3396 (
            .O(N__20291),
            .I(N__20288));
    Odrv4 I__3395 (
            .O(N__20288),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_12 ));
    InMux I__3394 (
            .O(N__20285),
            .I(N__20282));
    LocalMux I__3393 (
            .O(N__20282),
            .I(\POWERLED.un1_dutycycle_53_4_1 ));
    CascadeMux I__3392 (
            .O(N__20279),
            .I(\POWERLED.dutycycleZ0Z_3_cascade_ ));
    CascadeMux I__3391 (
            .O(N__20276),
            .I(N__20273));
    InMux I__3390 (
            .O(N__20273),
            .I(N__20270));
    LocalMux I__3389 (
            .O(N__20270),
            .I(\POWERLED.un1_dutycycle_53_45_a0_1 ));
    CascadeMux I__3388 (
            .O(N__20267),
            .I(\POWERLED.un1_dutycycle_53_45_a0_1_cascade_ ));
    InMux I__3387 (
            .O(N__20264),
            .I(N__20261));
    LocalMux I__3386 (
            .O(N__20261),
            .I(N__20258));
    Span4Mux_v I__3385 (
            .O(N__20258),
            .I(N__20255));
    Odrv4 I__3384 (
            .O(N__20255),
            .I(\POWERLED.un1_dutycycle_53_10_1 ));
    CascadeMux I__3383 (
            .O(N__20252),
            .I(N__20249));
    InMux I__3382 (
            .O(N__20249),
            .I(N__20246));
    LocalMux I__3381 (
            .O(N__20246),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__3380 (
            .O(N__20243),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    CascadeMux I__3379 (
            .O(N__20240),
            .I(N__20237));
    InMux I__3378 (
            .O(N__20237),
            .I(N__20234));
    LocalMux I__3377 (
            .O(N__20234),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    CascadeMux I__3376 (
            .O(N__20231),
            .I(N__20228));
    InMux I__3375 (
            .O(N__20228),
            .I(N__20225));
    LocalMux I__3374 (
            .O(N__20225),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__3373 (
            .O(N__20222),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    InMux I__3372 (
            .O(N__20219),
            .I(N__20216));
    LocalMux I__3371 (
            .O(N__20216),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__3370 (
            .O(N__20213),
            .I(N__20210));
    LocalMux I__3369 (
            .O(N__20210),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__3368 (
            .O(N__20207),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    InMux I__3367 (
            .O(N__20204),
            .I(N__20200));
    CascadeMux I__3366 (
            .O(N__20203),
            .I(N__20196));
    LocalMux I__3365 (
            .O(N__20200),
            .I(N__20192));
    InMux I__3364 (
            .O(N__20199),
            .I(N__20187));
    InMux I__3363 (
            .O(N__20196),
            .I(N__20187));
    InMux I__3362 (
            .O(N__20195),
            .I(N__20184));
    Odrv4 I__3361 (
            .O(N__20192),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3360 (
            .O(N__20187),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3359 (
            .O(N__20184),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    CascadeMux I__3358 (
            .O(N__20177),
            .I(N__20174));
    InMux I__3357 (
            .O(N__20174),
            .I(N__20171));
    LocalMux I__3356 (
            .O(N__20171),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__3355 (
            .O(N__20168),
            .I(N__20165));
    LocalMux I__3354 (
            .O(N__20165),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__3353 (
            .O(N__20162),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    InMux I__3352 (
            .O(N__20159),
            .I(N__20156));
    LocalMux I__3351 (
            .O(N__20156),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    CascadeMux I__3350 (
            .O(N__20153),
            .I(N__20149));
    CascadeMux I__3349 (
            .O(N__20152),
            .I(N__20145));
    InMux I__3348 (
            .O(N__20149),
            .I(N__20138));
    InMux I__3347 (
            .O(N__20148),
            .I(N__20138));
    InMux I__3346 (
            .O(N__20145),
            .I(N__20138));
    LocalMux I__3345 (
            .O(N__20138),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    CascadeMux I__3344 (
            .O(N__20135),
            .I(N__20132));
    InMux I__3343 (
            .O(N__20132),
            .I(N__20129));
    LocalMux I__3342 (
            .O(N__20129),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__3341 (
            .O(N__20126),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    CascadeMux I__3340 (
            .O(N__20123),
            .I(N__20120));
    InMux I__3339 (
            .O(N__20120),
            .I(N__20117));
    LocalMux I__3338 (
            .O(N__20117),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__3337 (
            .O(N__20114),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    InMux I__3336 (
            .O(N__20111),
            .I(N__20108));
    LocalMux I__3335 (
            .O(N__20108),
            .I(N__20104));
    CascadeMux I__3334 (
            .O(N__20107),
            .I(N__20100));
    Span4Mux_h I__3333 (
            .O(N__20104),
            .I(N__20095));
    InMux I__3332 (
            .O(N__20103),
            .I(N__20092));
    InMux I__3331 (
            .O(N__20100),
            .I(N__20085));
    InMux I__3330 (
            .O(N__20099),
            .I(N__20085));
    InMux I__3329 (
            .O(N__20098),
            .I(N__20085));
    Odrv4 I__3328 (
            .O(N__20095),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__3327 (
            .O(N__20092),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__3326 (
            .O(N__20085),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    InMux I__3325 (
            .O(N__20078),
            .I(N__20075));
    LocalMux I__3324 (
            .O(N__20075),
            .I(N__20071));
    InMux I__3323 (
            .O(N__20074),
            .I(N__20068));
    Span4Mux_v I__3322 (
            .O(N__20071),
            .I(N__20065));
    LocalMux I__3321 (
            .O(N__20068),
            .I(N__20062));
    Odrv4 I__3320 (
            .O(N__20065),
            .I(\POWERLED.mult1_un68_sum ));
    Odrv12 I__3319 (
            .O(N__20062),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__3318 (
            .O(N__20057),
            .I(N__20054));
    LocalMux I__3317 (
            .O(N__20054),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__3316 (
            .O(N__20051),
            .I(N__20048));
    LocalMux I__3315 (
            .O(N__20048),
            .I(N__20043));
    InMux I__3314 (
            .O(N__20047),
            .I(N__20040));
    InMux I__3313 (
            .O(N__20046),
            .I(N__20037));
    Odrv4 I__3312 (
            .O(N__20043),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__3311 (
            .O(N__20040),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__3310 (
            .O(N__20037),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    InMux I__3309 (
            .O(N__20030),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__3308 (
            .O(N__20027),
            .I(N__20024));
    InMux I__3307 (
            .O(N__20024),
            .I(N__20021));
    LocalMux I__3306 (
            .O(N__20021),
            .I(N__20018));
    Odrv4 I__3305 (
            .O(N__20018),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__3304 (
            .O(N__20015),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__3303 (
            .O(N__20012),
            .I(N__20009));
    InMux I__3302 (
            .O(N__20009),
            .I(N__20006));
    LocalMux I__3301 (
            .O(N__20006),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__3300 (
            .O(N__20003),
            .I(N__20000));
    InMux I__3299 (
            .O(N__20000),
            .I(N__19997));
    LocalMux I__3298 (
            .O(N__19997),
            .I(N__19994));
    Odrv4 I__3297 (
            .O(N__19994),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__3296 (
            .O(N__19991),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__3295 (
            .O(N__19988),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    CascadeMux I__3294 (
            .O(N__19985),
            .I(N__19982));
    InMux I__3293 (
            .O(N__19982),
            .I(N__19979));
    LocalMux I__3292 (
            .O(N__19979),
            .I(\POWERLED.un1_dutycycle_53_i_29 ));
    CascadeMux I__3291 (
            .O(N__19976),
            .I(N__19971));
    CascadeMux I__3290 (
            .O(N__19975),
            .I(N__19967));
    InMux I__3289 (
            .O(N__19974),
            .I(N__19962));
    InMux I__3288 (
            .O(N__19971),
            .I(N__19962));
    InMux I__3287 (
            .O(N__19970),
            .I(N__19957));
    InMux I__3286 (
            .O(N__19967),
            .I(N__19957));
    LocalMux I__3285 (
            .O(N__19962),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    LocalMux I__3284 (
            .O(N__19957),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    InMux I__3283 (
            .O(N__19952),
            .I(N__19945));
    InMux I__3282 (
            .O(N__19951),
            .I(N__19945));
    InMux I__3281 (
            .O(N__19950),
            .I(N__19942));
    LocalMux I__3280 (
            .O(N__19945),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    LocalMux I__3279 (
            .O(N__19942),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    CascadeMux I__3278 (
            .O(N__19937),
            .I(N__19934));
    InMux I__3277 (
            .O(N__19934),
            .I(N__19931));
    LocalMux I__3276 (
            .O(N__19931),
            .I(\POWERLED.mult1_un47_sum_s_4_sf ));
    CascadeMux I__3275 (
            .O(N__19928),
            .I(N__19924));
    InMux I__3274 (
            .O(N__19927),
            .I(N__19921));
    InMux I__3273 (
            .O(N__19924),
            .I(N__19918));
    LocalMux I__3272 (
            .O(N__19921),
            .I(N__19915));
    LocalMux I__3271 (
            .O(N__19918),
            .I(N__19912));
    Span4Mux_h I__3270 (
            .O(N__19915),
            .I(N__19909));
    Odrv4 I__3269 (
            .O(N__19912),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    Odrv4 I__3268 (
            .O(N__19909),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    CascadeMux I__3267 (
            .O(N__19904),
            .I(N__19900));
    InMux I__3266 (
            .O(N__19903),
            .I(N__19897));
    InMux I__3265 (
            .O(N__19900),
            .I(N__19894));
    LocalMux I__3264 (
            .O(N__19897),
            .I(N__19891));
    LocalMux I__3263 (
            .O(N__19894),
            .I(N__19888));
    Span4Mux_h I__3262 (
            .O(N__19891),
            .I(N__19885));
    Odrv4 I__3261 (
            .O(N__19888),
            .I(\POWERLED.dutycycle_en_12 ));
    Odrv4 I__3260 (
            .O(N__19885),
            .I(\POWERLED.dutycycle_en_12 ));
    InMux I__3259 (
            .O(N__19880),
            .I(N__19876));
    InMux I__3258 (
            .O(N__19879),
            .I(N__19873));
    LocalMux I__3257 (
            .O(N__19876),
            .I(N__19870));
    LocalMux I__3256 (
            .O(N__19873),
            .I(\POWERLED.mult1_un75_sum ));
    Odrv4 I__3255 (
            .O(N__19870),
            .I(\POWERLED.mult1_un75_sum ));
    CascadeMux I__3254 (
            .O(N__19865),
            .I(\POWERLED.un1_dutycycle_53_axb_10_1_cascade_ ));
    CascadeMux I__3253 (
            .O(N__19862),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_9_cascade_ ));
    CascadeMux I__3252 (
            .O(N__19859),
            .I(N__19856));
    InMux I__3251 (
            .O(N__19856),
            .I(N__19853));
    LocalMux I__3250 (
            .O(N__19853),
            .I(\POWERLED.dutycycle_RNIZ0Z_13 ));
    InMux I__3249 (
            .O(N__19850),
            .I(N__19844));
    InMux I__3248 (
            .O(N__19849),
            .I(N__19844));
    LocalMux I__3247 (
            .O(N__19844),
            .I(\POWERLED.dutycycleZ1Z_10 ));
    CascadeMux I__3246 (
            .O(N__19841),
            .I(\POWERLED.dutycycleZ0Z_2_cascade_ ));
    InMux I__3245 (
            .O(N__19838),
            .I(N__19835));
    LocalMux I__3244 (
            .O(N__19835),
            .I(\POWERLED.dutycycle_RNIZ0Z_10 ));
    CascadeMux I__3243 (
            .O(N__19832),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_9_cascade_ ));
    CascadeMux I__3242 (
            .O(N__19829),
            .I(N__19825));
    InMux I__3241 (
            .O(N__19828),
            .I(N__19822));
    InMux I__3240 (
            .O(N__19825),
            .I(N__19819));
    LocalMux I__3239 (
            .O(N__19822),
            .I(\POWERLED.mult1_un47_sum ));
    LocalMux I__3238 (
            .O(N__19819),
            .I(\POWERLED.mult1_un47_sum ));
    InMux I__3237 (
            .O(N__19814),
            .I(N__19811));
    LocalMux I__3236 (
            .O(N__19811),
            .I(\POWERLED.N_353_0 ));
    CascadeMux I__3235 (
            .O(N__19808),
            .I(\POWERLED.dutycycleZ0Z_10_cascade_ ));
    CascadeMux I__3234 (
            .O(N__19805),
            .I(N__19802));
    InMux I__3233 (
            .O(N__19802),
            .I(N__19799));
    LocalMux I__3232 (
            .O(N__19799),
            .I(N__19796));
    Odrv4 I__3231 (
            .O(N__19796),
            .I(\POWERLED.dutycycle_RNIZ0Z_14 ));
    CascadeMux I__3230 (
            .O(N__19793),
            .I(\POWERLED.N_86_f0_cascade_ ));
    InMux I__3229 (
            .O(N__19790),
            .I(N__19787));
    LocalMux I__3228 (
            .O(N__19787),
            .I(\POWERLED.dutycycle_en_11 ));
    CascadeMux I__3227 (
            .O(N__19784),
            .I(\POWERLED.dutycycle_en_11_cascade_ ));
    InMux I__3226 (
            .O(N__19781),
            .I(N__19778));
    LocalMux I__3225 (
            .O(N__19778),
            .I(N__19774));
    InMux I__3224 (
            .O(N__19777),
            .I(N__19771));
    Span4Mux_h I__3223 (
            .O(N__19774),
            .I(N__19768));
    LocalMux I__3222 (
            .O(N__19771),
            .I(\POWERLED.dutycycleZ1Z_14 ));
    Odrv4 I__3221 (
            .O(N__19768),
            .I(\POWERLED.dutycycleZ1Z_14 ));
    CascadeMux I__3220 (
            .O(N__19763),
            .I(N__19760));
    InMux I__3219 (
            .O(N__19760),
            .I(N__19757));
    LocalMux I__3218 (
            .O(N__19757),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_15 ));
    CascadeMux I__3217 (
            .O(N__19754),
            .I(N__19750));
    InMux I__3216 (
            .O(N__19753),
            .I(N__19747));
    InMux I__3215 (
            .O(N__19750),
            .I(N__19744));
    LocalMux I__3214 (
            .O(N__19747),
            .I(N__19741));
    LocalMux I__3213 (
            .O(N__19744),
            .I(N__19738));
    Span4Mux_v I__3212 (
            .O(N__19741),
            .I(N__19735));
    Span12Mux_s10_h I__3211 (
            .O(N__19738),
            .I(N__19732));
    Odrv4 I__3210 (
            .O(N__19735),
            .I(\POWERLED.N_2215_i ));
    Odrv12 I__3209 (
            .O(N__19732),
            .I(\POWERLED.N_2215_i ));
    CascadeMux I__3208 (
            .O(N__19727),
            .I(\POWERLED.N_84_f0_cascade_ ));
    CascadeMux I__3207 (
            .O(N__19724),
            .I(\POWERLED.N_108_f0_1_cascade_ ));
    InMux I__3206 (
            .O(N__19721),
            .I(N__19718));
    LocalMux I__3205 (
            .O(N__19718),
            .I(\POWERLED.dutycycle_eena_0 ));
    CascadeMux I__3204 (
            .O(N__19715),
            .I(\POWERLED.dutycycle_eena_0_cascade_ ));
    InMux I__3203 (
            .O(N__19712),
            .I(N__19706));
    InMux I__3202 (
            .O(N__19711),
            .I(N__19706));
    LocalMux I__3201 (
            .O(N__19706),
            .I(\POWERLED.dutycycleZ1Z_1 ));
    InMux I__3200 (
            .O(N__19703),
            .I(N__19700));
    LocalMux I__3199 (
            .O(N__19700),
            .I(\POWERLED.dutycycle_eena_1 ));
    CascadeMux I__3198 (
            .O(N__19697),
            .I(N__19694));
    InMux I__3197 (
            .O(N__19694),
            .I(N__19690));
    InMux I__3196 (
            .O(N__19693),
            .I(N__19687));
    LocalMux I__3195 (
            .O(N__19690),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    LocalMux I__3194 (
            .O(N__19687),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    CascadeMux I__3193 (
            .O(N__19682),
            .I(\POWERLED.func_state_0_sqmuxa_0_o2_xZ0Z1_cascade_ ));
    CascadeMux I__3192 (
            .O(N__19679),
            .I(\POWERLED.g1_1_cascade_ ));
    CascadeMux I__3191 (
            .O(N__19676),
            .I(\POWERLED.N_300_N_0_cascade_ ));
    InMux I__3190 (
            .O(N__19673),
            .I(N__19670));
    LocalMux I__3189 (
            .O(N__19670),
            .I(\POWERLED.N_4548_0 ));
    InMux I__3188 (
            .O(N__19667),
            .I(N__19664));
    LocalMux I__3187 (
            .O(N__19664),
            .I(\POWERLED.N_217_N_0 ));
    InMux I__3186 (
            .O(N__19661),
            .I(\POWERLED.un1_count_cry_12 ));
    InMux I__3185 (
            .O(N__19658),
            .I(\POWERLED.un1_count_cry_13 ));
    InMux I__3184 (
            .O(N__19655),
            .I(N__19652));
    LocalMux I__3183 (
            .O(N__19652),
            .I(N__19647));
    InMux I__3182 (
            .O(N__19651),
            .I(N__19644));
    InMux I__3181 (
            .O(N__19650),
            .I(N__19641));
    Span4Mux_v I__3180 (
            .O(N__19647),
            .I(N__19638));
    LocalMux I__3179 (
            .O(N__19644),
            .I(N__19633));
    LocalMux I__3178 (
            .O(N__19641),
            .I(N__19633));
    Odrv4 I__3177 (
            .O(N__19638),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv4 I__3176 (
            .O(N__19633),
            .I(\POWERLED.countZ0Z_15 ));
    InMux I__3175 (
            .O(N__19628),
            .I(\POWERLED.un1_count_cry_14 ));
    CascadeMux I__3174 (
            .O(N__19625),
            .I(N__19622));
    InMux I__3173 (
            .O(N__19622),
            .I(N__19616));
    InMux I__3172 (
            .O(N__19621),
            .I(N__19616));
    LocalMux I__3171 (
            .O(N__19616),
            .I(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ));
    InMux I__3170 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__3169 (
            .O(N__19610),
            .I(\POWERLED.count_0_9 ));
    InMux I__3168 (
            .O(N__19607),
            .I(N__19603));
    InMux I__3167 (
            .O(N__19606),
            .I(N__19600));
    LocalMux I__3166 (
            .O(N__19603),
            .I(\POWERLED.un1_count_cry_8_c_RNIIGZ0Z79 ));
    LocalMux I__3165 (
            .O(N__19600),
            .I(\POWERLED.un1_count_cry_8_c_RNIIGZ0Z79 ));
    InMux I__3164 (
            .O(N__19595),
            .I(N__19592));
    LocalMux I__3163 (
            .O(N__19592),
            .I(N__19588));
    InMux I__3162 (
            .O(N__19591),
            .I(N__19584));
    Span4Mux_v I__3161 (
            .O(N__19588),
            .I(N__19581));
    InMux I__3160 (
            .O(N__19587),
            .I(N__19578));
    LocalMux I__3159 (
            .O(N__19584),
            .I(N__19575));
    Odrv4 I__3158 (
            .O(N__19581),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__3157 (
            .O(N__19578),
            .I(\POWERLED.countZ0Z_9 ));
    Odrv4 I__3156 (
            .O(N__19575),
            .I(\POWERLED.countZ0Z_9 ));
    CascadeMux I__3155 (
            .O(N__19568),
            .I(\POWERLED.dutycycle_eena_1_cascade_ ));
    InMux I__3154 (
            .O(N__19565),
            .I(N__19562));
    LocalMux I__3153 (
            .O(N__19562),
            .I(\POWERLED.N_108_f0_1 ));
    InMux I__3152 (
            .O(N__19559),
            .I(\POWERLED.un1_count_cry_4 ));
    InMux I__3151 (
            .O(N__19556),
            .I(\POWERLED.un1_count_cry_5 ));
    InMux I__3150 (
            .O(N__19553),
            .I(N__19550));
    LocalMux I__3149 (
            .O(N__19550),
            .I(N__19545));
    InMux I__3148 (
            .O(N__19549),
            .I(N__19542));
    InMux I__3147 (
            .O(N__19548),
            .I(N__19539));
    Span4Mux_h I__3146 (
            .O(N__19545),
            .I(N__19532));
    LocalMux I__3145 (
            .O(N__19542),
            .I(N__19532));
    LocalMux I__3144 (
            .O(N__19539),
            .I(N__19532));
    Odrv4 I__3143 (
            .O(N__19532),
            .I(\POWERLED.countZ0Z_7 ));
    CascadeMux I__3142 (
            .O(N__19529),
            .I(N__19526));
    InMux I__3141 (
            .O(N__19526),
            .I(N__19520));
    InMux I__3140 (
            .O(N__19525),
            .I(N__19520));
    LocalMux I__3139 (
            .O(N__19520),
            .I(\POWERLED.un1_count_cry_6_c_RNIGCZ0Z59 ));
    InMux I__3138 (
            .O(N__19517),
            .I(\POWERLED.un1_count_cry_6 ));
    InMux I__3137 (
            .O(N__19514),
            .I(N__19510));
    InMux I__3136 (
            .O(N__19513),
            .I(N__19507));
    LocalMux I__3135 (
            .O(N__19510),
            .I(N__19503));
    LocalMux I__3134 (
            .O(N__19507),
            .I(N__19500));
    InMux I__3133 (
            .O(N__19506),
            .I(N__19497));
    Span4Mux_h I__3132 (
            .O(N__19503),
            .I(N__19492));
    Span4Mux_h I__3131 (
            .O(N__19500),
            .I(N__19492));
    LocalMux I__3130 (
            .O(N__19497),
            .I(\POWERLED.countZ0Z_8 ));
    Odrv4 I__3129 (
            .O(N__19492),
            .I(\POWERLED.countZ0Z_8 ));
    CascadeMux I__3128 (
            .O(N__19487),
            .I(N__19484));
    InMux I__3127 (
            .O(N__19484),
            .I(N__19478));
    InMux I__3126 (
            .O(N__19483),
            .I(N__19478));
    LocalMux I__3125 (
            .O(N__19478),
            .I(\POWERLED.un1_count_cry_7_c_RNIHEZ0Z69 ));
    InMux I__3124 (
            .O(N__19475),
            .I(\POWERLED.un1_count_cry_7 ));
    InMux I__3123 (
            .O(N__19472),
            .I(bfn_6_8_0_));
    InMux I__3122 (
            .O(N__19469),
            .I(N__19466));
    LocalMux I__3121 (
            .O(N__19466),
            .I(N__19461));
    CascadeMux I__3120 (
            .O(N__19465),
            .I(N__19458));
    CascadeMux I__3119 (
            .O(N__19464),
            .I(N__19455));
    Span4Mux_v I__3118 (
            .O(N__19461),
            .I(N__19452));
    InMux I__3117 (
            .O(N__19458),
            .I(N__19449));
    InMux I__3116 (
            .O(N__19455),
            .I(N__19446));
    Odrv4 I__3115 (
            .O(N__19452),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__3114 (
            .O(N__19449),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__3113 (
            .O(N__19446),
            .I(\POWERLED.countZ0Z_10 ));
    CascadeMux I__3112 (
            .O(N__19439),
            .I(N__19435));
    CascadeMux I__3111 (
            .O(N__19438),
            .I(N__19432));
    InMux I__3110 (
            .O(N__19435),
            .I(N__19429));
    InMux I__3109 (
            .O(N__19432),
            .I(N__19426));
    LocalMux I__3108 (
            .O(N__19429),
            .I(\POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ));
    LocalMux I__3107 (
            .O(N__19426),
            .I(\POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ));
    InMux I__3106 (
            .O(N__19421),
            .I(\POWERLED.un1_count_cry_9 ));
    InMux I__3105 (
            .O(N__19418),
            .I(N__19415));
    LocalMux I__3104 (
            .O(N__19415),
            .I(N__19412));
    Span4Mux_v I__3103 (
            .O(N__19412),
            .I(N__19407));
    InMux I__3102 (
            .O(N__19411),
            .I(N__19404));
    InMux I__3101 (
            .O(N__19410),
            .I(N__19401));
    Odrv4 I__3100 (
            .O(N__19407),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__3099 (
            .O(N__19404),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__3098 (
            .O(N__19401),
            .I(\POWERLED.countZ0Z_11 ));
    CascadeMux I__3097 (
            .O(N__19394),
            .I(N__19390));
    InMux I__3096 (
            .O(N__19393),
            .I(N__19385));
    InMux I__3095 (
            .O(N__19390),
            .I(N__19385));
    LocalMux I__3094 (
            .O(N__19385),
            .I(\POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7 ));
    InMux I__3093 (
            .O(N__19382),
            .I(\POWERLED.un1_count_cry_10 ));
    InMux I__3092 (
            .O(N__19379),
            .I(\POWERLED.un1_count_cry_11 ));
    CascadeMux I__3091 (
            .O(N__19376),
            .I(\POWERLED.un79_clk_100khzlt15_0_cascade_ ));
    SRMux I__3090 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__3089 (
            .O(N__19370),
            .I(N__19367));
    Span4Mux_v I__3088 (
            .O(N__19367),
            .I(N__19364));
    Span4Mux_s2_v I__3087 (
            .O(N__19364),
            .I(N__19361));
    Odrv4 I__3086 (
            .O(N__19361),
            .I(\POWERLED.pwm_out_1_sqmuxa ));
    InMux I__3085 (
            .O(N__19358),
            .I(N__19355));
    LocalMux I__3084 (
            .O(N__19355),
            .I(\POWERLED.un79_clk_100khzlto15_5 ));
    CascadeMux I__3083 (
            .O(N__19352),
            .I(\POWERLED.un79_clk_100khzlto15_6_cascade_ ));
    CascadeMux I__3082 (
            .O(N__19349),
            .I(\POWERLED.count_RNIZ0Z_15_cascade_ ));
    CascadeMux I__3081 (
            .O(N__19346),
            .I(N__19343));
    InMux I__3080 (
            .O(N__19343),
            .I(N__19337));
    InMux I__3079 (
            .O(N__19342),
            .I(N__19337));
    LocalMux I__3078 (
            .O(N__19337),
            .I(\POWERLED.N_8 ));
    InMux I__3077 (
            .O(N__19334),
            .I(N__19331));
    LocalMux I__3076 (
            .O(N__19331),
            .I(N__19328));
    Span4Mux_v I__3075 (
            .O(N__19328),
            .I(N__19323));
    InMux I__3074 (
            .O(N__19327),
            .I(N__19320));
    InMux I__3073 (
            .O(N__19326),
            .I(N__19317));
    Odrv4 I__3072 (
            .O(N__19323),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__3071 (
            .O(N__19320),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__3070 (
            .O(N__19317),
            .I(\POWERLED.countZ0Z_2 ));
    CascadeMux I__3069 (
            .O(N__19310),
            .I(N__19307));
    InMux I__3068 (
            .O(N__19307),
            .I(N__19301));
    InMux I__3067 (
            .O(N__19306),
            .I(N__19301));
    LocalMux I__3066 (
            .O(N__19301),
            .I(\POWERLED.un1_count_cry_1_c_RNIBZ0Z209 ));
    InMux I__3065 (
            .O(N__19298),
            .I(\POWERLED.un1_count_cry_1 ));
    InMux I__3064 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__3063 (
            .O(N__19292),
            .I(N__19289));
    Span4Mux_v I__3062 (
            .O(N__19289),
            .I(N__19284));
    InMux I__3061 (
            .O(N__19288),
            .I(N__19281));
    InMux I__3060 (
            .O(N__19287),
            .I(N__19278));
    Odrv4 I__3059 (
            .O(N__19284),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__3058 (
            .O(N__19281),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__3057 (
            .O(N__19278),
            .I(\POWERLED.countZ0Z_3 ));
    CascadeMux I__3056 (
            .O(N__19271),
            .I(N__19268));
    InMux I__3055 (
            .O(N__19268),
            .I(N__19262));
    InMux I__3054 (
            .O(N__19267),
            .I(N__19262));
    LocalMux I__3053 (
            .O(N__19262),
            .I(\POWERLED.un1_count_cry_2_c_RNICZ0Z419 ));
    InMux I__3052 (
            .O(N__19259),
            .I(\POWERLED.un1_count_cry_2 ));
    InMux I__3051 (
            .O(N__19256),
            .I(N__19253));
    LocalMux I__3050 (
            .O(N__19253),
            .I(N__19249));
    CascadeMux I__3049 (
            .O(N__19252),
            .I(N__19245));
    Span4Mux_v I__3048 (
            .O(N__19249),
            .I(N__19242));
    InMux I__3047 (
            .O(N__19248),
            .I(N__19239));
    InMux I__3046 (
            .O(N__19245),
            .I(N__19236));
    Odrv4 I__3045 (
            .O(N__19242),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__3044 (
            .O(N__19239),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__3043 (
            .O(N__19236),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__3042 (
            .O(N__19229),
            .I(N__19226));
    LocalMux I__3041 (
            .O(N__19226),
            .I(N__19223));
    Span4Mux_h I__3040 (
            .O(N__19223),
            .I(N__19219));
    InMux I__3039 (
            .O(N__19222),
            .I(N__19216));
    Odrv4 I__3038 (
            .O(N__19219),
            .I(\POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ));
    LocalMux I__3037 (
            .O(N__19216),
            .I(\POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ));
    InMux I__3036 (
            .O(N__19211),
            .I(\POWERLED.un1_count_cry_3 ));
    InMux I__3035 (
            .O(N__19208),
            .I(N__19204));
    InMux I__3034 (
            .O(N__19207),
            .I(N__19201));
    LocalMux I__3033 (
            .O(N__19204),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__3032 (
            .O(N__19201),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__3031 (
            .O(N__19196),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    CascadeMux I__3030 (
            .O(N__19193),
            .I(N__19189));
    InMux I__3029 (
            .O(N__19192),
            .I(N__19186));
    InMux I__3028 (
            .O(N__19189),
            .I(N__19183));
    LocalMux I__3027 (
            .O(N__19186),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    LocalMux I__3026 (
            .O(N__19183),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__3025 (
            .O(N__19178),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    CascadeMux I__3024 (
            .O(N__19175),
            .I(N__19171));
    InMux I__3023 (
            .O(N__19174),
            .I(N__19168));
    InMux I__3022 (
            .O(N__19171),
            .I(N__19165));
    LocalMux I__3021 (
            .O(N__19168),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__3020 (
            .O(N__19165),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__3019 (
            .O(N__19160),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__3018 (
            .O(N__19157),
            .I(N__19153));
    InMux I__3017 (
            .O(N__19156),
            .I(N__19150));
    LocalMux I__3016 (
            .O(N__19153),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    LocalMux I__3015 (
            .O(N__19150),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__3014 (
            .O(N__19145),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    InMux I__3013 (
            .O(N__19142),
            .I(bfn_6_5_0_));
    InMux I__3012 (
            .O(N__19139),
            .I(N__19135));
    InMux I__3011 (
            .O(N__19138),
            .I(N__19132));
    LocalMux I__3010 (
            .O(N__19135),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    LocalMux I__3009 (
            .O(N__19132),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    CEMux I__3008 (
            .O(N__19127),
            .I(N__19124));
    LocalMux I__3007 (
            .O(N__19124),
            .I(N__19121));
    Span4Mux_h I__3006 (
            .O(N__19121),
            .I(N__19118));
    Odrv4 I__3005 (
            .O(N__19118),
            .I(\RSMRST_PWRGD.N_27_2 ));
    SRMux I__3004 (
            .O(N__19115),
            .I(N__19111));
    SRMux I__3003 (
            .O(N__19114),
            .I(N__19108));
    LocalMux I__3002 (
            .O(N__19111),
            .I(N__19105));
    LocalMux I__3001 (
            .O(N__19108),
            .I(N__19101));
    Span4Mux_h I__3000 (
            .O(N__19105),
            .I(N__19098));
    SRMux I__2999 (
            .O(N__19104),
            .I(N__19095));
    Odrv4 I__2998 (
            .O(N__19101),
            .I(G_11));
    Odrv4 I__2997 (
            .O(N__19098),
            .I(G_11));
    LocalMux I__2996 (
            .O(N__19095),
            .I(G_11));
    CascadeMux I__2995 (
            .O(N__19088),
            .I(\POWERLED.un79_clk_100khzlto4_0_cascade_ ));
    InMux I__2994 (
            .O(N__19085),
            .I(N__19081));
    InMux I__2993 (
            .O(N__19084),
            .I(N__19078));
    LocalMux I__2992 (
            .O(N__19081),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__2991 (
            .O(N__19078),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    InMux I__2990 (
            .O(N__19073),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    CascadeMux I__2989 (
            .O(N__19070),
            .I(N__19066));
    InMux I__2988 (
            .O(N__19069),
            .I(N__19063));
    InMux I__2987 (
            .O(N__19066),
            .I(N__19060));
    LocalMux I__2986 (
            .O(N__19063),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__2985 (
            .O(N__19060),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__2984 (
            .O(N__19055),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__2983 (
            .O(N__19052),
            .I(N__19048));
    InMux I__2982 (
            .O(N__19051),
            .I(N__19045));
    LocalMux I__2981 (
            .O(N__19048),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__2980 (
            .O(N__19045),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    InMux I__2979 (
            .O(N__19040),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    InMux I__2978 (
            .O(N__19037),
            .I(N__19033));
    InMux I__2977 (
            .O(N__19036),
            .I(N__19030));
    LocalMux I__2976 (
            .O(N__19033),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    LocalMux I__2975 (
            .O(N__19030),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    InMux I__2974 (
            .O(N__19025),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__2973 (
            .O(N__19022),
            .I(N__19018));
    InMux I__2972 (
            .O(N__19021),
            .I(N__19015));
    LocalMux I__2971 (
            .O(N__19018),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__2970 (
            .O(N__19015),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__2969 (
            .O(N__19010),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__2968 (
            .O(N__19007),
            .I(N__19003));
    InMux I__2967 (
            .O(N__19006),
            .I(N__19000));
    LocalMux I__2966 (
            .O(N__19003),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__2965 (
            .O(N__19000),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    InMux I__2964 (
            .O(N__18995),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    CascadeMux I__2963 (
            .O(N__18992),
            .I(N__18988));
    InMux I__2962 (
            .O(N__18991),
            .I(N__18985));
    InMux I__2961 (
            .O(N__18988),
            .I(N__18982));
    LocalMux I__2960 (
            .O(N__18985),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__2959 (
            .O(N__18982),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__2958 (
            .O(N__18977),
            .I(bfn_6_4_0_));
    InMux I__2957 (
            .O(N__18974),
            .I(N__18970));
    InMux I__2956 (
            .O(N__18973),
            .I(N__18967));
    LocalMux I__2955 (
            .O(N__18970),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    LocalMux I__2954 (
            .O(N__18967),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__2953 (
            .O(N__18962),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__2952 (
            .O(N__18959),
            .I(N__18955));
    InMux I__2951 (
            .O(N__18958),
            .I(N__18952));
    LocalMux I__2950 (
            .O(N__18955),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    LocalMux I__2949 (
            .O(N__18952),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    InMux I__2948 (
            .O(N__18947),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__2947 (
            .O(N__18944),
            .I(N__18941));
    LocalMux I__2946 (
            .O(N__18941),
            .I(\PCH_PWRGD.un2_count_1_axb_2 ));
    SRMux I__2945 (
            .O(N__18938),
            .I(N__18932));
    SRMux I__2944 (
            .O(N__18937),
            .I(N__18929));
    SRMux I__2943 (
            .O(N__18936),
            .I(N__18923));
    SRMux I__2942 (
            .O(N__18935),
            .I(N__18920));
    LocalMux I__2941 (
            .O(N__18932),
            .I(N__18917));
    LocalMux I__2940 (
            .O(N__18929),
            .I(N__18914));
    SRMux I__2939 (
            .O(N__18928),
            .I(N__18910));
    SRMux I__2938 (
            .O(N__18927),
            .I(N__18907));
    InMux I__2937 (
            .O(N__18926),
            .I(N__18904));
    LocalMux I__2936 (
            .O(N__18923),
            .I(N__18901));
    LocalMux I__2935 (
            .O(N__18920),
            .I(N__18898));
    IoSpan4Mux I__2934 (
            .O(N__18917),
            .I(N__18893));
    Span4Mux_v I__2933 (
            .O(N__18914),
            .I(N__18893));
    SRMux I__2932 (
            .O(N__18913),
            .I(N__18890));
    LocalMux I__2931 (
            .O(N__18910),
            .I(N__18883));
    LocalMux I__2930 (
            .O(N__18907),
            .I(N__18883));
    LocalMux I__2929 (
            .O(N__18904),
            .I(N__18883));
    Span4Mux_s1_v I__2928 (
            .O(N__18901),
            .I(N__18876));
    Span4Mux_h I__2927 (
            .O(N__18898),
            .I(N__18867));
    Span4Mux_s1_v I__2926 (
            .O(N__18893),
            .I(N__18867));
    LocalMux I__2925 (
            .O(N__18890),
            .I(N__18867));
    Span4Mux_v I__2924 (
            .O(N__18883),
            .I(N__18867));
    InMux I__2923 (
            .O(N__18882),
            .I(N__18860));
    InMux I__2922 (
            .O(N__18881),
            .I(N__18860));
    InMux I__2921 (
            .O(N__18880),
            .I(N__18860));
    SRMux I__2920 (
            .O(N__18879),
            .I(N__18857));
    Sp12to4 I__2919 (
            .O(N__18876),
            .I(N__18850));
    Sp12to4 I__2918 (
            .O(N__18867),
            .I(N__18850));
    LocalMux I__2917 (
            .O(N__18860),
            .I(N__18850));
    LocalMux I__2916 (
            .O(N__18857),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv12 I__2915 (
            .O(N__18850),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    CascadeMux I__2914 (
            .O(N__18845),
            .I(N__18842));
    InMux I__2913 (
            .O(N__18842),
            .I(N__18833));
    InMux I__2912 (
            .O(N__18841),
            .I(N__18833));
    InMux I__2911 (
            .O(N__18840),
            .I(N__18833));
    LocalMux I__2910 (
            .O(N__18833),
            .I(\PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSCZ0 ));
    InMux I__2909 (
            .O(N__18830),
            .I(N__18824));
    InMux I__2908 (
            .O(N__18829),
            .I(N__18824));
    LocalMux I__2907 (
            .O(N__18824),
            .I(\PCH_PWRGD.count_0_2 ));
    CascadeMux I__2906 (
            .O(N__18821),
            .I(\PCH_PWRGD.count_rst_12_cascade_ ));
    InMux I__2905 (
            .O(N__18818),
            .I(N__18815));
    LocalMux I__2904 (
            .O(N__18815),
            .I(N__18811));
    InMux I__2903 (
            .O(N__18814),
            .I(N__18808));
    Span4Mux_s1_v I__2902 (
            .O(N__18811),
            .I(N__18805));
    LocalMux I__2901 (
            .O(N__18808),
            .I(N__18802));
    Odrv4 I__2900 (
            .O(N__18805),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    Odrv12 I__2899 (
            .O(N__18802),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__2898 (
            .O(N__18797),
            .I(N__18794));
    LocalMux I__2897 (
            .O(N__18794),
            .I(N__18791));
    Span4Mux_v I__2896 (
            .O(N__18791),
            .I(N__18788));
    Odrv4 I__2895 (
            .O(N__18788),
            .I(\PCH_PWRGD.un12_clk_100khz_3 ));
    InMux I__2894 (
            .O(N__18785),
            .I(N__18782));
    LocalMux I__2893 (
            .O(N__18782),
            .I(\PCH_PWRGD.count_0_12 ));
    InMux I__2892 (
            .O(N__18779),
            .I(N__18776));
    LocalMux I__2891 (
            .O(N__18776),
            .I(N__18772));
    InMux I__2890 (
            .O(N__18775),
            .I(N__18769));
    Odrv4 I__2889 (
            .O(N__18772),
            .I(\PCH_PWRGD.count_rst_2 ));
    LocalMux I__2888 (
            .O(N__18769),
            .I(\PCH_PWRGD.count_rst_2 ));
    InMux I__2887 (
            .O(N__18764),
            .I(N__18761));
    LocalMux I__2886 (
            .O(N__18761),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    InMux I__2885 (
            .O(N__18758),
            .I(N__18751));
    InMux I__2884 (
            .O(N__18757),
            .I(N__18751));
    InMux I__2883 (
            .O(N__18756),
            .I(N__18748));
    LocalMux I__2882 (
            .O(N__18751),
            .I(N__18745));
    LocalMux I__2881 (
            .O(N__18748),
            .I(\PCH_PWRGD.count_rst_4 ));
    Odrv12 I__2880 (
            .O(N__18745),
            .I(\PCH_PWRGD.count_rst_4 ));
    InMux I__2879 (
            .O(N__18740),
            .I(N__18737));
    LocalMux I__2878 (
            .O(N__18737),
            .I(N__18733));
    InMux I__2877 (
            .O(N__18736),
            .I(N__18730));
    Span4Mux_s1_v I__2876 (
            .O(N__18733),
            .I(N__18727));
    LocalMux I__2875 (
            .O(N__18730),
            .I(\PCH_PWRGD.count_0_10 ));
    Odrv4 I__2874 (
            .O(N__18727),
            .I(\PCH_PWRGD.count_0_10 ));
    CascadeMux I__2873 (
            .O(N__18722),
            .I(\PCH_PWRGD.countZ0Z_12_cascade_ ));
    CEMux I__2872 (
            .O(N__18719),
            .I(N__18710));
    CEMux I__2871 (
            .O(N__18718),
            .I(N__18707));
    CEMux I__2870 (
            .O(N__18717),
            .I(N__18704));
    CEMux I__2869 (
            .O(N__18716),
            .I(N__18698));
    CascadeMux I__2868 (
            .O(N__18715),
            .I(N__18694));
    CEMux I__2867 (
            .O(N__18714),
            .I(N__18685));
    CascadeMux I__2866 (
            .O(N__18713),
            .I(N__18682));
    LocalMux I__2865 (
            .O(N__18710),
            .I(N__18673));
    LocalMux I__2864 (
            .O(N__18707),
            .I(N__18670));
    LocalMux I__2863 (
            .O(N__18704),
            .I(N__18667));
    InMux I__2862 (
            .O(N__18703),
            .I(N__18658));
    InMux I__2861 (
            .O(N__18702),
            .I(N__18658));
    CEMux I__2860 (
            .O(N__18701),
            .I(N__18655));
    LocalMux I__2859 (
            .O(N__18698),
            .I(N__18652));
    CEMux I__2858 (
            .O(N__18697),
            .I(N__18647));
    InMux I__2857 (
            .O(N__18694),
            .I(N__18647));
    InMux I__2856 (
            .O(N__18693),
            .I(N__18642));
    InMux I__2855 (
            .O(N__18692),
            .I(N__18642));
    InMux I__2854 (
            .O(N__18691),
            .I(N__18637));
    InMux I__2853 (
            .O(N__18690),
            .I(N__18637));
    InMux I__2852 (
            .O(N__18689),
            .I(N__18629));
    InMux I__2851 (
            .O(N__18688),
            .I(N__18629));
    LocalMux I__2850 (
            .O(N__18685),
            .I(N__18626));
    InMux I__2849 (
            .O(N__18682),
            .I(N__18623));
    InMux I__2848 (
            .O(N__18681),
            .I(N__18618));
    InMux I__2847 (
            .O(N__18680),
            .I(N__18618));
    InMux I__2846 (
            .O(N__18679),
            .I(N__18609));
    InMux I__2845 (
            .O(N__18678),
            .I(N__18609));
    InMux I__2844 (
            .O(N__18677),
            .I(N__18609));
    InMux I__2843 (
            .O(N__18676),
            .I(N__18609));
    Span4Mux_s3_v I__2842 (
            .O(N__18673),
            .I(N__18606));
    Span4Mux_v I__2841 (
            .O(N__18670),
            .I(N__18601));
    Span4Mux_s3_v I__2840 (
            .O(N__18667),
            .I(N__18601));
    CEMux I__2839 (
            .O(N__18666),
            .I(N__18592));
    InMux I__2838 (
            .O(N__18665),
            .I(N__18592));
    InMux I__2837 (
            .O(N__18664),
            .I(N__18592));
    InMux I__2836 (
            .O(N__18663),
            .I(N__18592));
    LocalMux I__2835 (
            .O(N__18658),
            .I(N__18589));
    LocalMux I__2834 (
            .O(N__18655),
            .I(N__18586));
    Span4Mux_h I__2833 (
            .O(N__18652),
            .I(N__18577));
    LocalMux I__2832 (
            .O(N__18647),
            .I(N__18577));
    LocalMux I__2831 (
            .O(N__18642),
            .I(N__18577));
    LocalMux I__2830 (
            .O(N__18637),
            .I(N__18577));
    InMux I__2829 (
            .O(N__18636),
            .I(N__18570));
    InMux I__2828 (
            .O(N__18635),
            .I(N__18570));
    InMux I__2827 (
            .O(N__18634),
            .I(N__18570));
    LocalMux I__2826 (
            .O(N__18629),
            .I(N__18567));
    Span4Mux_s1_v I__2825 (
            .O(N__18626),
            .I(N__18560));
    LocalMux I__2824 (
            .O(N__18623),
            .I(N__18560));
    LocalMux I__2823 (
            .O(N__18618),
            .I(N__18560));
    LocalMux I__2822 (
            .O(N__18609),
            .I(N__18557));
    Span4Mux_h I__2821 (
            .O(N__18606),
            .I(N__18554));
    Span4Mux_h I__2820 (
            .O(N__18601),
            .I(N__18547));
    LocalMux I__2819 (
            .O(N__18592),
            .I(N__18547));
    Span4Mux_s3_v I__2818 (
            .O(N__18589),
            .I(N__18547));
    Span4Mux_s0_v I__2817 (
            .O(N__18586),
            .I(N__18542));
    Span4Mux_h I__2816 (
            .O(N__18577),
            .I(N__18542));
    LocalMux I__2815 (
            .O(N__18570),
            .I(N__18539));
    Span4Mux_h I__2814 (
            .O(N__18567),
            .I(N__18532));
    Span4Mux_h I__2813 (
            .O(N__18560),
            .I(N__18532));
    Span4Mux_h I__2812 (
            .O(N__18557),
            .I(N__18532));
    Odrv4 I__2811 (
            .O(N__18554),
            .I(\PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0 ));
    Odrv4 I__2810 (
            .O(N__18547),
            .I(\PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0 ));
    Odrv4 I__2809 (
            .O(N__18542),
            .I(\PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0 ));
    Odrv4 I__2808 (
            .O(N__18539),
            .I(\PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0 ));
    Odrv4 I__2807 (
            .O(N__18532),
            .I(\PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0 ));
    InMux I__2806 (
            .O(N__18521),
            .I(N__18518));
    LocalMux I__2805 (
            .O(N__18518),
            .I(N__18515));
    Span4Mux_h I__2804 (
            .O(N__18515),
            .I(N__18512));
    Odrv4 I__2803 (
            .O(N__18512),
            .I(\PCH_PWRGD.un12_clk_100khz_2 ));
    CascadeMux I__2802 (
            .O(N__18509),
            .I(N__18505));
    InMux I__2801 (
            .O(N__18508),
            .I(N__18502));
    InMux I__2800 (
            .O(N__18505),
            .I(N__18499));
    LocalMux I__2799 (
            .O(N__18502),
            .I(N__18494));
    LocalMux I__2798 (
            .O(N__18499),
            .I(N__18494));
    Span4Mux_v I__2797 (
            .O(N__18494),
            .I(N__18491));
    Odrv4 I__2796 (
            .O(N__18491),
            .I(\RSMRST_PWRGD.N_256_i ));
    InMux I__2795 (
            .O(N__18488),
            .I(N__18484));
    InMux I__2794 (
            .O(N__18487),
            .I(N__18481));
    LocalMux I__2793 (
            .O(N__18484),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__2792 (
            .O(N__18481),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__2791 (
            .O(N__18476),
            .I(N__18472));
    InMux I__2790 (
            .O(N__18475),
            .I(N__18469));
    LocalMux I__2789 (
            .O(N__18472),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__2788 (
            .O(N__18469),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    InMux I__2787 (
            .O(N__18464),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    InMux I__2786 (
            .O(N__18461),
            .I(N__18458));
    LocalMux I__2785 (
            .O(N__18458),
            .I(N__18455));
    Odrv4 I__2784 (
            .O(N__18455),
            .I(\POWERLED.mult1_un75_sum_i ));
    CascadeMux I__2783 (
            .O(N__18452),
            .I(N__18449));
    InMux I__2782 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__2781 (
            .O(N__18446),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__2780 (
            .O(N__18443),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    CascadeMux I__2779 (
            .O(N__18440),
            .I(N__18437));
    InMux I__2778 (
            .O(N__18437),
            .I(N__18434));
    LocalMux I__2777 (
            .O(N__18434),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__2776 (
            .O(N__18431),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    InMux I__2775 (
            .O(N__18428),
            .I(N__18425));
    LocalMux I__2774 (
            .O(N__18425),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__2773 (
            .O(N__18422),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__2772 (
            .O(N__18419),
            .I(N__18416));
    LocalMux I__2771 (
            .O(N__18416),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__2770 (
            .O(N__18413),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    CascadeMux I__2769 (
            .O(N__18410),
            .I(N__18407));
    InMux I__2768 (
            .O(N__18407),
            .I(N__18404));
    LocalMux I__2767 (
            .O(N__18404),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__2766 (
            .O(N__18401),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__2765 (
            .O(N__18398),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    InMux I__2764 (
            .O(N__18395),
            .I(N__18392));
    LocalMux I__2763 (
            .O(N__18392),
            .I(N__18388));
    CascadeMux I__2762 (
            .O(N__18391),
            .I(N__18384));
    Span4Mux_h I__2761 (
            .O(N__18388),
            .I(N__18379));
    InMux I__2760 (
            .O(N__18387),
            .I(N__18376));
    InMux I__2759 (
            .O(N__18384),
            .I(N__18369));
    InMux I__2758 (
            .O(N__18383),
            .I(N__18369));
    InMux I__2757 (
            .O(N__18382),
            .I(N__18369));
    Odrv4 I__2756 (
            .O(N__18379),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2755 (
            .O(N__18376),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2754 (
            .O(N__18369),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    CascadeMux I__2753 (
            .O(N__18362),
            .I(N__18358));
    CascadeMux I__2752 (
            .O(N__18361),
            .I(N__18354));
    InMux I__2751 (
            .O(N__18358),
            .I(N__18347));
    InMux I__2750 (
            .O(N__18357),
            .I(N__18347));
    InMux I__2749 (
            .O(N__18354),
            .I(N__18347));
    LocalMux I__2748 (
            .O(N__18347),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    InMux I__2747 (
            .O(N__18344),
            .I(N__18341));
    LocalMux I__2746 (
            .O(N__18341),
            .I(\POWERLED.mult1_un61_sum_i ));
    InMux I__2745 (
            .O(N__18338),
            .I(\POWERLED.mult1_un68_sum_cry_2_c ));
    CascadeMux I__2744 (
            .O(N__18335),
            .I(N__18332));
    InMux I__2743 (
            .O(N__18332),
            .I(N__18329));
    LocalMux I__2742 (
            .O(N__18329),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__2741 (
            .O(N__18326),
            .I(\POWERLED.mult1_un68_sum_cry_3_c ));
    InMux I__2740 (
            .O(N__18323),
            .I(N__18320));
    LocalMux I__2739 (
            .O(N__18320),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__2738 (
            .O(N__18317),
            .I(\POWERLED.mult1_un68_sum_cry_4_c ));
    InMux I__2737 (
            .O(N__18314),
            .I(N__18310));
    CascadeMux I__2736 (
            .O(N__18313),
            .I(N__18306));
    LocalMux I__2735 (
            .O(N__18310),
            .I(N__18302));
    InMux I__2734 (
            .O(N__18309),
            .I(N__18297));
    InMux I__2733 (
            .O(N__18306),
            .I(N__18297));
    InMux I__2732 (
            .O(N__18305),
            .I(N__18294));
    Odrv4 I__2731 (
            .O(N__18302),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__2730 (
            .O(N__18297),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__2729 (
            .O(N__18294),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__2728 (
            .O(N__18287),
            .I(N__18284));
    InMux I__2727 (
            .O(N__18284),
            .I(N__18281));
    LocalMux I__2726 (
            .O(N__18281),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__2725 (
            .O(N__18278),
            .I(\POWERLED.mult1_un68_sum_cry_5_c ));
    InMux I__2724 (
            .O(N__18275),
            .I(N__18272));
    LocalMux I__2723 (
            .O(N__18272),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    CascadeMux I__2722 (
            .O(N__18269),
            .I(N__18265));
    CascadeMux I__2721 (
            .O(N__18268),
            .I(N__18261));
    InMux I__2720 (
            .O(N__18265),
            .I(N__18254));
    InMux I__2719 (
            .O(N__18264),
            .I(N__18254));
    InMux I__2718 (
            .O(N__18261),
            .I(N__18254));
    LocalMux I__2717 (
            .O(N__18254),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    InMux I__2716 (
            .O(N__18251),
            .I(\POWERLED.mult1_un68_sum_cry_6_c ));
    CascadeMux I__2715 (
            .O(N__18248),
            .I(N__18245));
    InMux I__2714 (
            .O(N__18245),
            .I(N__18242));
    LocalMux I__2713 (
            .O(N__18242),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__2712 (
            .O(N__18239),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__2711 (
            .O(N__18236),
            .I(\POWERLED.mult1_un68_sum_s_8_cascade_ ));
    InMux I__2710 (
            .O(N__18233),
            .I(N__18229));
    InMux I__2709 (
            .O(N__18232),
            .I(N__18226));
    LocalMux I__2708 (
            .O(N__18229),
            .I(N__18223));
    LocalMux I__2707 (
            .O(N__18226),
            .I(\POWERLED.mult1_un82_sum ));
    Odrv12 I__2706 (
            .O(N__18223),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__2705 (
            .O(N__18218),
            .I(\POWERLED.un1_dutycycle_53_cry_14 ));
    InMux I__2704 (
            .O(N__18215),
            .I(bfn_5_13_0_));
    InMux I__2703 (
            .O(N__18212),
            .I(\POWERLED.CO2 ));
    InMux I__2702 (
            .O(N__18209),
            .I(N__18206));
    LocalMux I__2701 (
            .O(N__18206),
            .I(N__18203));
    Span4Mux_s3_v I__2700 (
            .O(N__18203),
            .I(N__18200));
    Odrv4 I__2699 (
            .O(N__18200),
            .I(\POWERLED.mult1_un82_sum_i ));
    CascadeMux I__2698 (
            .O(N__18197),
            .I(N__18194));
    InMux I__2697 (
            .O(N__18194),
            .I(N__18191));
    LocalMux I__2696 (
            .O(N__18191),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    InMux I__2695 (
            .O(N__18188),
            .I(N__18184));
    InMux I__2694 (
            .O(N__18187),
            .I(N__18181));
    LocalMux I__2693 (
            .O(N__18184),
            .I(N__18178));
    LocalMux I__2692 (
            .O(N__18181),
            .I(\POWERLED.mult1_un61_sum ));
    Odrv4 I__2691 (
            .O(N__18178),
            .I(\POWERLED.mult1_un61_sum ));
    CascadeMux I__2690 (
            .O(N__18173),
            .I(N__18170));
    InMux I__2689 (
            .O(N__18170),
            .I(N__18164));
    InMux I__2688 (
            .O(N__18169),
            .I(N__18164));
    LocalMux I__2687 (
            .O(N__18164),
            .I(\POWERLED.CO2_THRU_CO ));
    InMux I__2686 (
            .O(N__18161),
            .I(N__18157));
    InMux I__2685 (
            .O(N__18160),
            .I(N__18154));
    LocalMux I__2684 (
            .O(N__18157),
            .I(N__18151));
    LocalMux I__2683 (
            .O(N__18154),
            .I(N__18148));
    Span4Mux_s2_v I__2682 (
            .O(N__18151),
            .I(N__18145));
    Span4Mux_s1_v I__2681 (
            .O(N__18148),
            .I(N__18142));
    Span4Mux_h I__2680 (
            .O(N__18145),
            .I(N__18139));
    Span4Mux_v I__2679 (
            .O(N__18142),
            .I(N__18136));
    Odrv4 I__2678 (
            .O(N__18139),
            .I(\POWERLED.mult1_un103_sum ));
    Odrv4 I__2677 (
            .O(N__18136),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__2676 (
            .O(N__18131),
            .I(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ));
    InMux I__2675 (
            .O(N__18128),
            .I(N__18125));
    LocalMux I__2674 (
            .O(N__18125),
            .I(N__18121));
    InMux I__2673 (
            .O(N__18124),
            .I(N__18118));
    Span4Mux_s1_v I__2672 (
            .O(N__18121),
            .I(N__18113));
    LocalMux I__2671 (
            .O(N__18118),
            .I(N__18113));
    Span4Mux_v I__2670 (
            .O(N__18113),
            .I(N__18110));
    Odrv4 I__2669 (
            .O(N__18110),
            .I(\POWERLED.mult1_un96_sum ));
    InMux I__2668 (
            .O(N__18107),
            .I(\POWERLED.un1_dutycycle_53_cry_6_cZ0 ));
    InMux I__2667 (
            .O(N__18104),
            .I(N__18101));
    LocalMux I__2666 (
            .O(N__18101),
            .I(N__18097));
    InMux I__2665 (
            .O(N__18100),
            .I(N__18094));
    Span4Mux_h I__2664 (
            .O(N__18097),
            .I(N__18089));
    LocalMux I__2663 (
            .O(N__18094),
            .I(N__18089));
    Span4Mux_s2_v I__2662 (
            .O(N__18089),
            .I(N__18086));
    Odrv4 I__2661 (
            .O(N__18086),
            .I(\POWERLED.mult1_un89_sum ));
    InMux I__2660 (
            .O(N__18083),
            .I(bfn_5_12_0_));
    InMux I__2659 (
            .O(N__18080),
            .I(\POWERLED.un1_dutycycle_53_cry_8_cZ0 ));
    InMux I__2658 (
            .O(N__18077),
            .I(\POWERLED.un1_dutycycle_53_cry_9_cZ0 ));
    InMux I__2657 (
            .O(N__18074),
            .I(N__18071));
    LocalMux I__2656 (
            .O(N__18071),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_14 ));
    InMux I__2655 (
            .O(N__18068),
            .I(\POWERLED.un1_dutycycle_53_cry_10 ));
    InMux I__2654 (
            .O(N__18065),
            .I(\POWERLED.un1_dutycycle_53_cry_11 ));
    CascadeMux I__2653 (
            .O(N__18062),
            .I(N__18058));
    InMux I__2652 (
            .O(N__18061),
            .I(N__18055));
    InMux I__2651 (
            .O(N__18058),
            .I(N__18052));
    LocalMux I__2650 (
            .O(N__18055),
            .I(\POWERLED.mult1_un54_sum ));
    LocalMux I__2649 (
            .O(N__18052),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__2648 (
            .O(N__18047),
            .I(\POWERLED.un1_dutycycle_53_cry_12 ));
    InMux I__2647 (
            .O(N__18044),
            .I(\POWERLED.un1_dutycycle_53_cry_13 ));
    InMux I__2646 (
            .O(N__18041),
            .I(N__18038));
    LocalMux I__2645 (
            .O(N__18038),
            .I(N__18035));
    Odrv12 I__2644 (
            .O(N__18035),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__2643 (
            .O(N__18032),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    CascadeMux I__2642 (
            .O(N__18029),
            .I(N__18024));
    InMux I__2641 (
            .O(N__18028),
            .I(N__18017));
    InMux I__2640 (
            .O(N__18027),
            .I(N__18017));
    InMux I__2639 (
            .O(N__18024),
            .I(N__18012));
    InMux I__2638 (
            .O(N__18023),
            .I(N__18012));
    InMux I__2637 (
            .O(N__18022),
            .I(N__18009));
    LocalMux I__2636 (
            .O(N__18017),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__2635 (
            .O(N__18012),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__2634 (
            .O(N__18009),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    InMux I__2633 (
            .O(N__18002),
            .I(N__17999));
    LocalMux I__2632 (
            .O(N__17999),
            .I(N__17996));
    Span4Mux_v I__2631 (
            .O(N__17996),
            .I(N__17993));
    Span4Mux_h I__2630 (
            .O(N__17993),
            .I(N__17989));
    InMux I__2629 (
            .O(N__17992),
            .I(N__17986));
    Odrv4 I__2628 (
            .O(N__17989),
            .I(\POWERLED.mult1_un145_sum ));
    LocalMux I__2627 (
            .O(N__17986),
            .I(\POWERLED.mult1_un145_sum ));
    InMux I__2626 (
            .O(N__17981),
            .I(N__17978));
    LocalMux I__2625 (
            .O(N__17978),
            .I(N__17974));
    InMux I__2624 (
            .O(N__17977),
            .I(N__17971));
    Span4Mux_v I__2623 (
            .O(N__17974),
            .I(N__17968));
    LocalMux I__2622 (
            .O(N__17971),
            .I(N__17965));
    Odrv4 I__2621 (
            .O(N__17968),
            .I(\POWERLED.mult1_un138_sum ));
    Odrv12 I__2620 (
            .O(N__17965),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__2619 (
            .O(N__17960),
            .I(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ));
    InMux I__2618 (
            .O(N__17957),
            .I(N__17954));
    LocalMux I__2617 (
            .O(N__17954),
            .I(N__17950));
    InMux I__2616 (
            .O(N__17953),
            .I(N__17947));
    Span4Mux_v I__2615 (
            .O(N__17950),
            .I(N__17942));
    LocalMux I__2614 (
            .O(N__17947),
            .I(N__17942));
    Odrv4 I__2613 (
            .O(N__17942),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__2612 (
            .O(N__17939),
            .I(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ));
    InMux I__2611 (
            .O(N__17936),
            .I(N__17932));
    InMux I__2610 (
            .O(N__17935),
            .I(N__17929));
    LocalMux I__2609 (
            .O(N__17932),
            .I(N__17924));
    LocalMux I__2608 (
            .O(N__17929),
            .I(N__17924));
    Span4Mux_v I__2607 (
            .O(N__17924),
            .I(N__17921));
    Odrv4 I__2606 (
            .O(N__17921),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__2605 (
            .O(N__17918),
            .I(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ));
    InMux I__2604 (
            .O(N__17915),
            .I(N__17911));
    InMux I__2603 (
            .O(N__17914),
            .I(N__17908));
    LocalMux I__2602 (
            .O(N__17911),
            .I(N__17905));
    LocalMux I__2601 (
            .O(N__17908),
            .I(N__17902));
    Span4Mux_v I__2600 (
            .O(N__17905),
            .I(N__17899));
    Span4Mux_v I__2599 (
            .O(N__17902),
            .I(N__17896));
    Odrv4 I__2598 (
            .O(N__17899),
            .I(\POWERLED.mult1_un117_sum ));
    Odrv4 I__2597 (
            .O(N__17896),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__2596 (
            .O(N__17891),
            .I(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ));
    InMux I__2595 (
            .O(N__17888),
            .I(N__17885));
    LocalMux I__2594 (
            .O(N__17885),
            .I(N__17881));
    InMux I__2593 (
            .O(N__17884),
            .I(N__17878));
    Span4Mux_s2_h I__2592 (
            .O(N__17881),
            .I(N__17873));
    LocalMux I__2591 (
            .O(N__17878),
            .I(N__17873));
    Span4Mux_v I__2590 (
            .O(N__17873),
            .I(N__17870));
    Odrv4 I__2589 (
            .O(N__17870),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__2588 (
            .O(N__17867),
            .I(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ));
    InMux I__2587 (
            .O(N__17864),
            .I(N__17861));
    LocalMux I__2586 (
            .O(N__17861),
            .I(\POWERLED.count_0_8 ));
    InMux I__2585 (
            .O(N__17858),
            .I(N__17855));
    LocalMux I__2584 (
            .O(N__17855),
            .I(N__17852));
    Odrv4 I__2583 (
            .O(N__17852),
            .I(\POWERLED.count_0_10 ));
    CascadeMux I__2582 (
            .O(N__17849),
            .I(N__17846));
    InMux I__2581 (
            .O(N__17846),
            .I(N__17843));
    LocalMux I__2580 (
            .O(N__17843),
            .I(\POWERLED.mult1_un145_sum_i ));
    InMux I__2579 (
            .O(N__17840),
            .I(N__17837));
    LocalMux I__2578 (
            .O(N__17837),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    InMux I__2577 (
            .O(N__17834),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    InMux I__2576 (
            .O(N__17831),
            .I(N__17828));
    LocalMux I__2575 (
            .O(N__17828),
            .I(N__17825));
    Odrv12 I__2574 (
            .O(N__17825),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    CascadeMux I__2573 (
            .O(N__17822),
            .I(N__17819));
    InMux I__2572 (
            .O(N__17819),
            .I(N__17816));
    LocalMux I__2571 (
            .O(N__17816),
            .I(N__17813));
    Odrv4 I__2570 (
            .O(N__17813),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__2569 (
            .O(N__17810),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    InMux I__2568 (
            .O(N__17807),
            .I(N__17804));
    LocalMux I__2567 (
            .O(N__17804),
            .I(N__17801));
    Odrv12 I__2566 (
            .O(N__17801),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__2565 (
            .O(N__17798),
            .I(N__17795));
    LocalMux I__2564 (
            .O(N__17795),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    InMux I__2563 (
            .O(N__17792),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    CascadeMux I__2562 (
            .O(N__17789),
            .I(N__17785));
    InMux I__2561 (
            .O(N__17788),
            .I(N__17780));
    InMux I__2560 (
            .O(N__17785),
            .I(N__17780));
    LocalMux I__2559 (
            .O(N__17780),
            .I(N__17774));
    InMux I__2558 (
            .O(N__17779),
            .I(N__17769));
    InMux I__2557 (
            .O(N__17778),
            .I(N__17769));
    InMux I__2556 (
            .O(N__17777),
            .I(N__17766));
    Odrv12 I__2555 (
            .O(N__17774),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__2554 (
            .O(N__17769),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__2553 (
            .O(N__17766),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    CascadeMux I__2552 (
            .O(N__17759),
            .I(N__17756));
    InMux I__2551 (
            .O(N__17756),
            .I(N__17753));
    LocalMux I__2550 (
            .O(N__17753),
            .I(N__17750));
    Odrv12 I__2549 (
            .O(N__17750),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    CascadeMux I__2548 (
            .O(N__17747),
            .I(N__17744));
    InMux I__2547 (
            .O(N__17744),
            .I(N__17741));
    LocalMux I__2546 (
            .O(N__17741),
            .I(N__17738));
    Odrv4 I__2545 (
            .O(N__17738),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__2544 (
            .O(N__17735),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    CascadeMux I__2543 (
            .O(N__17732),
            .I(N__17728));
    InMux I__2542 (
            .O(N__17731),
            .I(N__17720));
    InMux I__2541 (
            .O(N__17728),
            .I(N__17720));
    InMux I__2540 (
            .O(N__17727),
            .I(N__17720));
    LocalMux I__2539 (
            .O(N__17720),
            .I(N__17717));
    Span4Mux_h I__2538 (
            .O(N__17717),
            .I(N__17714));
    Odrv4 I__2537 (
            .O(N__17714),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    CascadeMux I__2536 (
            .O(N__17711),
            .I(N__17708));
    InMux I__2535 (
            .O(N__17708),
            .I(N__17705));
    LocalMux I__2534 (
            .O(N__17705),
            .I(N__17702));
    Odrv12 I__2533 (
            .O(N__17702),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    InMux I__2532 (
            .O(N__17699),
            .I(N__17696));
    LocalMux I__2531 (
            .O(N__17696),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__2530 (
            .O(N__17693),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__2529 (
            .O(N__17690),
            .I(N__17687));
    LocalMux I__2528 (
            .O(N__17687),
            .I(\POWERLED.count_0_11 ));
    InMux I__2527 (
            .O(N__17684),
            .I(N__17681));
    LocalMux I__2526 (
            .O(N__17681),
            .I(\POWERLED.count_0_3 ));
    InMux I__2525 (
            .O(N__17678),
            .I(N__17675));
    LocalMux I__2524 (
            .O(N__17675),
            .I(\POWERLED.count_0_15 ));
    InMux I__2523 (
            .O(N__17672),
            .I(N__17669));
    LocalMux I__2522 (
            .O(N__17669),
            .I(\POWERLED.count_0_7 ));
    InMux I__2521 (
            .O(N__17666),
            .I(N__17663));
    LocalMux I__2520 (
            .O(N__17663),
            .I(\PCH_PWRGD.count_0_6 ));
    InMux I__2519 (
            .O(N__17660),
            .I(N__17657));
    LocalMux I__2518 (
            .O(N__17657),
            .I(N__17654));
    Odrv4 I__2517 (
            .O(N__17654),
            .I(\PCH_PWRGD.un2_count_1_axb_10 ));
    InMux I__2516 (
            .O(N__17651),
            .I(N__17647));
    CascadeMux I__2515 (
            .O(N__17650),
            .I(N__17643));
    LocalMux I__2514 (
            .O(N__17647),
            .I(N__17637));
    InMux I__2513 (
            .O(N__17646),
            .I(N__17626));
    InMux I__2512 (
            .O(N__17643),
            .I(N__17626));
    InMux I__2511 (
            .O(N__17642),
            .I(N__17626));
    InMux I__2510 (
            .O(N__17641),
            .I(N__17626));
    InMux I__2509 (
            .O(N__17640),
            .I(N__17626));
    Odrv4 I__2508 (
            .O(N__17637),
            .I(RSMRST_PWRGD_curr_state_0));
    LocalMux I__2507 (
            .O(N__17626),
            .I(RSMRST_PWRGD_curr_state_0));
    InMux I__2506 (
            .O(N__17621),
            .I(N__17618));
    LocalMux I__2505 (
            .O(N__17618),
            .I(N_187));
    CascadeMux I__2504 (
            .O(N__17615),
            .I(G_11_cascade_));
    InMux I__2503 (
            .O(N__17612),
            .I(N__17609));
    LocalMux I__2502 (
            .O(N__17609),
            .I(\POWERLED.count_0_4 ));
    InMux I__2501 (
            .O(N__17606),
            .I(N__17603));
    LocalMux I__2500 (
            .O(N__17603),
            .I(\POWERLED.count_0_2 ));
    CascadeMux I__2499 (
            .O(N__17600),
            .I(\POWERLED.g0_i_o3_0_cascade_ ));
    InMux I__2498 (
            .O(N__17597),
            .I(N__17591));
    InMux I__2497 (
            .O(N__17596),
            .I(N__17591));
    LocalMux I__2496 (
            .O(N__17591),
            .I(\POWERLED.pwm_outZ0 ));
    InMux I__2495 (
            .O(N__17588),
            .I(N__17585));
    LocalMux I__2494 (
            .O(N__17585),
            .I(\POWERLED.g0_i_o3_0 ));
    IoInMux I__2493 (
            .O(N__17582),
            .I(N__17579));
    LocalMux I__2492 (
            .O(N__17579),
            .I(N__17576));
    Span4Mux_s3_v I__2491 (
            .O(N__17576),
            .I(N__17573));
    Span4Mux_v I__2490 (
            .O(N__17573),
            .I(N__17570));
    Span4Mux_v I__2489 (
            .O(N__17570),
            .I(N__17567));
    Odrv4 I__2488 (
            .O(N__17567),
            .I(pwrbtn_led));
    CascadeMux I__2487 (
            .O(N__17564),
            .I(\POWERLED.curr_state_3_0_cascade_ ));
    CascadeMux I__2486 (
            .O(N__17561),
            .I(\POWERLED.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__2485 (
            .O(N__17558),
            .I(\POWERLED.count_0_sqmuxa_i_cascade_ ));
    CascadeMux I__2484 (
            .O(N__17555),
            .I(\POWERLED.count_RNIZ0Z_0_cascade_ ));
    InMux I__2483 (
            .O(N__17552),
            .I(N__17546));
    InMux I__2482 (
            .O(N__17551),
            .I(N__17546));
    LocalMux I__2481 (
            .O(N__17546),
            .I(N__17543));
    Odrv12 I__2480 (
            .O(N__17543),
            .I(\PCH_PWRGD.count_rst_8 ));
    InMux I__2479 (
            .O(N__17540),
            .I(N__17536));
    InMux I__2478 (
            .O(N__17539),
            .I(N__17533));
    LocalMux I__2477 (
            .O(N__17536),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    LocalMux I__2476 (
            .O(N__17533),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    CascadeMux I__2475 (
            .O(N__17528),
            .I(N__17524));
    InMux I__2474 (
            .O(N__17527),
            .I(N__17519));
    InMux I__2473 (
            .O(N__17524),
            .I(N__17519));
    LocalMux I__2472 (
            .O(N__17519),
            .I(\PCH_PWRGD.count_rst_0 ));
    InMux I__2471 (
            .O(N__17516),
            .I(\PCH_PWRGD.un2_count_1_cry_13 ));
    InMux I__2470 (
            .O(N__17513),
            .I(N__17510));
    LocalMux I__2469 (
            .O(N__17510),
            .I(N__17507));
    Odrv4 I__2468 (
            .O(N__17507),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    InMux I__2467 (
            .O(N__17504),
            .I(\PCH_PWRGD.un2_count_1_cry_14 ));
    InMux I__2466 (
            .O(N__17501),
            .I(N__17495));
    InMux I__2465 (
            .O(N__17500),
            .I(N__17495));
    LocalMux I__2464 (
            .O(N__17495),
            .I(\PCH_PWRGD.count_rst ));
    CascadeMux I__2463 (
            .O(N__17492),
            .I(N__17489));
    InMux I__2462 (
            .O(N__17489),
            .I(N__17467));
    InMux I__2461 (
            .O(N__17488),
            .I(N__17467));
    InMux I__2460 (
            .O(N__17487),
            .I(N__17467));
    InMux I__2459 (
            .O(N__17486),
            .I(N__17467));
    InMux I__2458 (
            .O(N__17485),
            .I(N__17467));
    InMux I__2457 (
            .O(N__17484),
            .I(N__17460));
    InMux I__2456 (
            .O(N__17483),
            .I(N__17460));
    InMux I__2455 (
            .O(N__17482),
            .I(N__17460));
    InMux I__2454 (
            .O(N__17481),
            .I(N__17456));
    CascadeMux I__2453 (
            .O(N__17480),
            .I(N__17453));
    InMux I__2452 (
            .O(N__17479),
            .I(N__17450));
    CascadeMux I__2451 (
            .O(N__17478),
            .I(N__17443));
    LocalMux I__2450 (
            .O(N__17467),
            .I(N__17440));
    LocalMux I__2449 (
            .O(N__17460),
            .I(N__17437));
    InMux I__2448 (
            .O(N__17459),
            .I(N__17434));
    LocalMux I__2447 (
            .O(N__17456),
            .I(N__17431));
    InMux I__2446 (
            .O(N__17453),
            .I(N__17428));
    LocalMux I__2445 (
            .O(N__17450),
            .I(N__17425));
    InMux I__2444 (
            .O(N__17449),
            .I(N__17414));
    InMux I__2443 (
            .O(N__17448),
            .I(N__17414));
    InMux I__2442 (
            .O(N__17447),
            .I(N__17414));
    InMux I__2441 (
            .O(N__17446),
            .I(N__17414));
    InMux I__2440 (
            .O(N__17443),
            .I(N__17414));
    Span4Mux_h I__2439 (
            .O(N__17440),
            .I(N__17409));
    Span4Mux_s3_h I__2438 (
            .O(N__17437),
            .I(N__17409));
    LocalMux I__2437 (
            .O(N__17434),
            .I(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ));
    Odrv4 I__2436 (
            .O(N__17431),
            .I(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ));
    LocalMux I__2435 (
            .O(N__17428),
            .I(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ));
    Odrv4 I__2434 (
            .O(N__17425),
            .I(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ));
    LocalMux I__2433 (
            .O(N__17414),
            .I(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ));
    Odrv4 I__2432 (
            .O(N__17409),
            .I(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ));
    InMux I__2431 (
            .O(N__17396),
            .I(N__17370));
    InMux I__2430 (
            .O(N__17395),
            .I(N__17370));
    InMux I__2429 (
            .O(N__17394),
            .I(N__17370));
    InMux I__2428 (
            .O(N__17393),
            .I(N__17367));
    InMux I__2427 (
            .O(N__17392),
            .I(N__17364));
    InMux I__2426 (
            .O(N__17391),
            .I(N__17359));
    InMux I__2425 (
            .O(N__17390),
            .I(N__17359));
    InMux I__2424 (
            .O(N__17389),
            .I(N__17356));
    InMux I__2423 (
            .O(N__17388),
            .I(N__17347));
    InMux I__2422 (
            .O(N__17387),
            .I(N__17347));
    InMux I__2421 (
            .O(N__17386),
            .I(N__17347));
    InMux I__2420 (
            .O(N__17385),
            .I(N__17347));
    InMux I__2419 (
            .O(N__17384),
            .I(N__17336));
    InMux I__2418 (
            .O(N__17383),
            .I(N__17336));
    InMux I__2417 (
            .O(N__17382),
            .I(N__17336));
    InMux I__2416 (
            .O(N__17381),
            .I(N__17336));
    InMux I__2415 (
            .O(N__17380),
            .I(N__17336));
    InMux I__2414 (
            .O(N__17379),
            .I(N__17323));
    InMux I__2413 (
            .O(N__17378),
            .I(N__17323));
    InMux I__2412 (
            .O(N__17377),
            .I(N__17323));
    LocalMux I__2411 (
            .O(N__17370),
            .I(N__17320));
    LocalMux I__2410 (
            .O(N__17367),
            .I(N__17307));
    LocalMux I__2409 (
            .O(N__17364),
            .I(N__17307));
    LocalMux I__2408 (
            .O(N__17359),
            .I(N__17307));
    LocalMux I__2407 (
            .O(N__17356),
            .I(N__17307));
    LocalMux I__2406 (
            .O(N__17347),
            .I(N__17307));
    LocalMux I__2405 (
            .O(N__17336),
            .I(N__17307));
    InMux I__2404 (
            .O(N__17335),
            .I(N__17295));
    InMux I__2403 (
            .O(N__17334),
            .I(N__17295));
    InMux I__2402 (
            .O(N__17333),
            .I(N__17295));
    InMux I__2401 (
            .O(N__17332),
            .I(N__17295));
    InMux I__2400 (
            .O(N__17331),
            .I(N__17295));
    InMux I__2399 (
            .O(N__17330),
            .I(N__17292));
    LocalMux I__2398 (
            .O(N__17323),
            .I(N__17285));
    Span4Mux_h I__2397 (
            .O(N__17320),
            .I(N__17285));
    Span4Mux_s2_v I__2396 (
            .O(N__17307),
            .I(N__17285));
    InMux I__2395 (
            .O(N__17306),
            .I(N__17282));
    LocalMux I__2394 (
            .O(N__17295),
            .I(N__17279));
    LocalMux I__2393 (
            .O(N__17292),
            .I(\PCH_PWRGD.N_386 ));
    Odrv4 I__2392 (
            .O(N__17285),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__2391 (
            .O(N__17282),
            .I(\PCH_PWRGD.N_386 ));
    Odrv4 I__2390 (
            .O(N__17279),
            .I(\PCH_PWRGD.N_386 ));
    CascadeMux I__2389 (
            .O(N__17270),
            .I(N__17267));
    InMux I__2388 (
            .O(N__17267),
            .I(N__17260));
    InMux I__2387 (
            .O(N__17266),
            .I(N__17260));
    InMux I__2386 (
            .O(N__17265),
            .I(N__17257));
    LocalMux I__2385 (
            .O(N__17260),
            .I(N__17254));
    LocalMux I__2384 (
            .O(N__17257),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    Odrv4 I__2383 (
            .O(N__17254),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    InMux I__2382 (
            .O(N__17249),
            .I(N__17246));
    LocalMux I__2381 (
            .O(N__17246),
            .I(N__17242));
    InMux I__2380 (
            .O(N__17245),
            .I(N__17239));
    Odrv4 I__2379 (
            .O(N__17242),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    LocalMux I__2378 (
            .O(N__17239),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    InMux I__2377 (
            .O(N__17234),
            .I(N__17231));
    LocalMux I__2376 (
            .O(N__17231),
            .I(N__17228));
    Odrv4 I__2375 (
            .O(N__17228),
            .I(\PCH_PWRGD.count_rst_5 ));
    CascadeMux I__2374 (
            .O(N__17225),
            .I(\RSMRST_PWRGD.un4_count_9_cascade_ ));
    InMux I__2373 (
            .O(N__17222),
            .I(N__17218));
    InMux I__2372 (
            .O(N__17221),
            .I(N__17215));
    LocalMux I__2371 (
            .O(N__17218),
            .I(\RSMRST_PWRGD.N_1_i ));
    LocalMux I__2370 (
            .O(N__17215),
            .I(\RSMRST_PWRGD.N_1_i ));
    InMux I__2369 (
            .O(N__17210),
            .I(N__17207));
    LocalMux I__2368 (
            .O(N__17207),
            .I(\RSMRST_PWRGD.un4_count_8 ));
    InMux I__2367 (
            .O(N__17204),
            .I(N__17201));
    LocalMux I__2366 (
            .O(N__17201),
            .I(\RSMRST_PWRGD.un4_count_10 ));
    InMux I__2365 (
            .O(N__17198),
            .I(N__17195));
    LocalMux I__2364 (
            .O(N__17195),
            .I(\RSMRST_PWRGD.un4_count_11 ));
    InMux I__2363 (
            .O(N__17192),
            .I(N__17186));
    InMux I__2362 (
            .O(N__17191),
            .I(N__17186));
    LocalMux I__2361 (
            .O(N__17186),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    InMux I__2360 (
            .O(N__17183),
            .I(\PCH_PWRGD.un2_count_1_cry_4 ));
    InMux I__2359 (
            .O(N__17180),
            .I(\PCH_PWRGD.un2_count_1_cry_5 ));
    InMux I__2358 (
            .O(N__17177),
            .I(N__17170));
    InMux I__2357 (
            .O(N__17176),
            .I(N__17170));
    InMux I__2356 (
            .O(N__17175),
            .I(N__17167));
    LocalMux I__2355 (
            .O(N__17170),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    LocalMux I__2354 (
            .O(N__17167),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    CascadeMux I__2353 (
            .O(N__17162),
            .I(N__17158));
    InMux I__2352 (
            .O(N__17161),
            .I(N__17155));
    InMux I__2351 (
            .O(N__17158),
            .I(N__17152));
    LocalMux I__2350 (
            .O(N__17155),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    LocalMux I__2349 (
            .O(N__17152),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    InMux I__2348 (
            .O(N__17147),
            .I(\PCH_PWRGD.un2_count_1_cry_6 ));
    InMux I__2347 (
            .O(N__17144),
            .I(N__17139));
    CascadeMux I__2346 (
            .O(N__17143),
            .I(N__17136));
    CascadeMux I__2345 (
            .O(N__17142),
            .I(N__17133));
    LocalMux I__2344 (
            .O(N__17139),
            .I(N__17130));
    InMux I__2343 (
            .O(N__17136),
            .I(N__17125));
    InMux I__2342 (
            .O(N__17133),
            .I(N__17125));
    Span4Mux_h I__2341 (
            .O(N__17130),
            .I(N__17122));
    LocalMux I__2340 (
            .O(N__17125),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    Odrv4 I__2339 (
            .O(N__17122),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    InMux I__2338 (
            .O(N__17117),
            .I(N__17111));
    InMux I__2337 (
            .O(N__17116),
            .I(N__17111));
    LocalMux I__2336 (
            .O(N__17111),
            .I(N__17108));
    Span4Mux_s1_v I__2335 (
            .O(N__17108),
            .I(N__17105));
    Odrv4 I__2334 (
            .O(N__17105),
            .I(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__2333 (
            .O(N__17102),
            .I(\PCH_PWRGD.un2_count_1_cry_7 ));
    InMux I__2332 (
            .O(N__17099),
            .I(bfn_5_3_0_));
    InMux I__2331 (
            .O(N__17096),
            .I(\PCH_PWRGD.un2_count_1_cry_9 ));
    InMux I__2330 (
            .O(N__17093),
            .I(N__17089));
    InMux I__2329 (
            .O(N__17092),
            .I(N__17086));
    LocalMux I__2328 (
            .O(N__17089),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    LocalMux I__2327 (
            .O(N__17086),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    InMux I__2326 (
            .O(N__17081),
            .I(N__17075));
    InMux I__2325 (
            .O(N__17080),
            .I(N__17075));
    LocalMux I__2324 (
            .O(N__17075),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    InMux I__2323 (
            .O(N__17072),
            .I(\PCH_PWRGD.un2_count_1_cry_10 ));
    InMux I__2322 (
            .O(N__17069),
            .I(\PCH_PWRGD.un2_count_1_cry_11 ));
    InMux I__2321 (
            .O(N__17066),
            .I(N__17062));
    InMux I__2320 (
            .O(N__17065),
            .I(N__17059));
    LocalMux I__2319 (
            .O(N__17062),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    LocalMux I__2318 (
            .O(N__17059),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    InMux I__2317 (
            .O(N__17054),
            .I(N__17048));
    InMux I__2316 (
            .O(N__17053),
            .I(N__17048));
    LocalMux I__2315 (
            .O(N__17048),
            .I(\PCH_PWRGD.count_rst_1 ));
    InMux I__2314 (
            .O(N__17045),
            .I(\PCH_PWRGD.un2_count_1_cry_12 ));
    CascadeMux I__2313 (
            .O(N__17042),
            .I(\PCH_PWRGD.count_rst_7_cascade_ ));
    CascadeMux I__2312 (
            .O(N__17039),
            .I(\PCH_PWRGD.countZ0Z_7_cascade_ ));
    InMux I__2311 (
            .O(N__17036),
            .I(N__17033));
    LocalMux I__2310 (
            .O(N__17033),
            .I(\PCH_PWRGD.count_0_7 ));
    InMux I__2309 (
            .O(N__17030),
            .I(N__17027));
    LocalMux I__2308 (
            .O(N__17027),
            .I(N__17024));
    Odrv4 I__2307 (
            .O(N__17024),
            .I(\PCH_PWRGD.count_0_9 ));
    InMux I__2306 (
            .O(N__17021),
            .I(N__17017));
    InMux I__2305 (
            .O(N__17020),
            .I(N__17014));
    LocalMux I__2304 (
            .O(N__17017),
            .I(N__17010));
    LocalMux I__2303 (
            .O(N__17014),
            .I(N__17007));
    InMux I__2302 (
            .O(N__17013),
            .I(N__17004));
    Span4Mux_h I__2301 (
            .O(N__17010),
            .I(N__17001));
    Span4Mux_h I__2300 (
            .O(N__17007),
            .I(N__16998));
    LocalMux I__2299 (
            .O(N__17004),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    Odrv4 I__2298 (
            .O(N__17001),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    Odrv4 I__2297 (
            .O(N__16998),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    CascadeMux I__2296 (
            .O(N__16991),
            .I(N__16986));
    InMux I__2295 (
            .O(N__16990),
            .I(N__16983));
    InMux I__2294 (
            .O(N__16989),
            .I(N__16980));
    InMux I__2293 (
            .O(N__16986),
            .I(N__16977));
    LocalMux I__2292 (
            .O(N__16983),
            .I(N__16973));
    LocalMux I__2291 (
            .O(N__16980),
            .I(N__16970));
    LocalMux I__2290 (
            .O(N__16977),
            .I(N__16967));
    InMux I__2289 (
            .O(N__16976),
            .I(N__16964));
    Span4Mux_v I__2288 (
            .O(N__16973),
            .I(N__16961));
    Span4Mux_h I__2287 (
            .O(N__16970),
            .I(N__16958));
    Span4Mux_v I__2286 (
            .O(N__16967),
            .I(N__16955));
    LocalMux I__2285 (
            .O(N__16964),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    Odrv4 I__2284 (
            .O(N__16961),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    Odrv4 I__2283 (
            .O(N__16958),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    Odrv4 I__2282 (
            .O(N__16955),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    InMux I__2281 (
            .O(N__16946),
            .I(\PCH_PWRGD.un2_count_1_cry_1 ));
    InMux I__2280 (
            .O(N__16943),
            .I(N__16939));
    InMux I__2279 (
            .O(N__16942),
            .I(N__16936));
    LocalMux I__2278 (
            .O(N__16939),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    LocalMux I__2277 (
            .O(N__16936),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    InMux I__2276 (
            .O(N__16931),
            .I(N__16928));
    LocalMux I__2275 (
            .O(N__16928),
            .I(N__16924));
    InMux I__2274 (
            .O(N__16927),
            .I(N__16921));
    Odrv4 I__2273 (
            .O(N__16924),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    LocalMux I__2272 (
            .O(N__16921),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    InMux I__2271 (
            .O(N__16916),
            .I(\PCH_PWRGD.un2_count_1_cry_2 ));
    CascadeMux I__2270 (
            .O(N__16913),
            .I(N__16910));
    InMux I__2269 (
            .O(N__16910),
            .I(N__16905));
    InMux I__2268 (
            .O(N__16909),
            .I(N__16902));
    InMux I__2267 (
            .O(N__16908),
            .I(N__16899));
    LocalMux I__2266 (
            .O(N__16905),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__2265 (
            .O(N__16902),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__2264 (
            .O(N__16899),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    InMux I__2263 (
            .O(N__16892),
            .I(N__16886));
    InMux I__2262 (
            .O(N__16891),
            .I(N__16886));
    LocalMux I__2261 (
            .O(N__16886),
            .I(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__2260 (
            .O(N__16883),
            .I(\PCH_PWRGD.un2_count_1_cry_3 ));
    CascadeMux I__2259 (
            .O(N__16880),
            .I(N__16877));
    InMux I__2258 (
            .O(N__16877),
            .I(N__16873));
    InMux I__2257 (
            .O(N__16876),
            .I(N__16870));
    LocalMux I__2256 (
            .O(N__16873),
            .I(\PCH_PWRGD.un2_count_1_axb_5 ));
    LocalMux I__2255 (
            .O(N__16870),
            .I(\PCH_PWRGD.un2_count_1_axb_5 ));
    InMux I__2254 (
            .O(N__16865),
            .I(N__16862));
    LocalMux I__2253 (
            .O(N__16862),
            .I(N__16859));
    Odrv4 I__2252 (
            .O(N__16859),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__2251 (
            .O(N__16856),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__2250 (
            .O(N__16853),
            .I(N__16850));
    LocalMux I__2249 (
            .O(N__16850),
            .I(N__16847));
    Odrv4 I__2248 (
            .O(N__16847),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    InMux I__2247 (
            .O(N__16844),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__2246 (
            .O(N__16841),
            .I(N__16838));
    LocalMux I__2245 (
            .O(N__16838),
            .I(N__16835));
    Odrv4 I__2244 (
            .O(N__16835),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__2243 (
            .O(N__16832),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__2242 (
            .O(N__16829),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    InMux I__2241 (
            .O(N__16826),
            .I(N__16823));
    LocalMux I__2240 (
            .O(N__16823),
            .I(N__16819));
    CascadeMux I__2239 (
            .O(N__16822),
            .I(N__16816));
    Span4Mux_h I__2238 (
            .O(N__16819),
            .I(N__16810));
    InMux I__2237 (
            .O(N__16816),
            .I(N__16803));
    InMux I__2236 (
            .O(N__16815),
            .I(N__16803));
    InMux I__2235 (
            .O(N__16814),
            .I(N__16803));
    InMux I__2234 (
            .O(N__16813),
            .I(N__16800));
    Span4Mux_v I__2233 (
            .O(N__16810),
            .I(N__16795));
    LocalMux I__2232 (
            .O(N__16803),
            .I(N__16795));
    LocalMux I__2231 (
            .O(N__16800),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    Odrv4 I__2230 (
            .O(N__16795),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__2229 (
            .O(N__16790),
            .I(N__16786));
    CascadeMux I__2228 (
            .O(N__16789),
            .I(N__16782));
    InMux I__2227 (
            .O(N__16786),
            .I(N__16775));
    InMux I__2226 (
            .O(N__16785),
            .I(N__16775));
    InMux I__2225 (
            .O(N__16782),
            .I(N__16775));
    LocalMux I__2224 (
            .O(N__16775),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    CascadeMux I__2223 (
            .O(N__16772),
            .I(\PCH_PWRGD.un2_count_1_axb_5_cascade_ ));
    InMux I__2222 (
            .O(N__16769),
            .I(N__16763));
    InMux I__2221 (
            .O(N__16768),
            .I(N__16763));
    LocalMux I__2220 (
            .O(N__16763),
            .I(\PCH_PWRGD.count_0_5 ));
    InMux I__2219 (
            .O(N__16760),
            .I(N__16757));
    LocalMux I__2218 (
            .O(N__16757),
            .I(N__16754));
    Span4Mux_v I__2217 (
            .O(N__16754),
            .I(N__16751));
    Odrv4 I__2216 (
            .O(N__16751),
            .I(\PCH_PWRGD.un12_clk_100khz_6 ));
    InMux I__2215 (
            .O(N__16748),
            .I(N__16742));
    InMux I__2214 (
            .O(N__16747),
            .I(N__16742));
    LocalMux I__2213 (
            .O(N__16742),
            .I(\PCH_PWRGD.count_rst_9 ));
    InMux I__2212 (
            .O(N__16739),
            .I(N__16736));
    LocalMux I__2211 (
            .O(N__16736),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    InMux I__2210 (
            .O(N__16733),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    CascadeMux I__2209 (
            .O(N__16730),
            .I(N__16726));
    InMux I__2208 (
            .O(N__16729),
            .I(N__16720));
    InMux I__2207 (
            .O(N__16726),
            .I(N__16720));
    InMux I__2206 (
            .O(N__16725),
            .I(N__16717));
    LocalMux I__2205 (
            .O(N__16720),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    LocalMux I__2204 (
            .O(N__16717),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__2203 (
            .O(N__16712),
            .I(N__16709));
    InMux I__2202 (
            .O(N__16709),
            .I(N__16706));
    LocalMux I__2201 (
            .O(N__16706),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__2200 (
            .O(N__16703),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__2199 (
            .O(N__16700),
            .I(N__16697));
    LocalMux I__2198 (
            .O(N__16697),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    CascadeMux I__2197 (
            .O(N__16694),
            .I(N__16690));
    CascadeMux I__2196 (
            .O(N__16693),
            .I(N__16686));
    InMux I__2195 (
            .O(N__16690),
            .I(N__16679));
    InMux I__2194 (
            .O(N__16689),
            .I(N__16679));
    InMux I__2193 (
            .O(N__16686),
            .I(N__16679));
    LocalMux I__2192 (
            .O(N__16679),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    InMux I__2191 (
            .O(N__16676),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    CascadeMux I__2190 (
            .O(N__16673),
            .I(N__16670));
    InMux I__2189 (
            .O(N__16670),
            .I(N__16667));
    LocalMux I__2188 (
            .O(N__16667),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__2187 (
            .O(N__16664),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__2186 (
            .O(N__16661),
            .I(\POWERLED.mult1_un61_sum_s_8_cascade_ ));
    CascadeMux I__2185 (
            .O(N__16658),
            .I(N__16655));
    InMux I__2184 (
            .O(N__16655),
            .I(N__16652));
    LocalMux I__2183 (
            .O(N__16652),
            .I(N__16649));
    Odrv4 I__2182 (
            .O(N__16649),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__2181 (
            .O(N__16646),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    CascadeMux I__2180 (
            .O(N__16643),
            .I(N__16640));
    InMux I__2179 (
            .O(N__16640),
            .I(N__16637));
    LocalMux I__2178 (
            .O(N__16637),
            .I(N__16634));
    Odrv12 I__2177 (
            .O(N__16634),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__2176 (
            .O(N__16631),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__2175 (
            .O(N__16628),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__2174 (
            .O(N__16625),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__2173 (
            .O(N__16622),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__2172 (
            .O(N__16619),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__2171 (
            .O(N__16616),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    CascadeMux I__2170 (
            .O(N__16613),
            .I(\POWERLED.mult1_un54_sum_s_8_cascade_ ));
    InMux I__2169 (
            .O(N__16610),
            .I(N__16607));
    LocalMux I__2168 (
            .O(N__16607),
            .I(N__16604));
    Odrv4 I__2167 (
            .O(N__16604),
            .I(\POWERLED.mult1_un54_sum_i ));
    InMux I__2166 (
            .O(N__16601),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__2165 (
            .O(N__16598),
            .I(N__16595));
    InMux I__2164 (
            .O(N__16595),
            .I(N__16592));
    LocalMux I__2163 (
            .O(N__16592),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__2162 (
            .O(N__16589),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    CascadeMux I__2161 (
            .O(N__16586),
            .I(\POWERLED.un2_count_clk_17_0_a2_5_cascade_ ));
    CascadeMux I__2160 (
            .O(N__16583),
            .I(\POWERLED.un1_dutycycle_53_46_0_cascade_ ));
    InMux I__2159 (
            .O(N__16580),
            .I(N__16577));
    LocalMux I__2158 (
            .O(N__16577),
            .I(N__16574));
    Odrv4 I__2157 (
            .O(N__16574),
            .I(\POWERLED.mult1_un47_sum_i ));
    InMux I__2156 (
            .O(N__16571),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    CascadeMux I__2155 (
            .O(N__16568),
            .I(N__16565));
    InMux I__2154 (
            .O(N__16565),
            .I(N__16562));
    LocalMux I__2153 (
            .O(N__16562),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__2152 (
            .O(N__16559),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    InMux I__2151 (
            .O(N__16556),
            .I(N__16553));
    LocalMux I__2150 (
            .O(N__16553),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    InMux I__2149 (
            .O(N__16550),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__2148 (
            .O(N__16547),
            .I(N__16544));
    LocalMux I__2147 (
            .O(N__16544),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    InMux I__2146 (
            .O(N__16541),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    InMux I__2145 (
            .O(N__16538),
            .I(N__16535));
    LocalMux I__2144 (
            .O(N__16535),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__2143 (
            .O(N__16532),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__2142 (
            .O(N__16529),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    InMux I__2141 (
            .O(N__16526),
            .I(N__16523));
    LocalMux I__2140 (
            .O(N__16523),
            .I(N__16519));
    CascadeMux I__2139 (
            .O(N__16522),
            .I(N__16516));
    Span4Mux_v I__2138 (
            .O(N__16519),
            .I(N__16510));
    InMux I__2137 (
            .O(N__16516),
            .I(N__16503));
    InMux I__2136 (
            .O(N__16515),
            .I(N__16503));
    InMux I__2135 (
            .O(N__16514),
            .I(N__16503));
    InMux I__2134 (
            .O(N__16513),
            .I(N__16500));
    Odrv4 I__2133 (
            .O(N__16510),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__2132 (
            .O(N__16503),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__2131 (
            .O(N__16500),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    CascadeMux I__2130 (
            .O(N__16493),
            .I(N__16490));
    InMux I__2129 (
            .O(N__16490),
            .I(N__16487));
    LocalMux I__2128 (
            .O(N__16487),
            .I(\POWERLED.mult1_un152_sum_i ));
    CascadeMux I__2127 (
            .O(N__16484),
            .I(N__16480));
    InMux I__2126 (
            .O(N__16483),
            .I(N__16472));
    InMux I__2125 (
            .O(N__16480),
            .I(N__16472));
    InMux I__2124 (
            .O(N__16479),
            .I(N__16472));
    LocalMux I__2123 (
            .O(N__16472),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    CascadeMux I__2122 (
            .O(N__16469),
            .I(N__16466));
    InMux I__2121 (
            .O(N__16466),
            .I(N__16463));
    LocalMux I__2120 (
            .O(N__16463),
            .I(N__16460));
    Span4Mux_v I__2119 (
            .O(N__16460),
            .I(N__16457));
    Span4Mux_v I__2118 (
            .O(N__16457),
            .I(N__16454));
    Odrv4 I__2117 (
            .O(N__16454),
            .I(\POWERLED.un85_clk_100khz_2 ));
    CascadeMux I__2116 (
            .O(N__16451),
            .I(N__16447));
    CascadeMux I__2115 (
            .O(N__16450),
            .I(N__16443));
    InMux I__2114 (
            .O(N__16447),
            .I(N__16436));
    InMux I__2113 (
            .O(N__16446),
            .I(N__16436));
    InMux I__2112 (
            .O(N__16443),
            .I(N__16436));
    LocalMux I__2111 (
            .O(N__16436),
            .I(G_2121));
    InMux I__2110 (
            .O(N__16433),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    CascadeMux I__2109 (
            .O(N__16430),
            .I(N__16427));
    InMux I__2108 (
            .O(N__16427),
            .I(N__16424));
    LocalMux I__2107 (
            .O(N__16424),
            .I(N__16421));
    Odrv12 I__2106 (
            .O(N__16421),
            .I(\POWERLED.un85_clk_100khz_0 ));
    InMux I__2105 (
            .O(N__16418),
            .I(N__16415));
    LocalMux I__2104 (
            .O(N__16415),
            .I(\POWERLED.mult1_un159_sum_i ));
    CascadeMux I__2103 (
            .O(N__16412),
            .I(N__16409));
    InMux I__2102 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__2101 (
            .O(N__16406),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    InMux I__2100 (
            .O(N__16403),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    CascadeMux I__2099 (
            .O(N__16400),
            .I(N__16397));
    InMux I__2098 (
            .O(N__16397),
            .I(N__16394));
    LocalMux I__2097 (
            .O(N__16394),
            .I(N__16391));
    Odrv4 I__2096 (
            .O(N__16391),
            .I(\COUNTER.un4_counter_3_and ));
    CascadeMux I__2095 (
            .O(N__16388),
            .I(N__16385));
    InMux I__2094 (
            .O(N__16385),
            .I(N__16382));
    LocalMux I__2093 (
            .O(N__16382),
            .I(N__16379));
    Odrv4 I__2092 (
            .O(N__16379),
            .I(\COUNTER.un4_counter_4_and ));
    CascadeMux I__2091 (
            .O(N__16376),
            .I(N__16373));
    InMux I__2090 (
            .O(N__16373),
            .I(N__16370));
    LocalMux I__2089 (
            .O(N__16370),
            .I(N__16367));
    Odrv4 I__2088 (
            .O(N__16367),
            .I(\COUNTER.un4_counter_5_and ));
    InMux I__2087 (
            .O(N__16364),
            .I(N__16361));
    LocalMux I__2086 (
            .O(N__16361),
            .I(N__16358));
    Odrv4 I__2085 (
            .O(N__16358),
            .I(\COUNTER.un4_counter_6_and ));
    CascadeMux I__2084 (
            .O(N__16355),
            .I(N__16352));
    InMux I__2083 (
            .O(N__16352),
            .I(N__16349));
    LocalMux I__2082 (
            .O(N__16349),
            .I(N__16346));
    Span4Mux_h I__2081 (
            .O(N__16346),
            .I(N__16343));
    Odrv4 I__2080 (
            .O(N__16343),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__2079 (
            .O(N__16340),
            .I(bfn_4_8_0_));
    IoInMux I__2078 (
            .O(N__16337),
            .I(N__16334));
    LocalMux I__2077 (
            .O(N__16334),
            .I(N__16330));
    IoInMux I__2076 (
            .O(N__16333),
            .I(N__16327));
    Span4Mux_s2_h I__2075 (
            .O(N__16330),
            .I(N__16324));
    LocalMux I__2074 (
            .O(N__16327),
            .I(N__16321));
    Span4Mux_v I__2073 (
            .O(N__16324),
            .I(N__16318));
    Span4Mux_s3_h I__2072 (
            .O(N__16321),
            .I(N__16315));
    Odrv4 I__2071 (
            .O(N__16318),
            .I(v5s_enn));
    Odrv4 I__2070 (
            .O(N__16315),
            .I(v5s_enn));
    CascadeMux I__2069 (
            .O(N__16310),
            .I(N_187_cascade_));
    IoInMux I__2068 (
            .O(N__16307),
            .I(N__16303));
    IoInMux I__2067 (
            .O(N__16306),
            .I(N__16300));
    LocalMux I__2066 (
            .O(N__16303),
            .I(N__16297));
    LocalMux I__2065 (
            .O(N__16300),
            .I(N__16293));
    Span4Mux_s3_h I__2064 (
            .O(N__16297),
            .I(N__16290));
    InMux I__2063 (
            .O(N__16296),
            .I(N__16287));
    IoSpan4Mux I__2062 (
            .O(N__16293),
            .I(N__16284));
    Sp12to4 I__2061 (
            .O(N__16290),
            .I(N__16279));
    LocalMux I__2060 (
            .O(N__16287),
            .I(N__16279));
    IoSpan4Mux I__2059 (
            .O(N__16284),
            .I(N__16276));
    Span12Mux_v I__2058 (
            .O(N__16279),
            .I(N__16273));
    IoSpan4Mux I__2057 (
            .O(N__16276),
            .I(N__16270));
    Odrv12 I__2056 (
            .O(N__16273),
            .I(v33a_ok));
    Odrv4 I__2055 (
            .O(N__16270),
            .I(v33a_ok));
    InMux I__2054 (
            .O(N__16265),
            .I(N__16262));
    LocalMux I__2053 (
            .O(N__16262),
            .I(N__16259));
    Odrv12 I__2052 (
            .O(N__16259),
            .I(v5a_ok));
    InMux I__2051 (
            .O(N__16256),
            .I(N__16252));
    CascadeMux I__2050 (
            .O(N__16255),
            .I(N__16249));
    LocalMux I__2049 (
            .O(N__16252),
            .I(N__16246));
    InMux I__2048 (
            .O(N__16249),
            .I(N__16243));
    Span4Mux_h I__2047 (
            .O(N__16246),
            .I(N__16240));
    LocalMux I__2046 (
            .O(N__16243),
            .I(N__16237));
    Span4Mux_v I__2045 (
            .O(N__16240),
            .I(N__16234));
    Span12Mux_s8_h I__2044 (
            .O(N__16237),
            .I(N__16231));
    Span4Mux_h I__2043 (
            .O(N__16234),
            .I(N__16228));
    Odrv12 I__2042 (
            .O(N__16231),
            .I(slp_susn));
    Odrv4 I__2041 (
            .O(N__16228),
            .I(slp_susn));
    IoInMux I__2040 (
            .O(N__16223),
            .I(N__16220));
    LocalMux I__2039 (
            .O(N__16220),
            .I(N__16216));
    InMux I__2038 (
            .O(N__16219),
            .I(N__16213));
    Span4Mux_s2_h I__2037 (
            .O(N__16216),
            .I(N__16210));
    LocalMux I__2036 (
            .O(N__16213),
            .I(N__16207));
    Sp12to4 I__2035 (
            .O(N__16210),
            .I(N__16204));
    Span4Mux_v I__2034 (
            .O(N__16207),
            .I(N__16201));
    Span12Mux_s11_v I__2033 (
            .O(N__16204),
            .I(N__16198));
    Span4Mux_v I__2032 (
            .O(N__16201),
            .I(N__16195));
    Odrv12 I__2031 (
            .O(N__16198),
            .I(v1p8a_ok));
    Odrv4 I__2030 (
            .O(N__16195),
            .I(v1p8a_ok));
    CascadeMux I__2029 (
            .O(N__16190),
            .I(rsmrst_pwrgd_signal_cascade_));
    InMux I__2028 (
            .O(N__16187),
            .I(N__16177));
    InMux I__2027 (
            .O(N__16186),
            .I(N__16177));
    InMux I__2026 (
            .O(N__16185),
            .I(N__16168));
    InMux I__2025 (
            .O(N__16184),
            .I(N__16168));
    InMux I__2024 (
            .O(N__16183),
            .I(N__16168));
    InMux I__2023 (
            .O(N__16182),
            .I(N__16168));
    LocalMux I__2022 (
            .O(N__16177),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__2021 (
            .O(N__16168),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__2020 (
            .O(N__16163),
            .I(N__16160));
    InMux I__2019 (
            .O(N__16160),
            .I(N__16157));
    LocalMux I__2018 (
            .O(N__16157),
            .I(N__16154));
    Span4Mux_v I__2017 (
            .O(N__16154),
            .I(N__16151));
    Odrv4 I__2016 (
            .O(N__16151),
            .I(\COUNTER.un4_counter_0_and ));
    CascadeMux I__2015 (
            .O(N__16148),
            .I(N__16145));
    InMux I__2014 (
            .O(N__16145),
            .I(N__16142));
    LocalMux I__2013 (
            .O(N__16142),
            .I(N__16139));
    Span4Mux_h I__2012 (
            .O(N__16139),
            .I(N__16136));
    Odrv4 I__2011 (
            .O(N__16136),
            .I(\COUNTER.un4_counter_1_and ));
    CascadeMux I__2010 (
            .O(N__16133),
            .I(N__16130));
    InMux I__2009 (
            .O(N__16130),
            .I(N__16127));
    LocalMux I__2008 (
            .O(N__16127),
            .I(N__16124));
    Odrv4 I__2007 (
            .O(N__16124),
            .I(\COUNTER.un4_counter_2_and ));
    InMux I__2006 (
            .O(N__16121),
            .I(N__16113));
    InMux I__2005 (
            .O(N__16120),
            .I(N__16110));
    InMux I__2004 (
            .O(N__16119),
            .I(N__16107));
    InMux I__2003 (
            .O(N__16118),
            .I(N__16104));
    InMux I__2002 (
            .O(N__16117),
            .I(N__16099));
    InMux I__2001 (
            .O(N__16116),
            .I(N__16099));
    LocalMux I__2000 (
            .O(N__16113),
            .I(N__16092));
    LocalMux I__1999 (
            .O(N__16110),
            .I(N__16092));
    LocalMux I__1998 (
            .O(N__16107),
            .I(N__16092));
    LocalMux I__1997 (
            .O(N__16104),
            .I(N__16089));
    LocalMux I__1996 (
            .O(N__16099),
            .I(N__16084));
    Span4Mux_v I__1995 (
            .O(N__16092),
            .I(N__16084));
    Odrv12 I__1994 (
            .O(N__16089),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__1993 (
            .O(N__16084),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    InMux I__1992 (
            .O(N__16079),
            .I(N__16076));
    LocalMux I__1991 (
            .O(N__16076),
            .I(N__16072));
    InMux I__1990 (
            .O(N__16075),
            .I(N__16069));
    Span4Mux_h I__1989 (
            .O(N__16072),
            .I(N__16062));
    LocalMux I__1988 (
            .O(N__16069),
            .I(N__16062));
    InMux I__1987 (
            .O(N__16068),
            .I(N__16057));
    InMux I__1986 (
            .O(N__16067),
            .I(N__16057));
    Span4Mux_s3_h I__1985 (
            .O(N__16062),
            .I(N__16054));
    LocalMux I__1984 (
            .O(N__16057),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__1983 (
            .O(N__16054),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__1982 (
            .O(N__16049),
            .I(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2_cascade_ ));
    InMux I__1981 (
            .O(N__16046),
            .I(N__16043));
    LocalMux I__1980 (
            .O(N__16043),
            .I(N__16040));
    Odrv4 I__1979 (
            .O(N__16040),
            .I(\PCH_PWRGD.curr_state_7_1 ));
    CascadeMux I__1978 (
            .O(N__16037),
            .I(\PCH_PWRGD.countZ0Z_15_cascade_ ));
    InMux I__1977 (
            .O(N__16034),
            .I(N__16031));
    LocalMux I__1976 (
            .O(N__16031),
            .I(\PCH_PWRGD.un12_clk_100khz_8 ));
    InMux I__1975 (
            .O(N__16028),
            .I(N__16025));
    LocalMux I__1974 (
            .O(N__16025),
            .I(\PCH_PWRGD.count_0_14 ));
    InMux I__1973 (
            .O(N__16022),
            .I(N__16019));
    LocalMux I__1972 (
            .O(N__16019),
            .I(\PCH_PWRGD.count_0_13 ));
    InMux I__1971 (
            .O(N__16016),
            .I(N__16013));
    LocalMux I__1970 (
            .O(N__16013),
            .I(\PCH_PWRGD.count_0_15 ));
    InMux I__1969 (
            .O(N__16010),
            .I(N__16007));
    LocalMux I__1968 (
            .O(N__16007),
            .I(N__16004));
    Span4Mux_s1_v I__1967 (
            .O(N__16004),
            .I(N__16001));
    Odrv4 I__1966 (
            .O(N__16001),
            .I(\PCH_PWRGD.count_0_0 ));
    CascadeMux I__1965 (
            .O(N__15998),
            .I(\PCH_PWRGD.count_rst_3_cascade_ ));
    CascadeMux I__1964 (
            .O(N__15995),
            .I(\PCH_PWRGD.un2_count_1_axb_11_cascade_ ));
    InMux I__1963 (
            .O(N__15992),
            .I(N__15989));
    LocalMux I__1962 (
            .O(N__15989),
            .I(\PCH_PWRGD.count_rst_3 ));
    CascadeMux I__1961 (
            .O(N__15986),
            .I(N__15983));
    InMux I__1960 (
            .O(N__15983),
            .I(N__15977));
    InMux I__1959 (
            .O(N__15982),
            .I(N__15977));
    LocalMux I__1958 (
            .O(N__15977),
            .I(\PCH_PWRGD.count_0_11 ));
    InMux I__1957 (
            .O(N__15974),
            .I(N__15971));
    LocalMux I__1956 (
            .O(N__15971),
            .I(\PCH_PWRGD.un12_clk_100khz_7 ));
    CascadeMux I__1955 (
            .O(N__15968),
            .I(\PCH_PWRGD.un12_clk_100khz_4_cascade_ ));
    InMux I__1954 (
            .O(N__15965),
            .I(N__15962));
    LocalMux I__1953 (
            .O(N__15962),
            .I(N__15959));
    Odrv4 I__1952 (
            .O(N__15959),
            .I(\PCH_PWRGD.un12_clk_100khz_5 ));
    CascadeMux I__1951 (
            .O(N__15956),
            .I(\PCH_PWRGD.un12_clk_100khz_13_cascade_ ));
    InMux I__1950 (
            .O(N__15953),
            .I(N__15947));
    InMux I__1949 (
            .O(N__15952),
            .I(N__15947));
    LocalMux I__1948 (
            .O(N__15947),
            .I(N__15944));
    Odrv4 I__1947 (
            .O(N__15944),
            .I(\PCH_PWRGD.N_1_i ));
    CascadeMux I__1946 (
            .O(N__15941),
            .I(\PCH_PWRGD.N_1_i_cascade_ ));
    InMux I__1945 (
            .O(N__15938),
            .I(N__15935));
    LocalMux I__1944 (
            .O(N__15935),
            .I(N__15931));
    InMux I__1943 (
            .O(N__15934),
            .I(N__15928));
    Odrv12 I__1942 (
            .O(N__15931),
            .I(\PCH_PWRGD.count_0_8 ));
    LocalMux I__1941 (
            .O(N__15928),
            .I(\PCH_PWRGD.count_0_8 ));
    CascadeMux I__1940 (
            .O(N__15923),
            .I(\PCH_PWRGD.countZ0Z_9_cascade_ ));
    InMux I__1939 (
            .O(N__15920),
            .I(N__15917));
    LocalMux I__1938 (
            .O(N__15917),
            .I(N__15914));
    Odrv4 I__1937 (
            .O(N__15914),
            .I(\PCH_PWRGD.count_rst_6 ));
    CascadeMux I__1936 (
            .O(N__15911),
            .I(N__15907));
    InMux I__1935 (
            .O(N__15910),
            .I(N__15902));
    InMux I__1934 (
            .O(N__15907),
            .I(N__15902));
    LocalMux I__1933 (
            .O(N__15902),
            .I(N__15899));
    Span4Mux_s1_v I__1932 (
            .O(N__15899),
            .I(N__15895));
    InMux I__1931 (
            .O(N__15898),
            .I(N__15892));
    Odrv4 I__1930 (
            .O(N__15895),
            .I(\PCH_PWRGD.curr_state_RNI3DJUZ0Z_0 ));
    LocalMux I__1929 (
            .O(N__15892),
            .I(\PCH_PWRGD.curr_state_RNI3DJUZ0Z_0 ));
    InMux I__1928 (
            .O(N__15887),
            .I(N__15884));
    LocalMux I__1927 (
            .O(N__15884),
            .I(\PCH_PWRGD.curr_state_0_0 ));
    InMux I__1926 (
            .O(N__15881),
            .I(N__15878));
    LocalMux I__1925 (
            .O(N__15878),
            .I(\PCH_PWRGD.count_rst_11 ));
    CascadeMux I__1924 (
            .O(N__15875),
            .I(\PCH_PWRGD.count_rst_11_cascade_ ));
    CascadeMux I__1923 (
            .O(N__15872),
            .I(\PCH_PWRGD.un2_count_1_axb_3_cascade_ ));
    InMux I__1922 (
            .O(N__15869),
            .I(N__15863));
    InMux I__1921 (
            .O(N__15868),
            .I(N__15863));
    LocalMux I__1920 (
            .O(N__15863),
            .I(\PCH_PWRGD.count_0_3 ));
    CascadeMux I__1919 (
            .O(N__15860),
            .I(\PCH_PWRGD.count_rst_10_cascade_ ));
    CascadeMux I__1918 (
            .O(N__15857),
            .I(\PCH_PWRGD.countZ0Z_4_cascade_ ));
    InMux I__1917 (
            .O(N__15854),
            .I(N__15851));
    LocalMux I__1916 (
            .O(N__15851),
            .I(\PCH_PWRGD.count_0_4 ));
    InMux I__1915 (
            .O(N__15848),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    CascadeMux I__1914 (
            .O(N__15845),
            .I(N__15841));
    CascadeMux I__1913 (
            .O(N__15844),
            .I(N__15837));
    InMux I__1912 (
            .O(N__15841),
            .I(N__15830));
    InMux I__1911 (
            .O(N__15840),
            .I(N__15830));
    InMux I__1910 (
            .O(N__15837),
            .I(N__15830));
    LocalMux I__1909 (
            .O(N__15830),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__1908 (
            .O(N__15827),
            .I(N__15824));
    LocalMux I__1907 (
            .O(N__15824),
            .I(\POWERLED.mult1_un103_sum_i ));
    CascadeMux I__1906 (
            .O(N__15821),
            .I(N__15817));
    CascadeMux I__1905 (
            .O(N__15820),
            .I(N__15813));
    InMux I__1904 (
            .O(N__15817),
            .I(N__15806));
    InMux I__1903 (
            .O(N__15816),
            .I(N__15806));
    InMux I__1902 (
            .O(N__15813),
            .I(N__15806));
    LocalMux I__1901 (
            .O(N__15806),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    InMux I__1900 (
            .O(N__15803),
            .I(N__15800));
    LocalMux I__1899 (
            .O(N__15800),
            .I(\POWERLED.mult1_un96_sum_i ));
    CascadeMux I__1898 (
            .O(N__15797),
            .I(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__1897 (
            .O(N__15794),
            .I(\PCH_PWRGD.m4_0_0_cascade_ ));
    CascadeMux I__1896 (
            .O(N__15791),
            .I(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ));
    InMux I__1895 (
            .O(N__15788),
            .I(N__15785));
    LocalMux I__1894 (
            .O(N__15785),
            .I(\PCH_PWRGD.curr_state_0_1 ));
    InMux I__1893 (
            .O(N__15782),
            .I(N__15779));
    LocalMux I__1892 (
            .O(N__15779),
            .I(N__15776));
    Odrv12 I__1891 (
            .O(N__15776),
            .I(\POWERLED.un85_clk_100khz_14 ));
    InMux I__1890 (
            .O(N__15773),
            .I(N__15770));
    LocalMux I__1889 (
            .O(N__15770),
            .I(N__15767));
    Span4Mux_s3_v I__1888 (
            .O(N__15767),
            .I(N__15764));
    Odrv4 I__1887 (
            .O(N__15764),
            .I(vpp_ok));
    IoInMux I__1886 (
            .O(N__15761),
            .I(N__15758));
    LocalMux I__1885 (
            .O(N__15758),
            .I(N__15755));
    Span4Mux_s2_v I__1884 (
            .O(N__15755),
            .I(N__15752));
    Odrv4 I__1883 (
            .O(N__15752),
            .I(vddq_en));
    InMux I__1882 (
            .O(N__15749),
            .I(N__15746));
    LocalMux I__1881 (
            .O(N__15746),
            .I(N__15743));
    Odrv4 I__1880 (
            .O(N__15743),
            .I(\POWERLED.mult1_un89_sum_i ));
    CascadeMux I__1879 (
            .O(N__15740),
            .I(N__15737));
    InMux I__1878 (
            .O(N__15737),
            .I(N__15734));
    LocalMux I__1877 (
            .O(N__15734),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__1876 (
            .O(N__15731),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    InMux I__1875 (
            .O(N__15728),
            .I(N__15725));
    LocalMux I__1874 (
            .O(N__15725),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    InMux I__1873 (
            .O(N__15722),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    InMux I__1872 (
            .O(N__15719),
            .I(N__15716));
    LocalMux I__1871 (
            .O(N__15716),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__1870 (
            .O(N__15713),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    InMux I__1869 (
            .O(N__15710),
            .I(N__15707));
    LocalMux I__1868 (
            .O(N__15707),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    InMux I__1867 (
            .O(N__15704),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    InMux I__1866 (
            .O(N__15701),
            .I(N__15698));
    LocalMux I__1865 (
            .O(N__15698),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__1864 (
            .O(N__15695),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    CascadeMux I__1863 (
            .O(N__15692),
            .I(N__15689));
    InMux I__1862 (
            .O(N__15689),
            .I(N__15686));
    LocalMux I__1861 (
            .O(N__15686),
            .I(N__15683));
    Span4Mux_v I__1860 (
            .O(N__15683),
            .I(N__15680));
    Odrv4 I__1859 (
            .O(N__15680),
            .I(\POWERLED.un85_clk_100khz_8 ));
    InMux I__1858 (
            .O(N__15677),
            .I(N__15674));
    LocalMux I__1857 (
            .O(N__15674),
            .I(\POWERLED.mult1_un117_sum_i ));
    CascadeMux I__1856 (
            .O(N__15671),
            .I(N__15666));
    CascadeMux I__1855 (
            .O(N__15670),
            .I(N__15663));
    InMux I__1854 (
            .O(N__15669),
            .I(N__15659));
    InMux I__1853 (
            .O(N__15666),
            .I(N__15656));
    InMux I__1852 (
            .O(N__15663),
            .I(N__15653));
    InMux I__1851 (
            .O(N__15662),
            .I(N__15650));
    LocalMux I__1850 (
            .O(N__15659),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1849 (
            .O(N__15656),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1848 (
            .O(N__15653),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1847 (
            .O(N__15650),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    CascadeMux I__1846 (
            .O(N__15641),
            .I(N__15638));
    InMux I__1845 (
            .O(N__15638),
            .I(N__15635));
    LocalMux I__1844 (
            .O(N__15635),
            .I(N__15632));
    Span4Mux_v I__1843 (
            .O(N__15632),
            .I(N__15629));
    Odrv4 I__1842 (
            .O(N__15629),
            .I(\POWERLED.un85_clk_100khz_7 ));
    CascadeMux I__1841 (
            .O(N__15626),
            .I(N__15623));
    InMux I__1840 (
            .O(N__15623),
            .I(N__15620));
    LocalMux I__1839 (
            .O(N__15620),
            .I(N__15617));
    Odrv4 I__1838 (
            .O(N__15617),
            .I(\POWERLED.un85_clk_100khz_12 ));
    InMux I__1837 (
            .O(N__15614),
            .I(N__15611));
    LocalMux I__1836 (
            .O(N__15611),
            .I(N__15608));
    Span4Mux_s2_h I__1835 (
            .O(N__15608),
            .I(N__15605));
    Odrv4 I__1834 (
            .O(N__15605),
            .I(\POWERLED.mult1_un61_sum_i_8 ));
    InMux I__1833 (
            .O(N__15602),
            .I(N__15599));
    LocalMux I__1832 (
            .O(N__15599),
            .I(\POWERLED.mult1_un110_sum_i ));
    InMux I__1831 (
            .O(N__15596),
            .I(N__15591));
    CascadeMux I__1830 (
            .O(N__15595),
            .I(N__15587));
    CascadeMux I__1829 (
            .O(N__15594),
            .I(N__15584));
    LocalMux I__1828 (
            .O(N__15591),
            .I(N__15580));
    InMux I__1827 (
            .O(N__15590),
            .I(N__15577));
    InMux I__1826 (
            .O(N__15587),
            .I(N__15574));
    InMux I__1825 (
            .O(N__15584),
            .I(N__15571));
    InMux I__1824 (
            .O(N__15583),
            .I(N__15568));
    Odrv4 I__1823 (
            .O(N__15580),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1822 (
            .O(N__15577),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1821 (
            .O(N__15574),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1820 (
            .O(N__15571),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1819 (
            .O(N__15568),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    CascadeMux I__1818 (
            .O(N__15557),
            .I(N__15552));
    CascadeMux I__1817 (
            .O(N__15556),
            .I(N__15549));
    CascadeMux I__1816 (
            .O(N__15555),
            .I(N__15546));
    InMux I__1815 (
            .O(N__15552),
            .I(N__15543));
    InMux I__1814 (
            .O(N__15549),
            .I(N__15538));
    InMux I__1813 (
            .O(N__15546),
            .I(N__15538));
    LocalMux I__1812 (
            .O(N__15543),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    LocalMux I__1811 (
            .O(N__15538),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    InMux I__1810 (
            .O(N__15533),
            .I(N__15530));
    LocalMux I__1809 (
            .O(N__15530),
            .I(N__15524));
    CascadeMux I__1808 (
            .O(N__15529),
            .I(N__15521));
    CascadeMux I__1807 (
            .O(N__15528),
            .I(N__15518));
    InMux I__1806 (
            .O(N__15527),
            .I(N__15515));
    Span4Mux_v I__1805 (
            .O(N__15524),
            .I(N__15512));
    InMux I__1804 (
            .O(N__15521),
            .I(N__15509));
    InMux I__1803 (
            .O(N__15518),
            .I(N__15506));
    LocalMux I__1802 (
            .O(N__15515),
            .I(N__15503));
    Odrv4 I__1801 (
            .O(N__15512),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1800 (
            .O(N__15509),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1799 (
            .O(N__15506),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    Odrv4 I__1798 (
            .O(N__15503),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__1797 (
            .O(N__15494),
            .I(N__15491));
    InMux I__1796 (
            .O(N__15491),
            .I(N__15488));
    LocalMux I__1795 (
            .O(N__15488),
            .I(N__15485));
    Odrv4 I__1794 (
            .O(N__15485),
            .I(\POWERLED.un85_clk_100khz_9 ));
    InMux I__1793 (
            .O(N__15482),
            .I(N__15479));
    LocalMux I__1792 (
            .O(N__15479),
            .I(\POWERLED.mult1_un131_sum_i ));
    CascadeMux I__1791 (
            .O(N__15476),
            .I(N__15473));
    InMux I__1790 (
            .O(N__15473),
            .I(N__15470));
    LocalMux I__1789 (
            .O(N__15470),
            .I(N__15467));
    Span4Mux_v I__1788 (
            .O(N__15467),
            .I(N__15464));
    Odrv4 I__1787 (
            .O(N__15464),
            .I(\POWERLED.un85_clk_100khz_5 ));
    CascadeMux I__1786 (
            .O(N__15461),
            .I(N__15458));
    InMux I__1785 (
            .O(N__15458),
            .I(N__15455));
    LocalMux I__1784 (
            .O(N__15455),
            .I(\POWERLED.un85_clk_100khz_11 ));
    IoInMux I__1783 (
            .O(N__15452),
            .I(N__15449));
    LocalMux I__1782 (
            .O(N__15449),
            .I(N__15446));
    Span4Mux_s1_h I__1781 (
            .O(N__15446),
            .I(N__15443));
    Odrv4 I__1780 (
            .O(N__15443),
            .I(v33a_enn));
    CascadeMux I__1779 (
            .O(N__15440),
            .I(N__15435));
    CascadeMux I__1778 (
            .O(N__15439),
            .I(N__15432));
    InMux I__1777 (
            .O(N__15438),
            .I(N__15427));
    InMux I__1776 (
            .O(N__15435),
            .I(N__15424));
    InMux I__1775 (
            .O(N__15432),
            .I(N__15421));
    InMux I__1774 (
            .O(N__15431),
            .I(N__15418));
    InMux I__1773 (
            .O(N__15430),
            .I(N__15415));
    LocalMux I__1772 (
            .O(N__15427),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1771 (
            .O(N__15424),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1770 (
            .O(N__15421),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1769 (
            .O(N__15418),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1768 (
            .O(N__15415),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    CascadeMux I__1767 (
            .O(N__15404),
            .I(N__15399));
    CascadeMux I__1766 (
            .O(N__15403),
            .I(N__15396));
    CascadeMux I__1765 (
            .O(N__15402),
            .I(N__15393));
    InMux I__1764 (
            .O(N__15399),
            .I(N__15390));
    InMux I__1763 (
            .O(N__15396),
            .I(N__15385));
    InMux I__1762 (
            .O(N__15393),
            .I(N__15385));
    LocalMux I__1761 (
            .O(N__15390),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    LocalMux I__1760 (
            .O(N__15385),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    CascadeMux I__1759 (
            .O(N__15380),
            .I(N__15377));
    InMux I__1758 (
            .O(N__15377),
            .I(N__15374));
    LocalMux I__1757 (
            .O(N__15374),
            .I(\POWERLED.mult1_un124_sum_i ));
    CascadeMux I__1756 (
            .O(N__15371),
            .I(N__15368));
    InMux I__1755 (
            .O(N__15368),
            .I(N__15365));
    LocalMux I__1754 (
            .O(N__15365),
            .I(N__15362));
    Span4Mux_s1_h I__1753 (
            .O(N__15362),
            .I(N__15359));
    Odrv4 I__1752 (
            .O(N__15359),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__1751 (
            .O(N__15356),
            .I(N__15353));
    LocalMux I__1750 (
            .O(N__15353),
            .I(N__15350));
    Odrv4 I__1749 (
            .O(N__15350),
            .I(\POWERLED.un85_clk_100khz_13 ));
    InMux I__1748 (
            .O(N__15347),
            .I(N__15344));
    LocalMux I__1747 (
            .O(N__15344),
            .I(\POWERLED.N_4535_i ));
    InMux I__1746 (
            .O(N__15341),
            .I(N__15338));
    LocalMux I__1745 (
            .O(N__15338),
            .I(\POWERLED.N_4536_i ));
    InMux I__1744 (
            .O(N__15335),
            .I(N__15332));
    LocalMux I__1743 (
            .O(N__15332),
            .I(\POWERLED.N_4537_i ));
    InMux I__1742 (
            .O(N__15329),
            .I(N__15326));
    LocalMux I__1741 (
            .O(N__15326),
            .I(\POWERLED.N_4538_i ));
    CascadeMux I__1740 (
            .O(N__15323),
            .I(N__15320));
    InMux I__1739 (
            .O(N__15320),
            .I(N__15317));
    LocalMux I__1738 (
            .O(N__15317),
            .I(\POWERLED.N_4539_i ));
    CascadeMux I__1737 (
            .O(N__15314),
            .I(N__15311));
    InMux I__1736 (
            .O(N__15311),
            .I(N__15308));
    LocalMux I__1735 (
            .O(N__15308),
            .I(\POWERLED.N_4540_i ));
    CascadeMux I__1734 (
            .O(N__15305),
            .I(N__15302));
    InMux I__1733 (
            .O(N__15302),
            .I(N__15299));
    LocalMux I__1732 (
            .O(N__15299),
            .I(N__15296));
    Odrv4 I__1731 (
            .O(N__15296),
            .I(\POWERLED.N_4541_i ));
    InMux I__1730 (
            .O(N__15293),
            .I(bfn_2_11_0_));
    InMux I__1729 (
            .O(N__15290),
            .I(N__15287));
    LocalMux I__1728 (
            .O(N__15287),
            .I(N__15284));
    Odrv12 I__1727 (
            .O(N__15284),
            .I(\POWERLED.un85_clk_100khz_1 ));
    CascadeMux I__1726 (
            .O(N__15281),
            .I(N__15278));
    InMux I__1725 (
            .O(N__15278),
            .I(N__15275));
    LocalMux I__1724 (
            .O(N__15275),
            .I(\POWERLED.N_4527_i ));
    InMux I__1723 (
            .O(N__15272),
            .I(N__15269));
    LocalMux I__1722 (
            .O(N__15269),
            .I(\POWERLED.N_4528_i ));
    CascadeMux I__1721 (
            .O(N__15266),
            .I(N__15263));
    InMux I__1720 (
            .O(N__15263),
            .I(N__15260));
    LocalMux I__1719 (
            .O(N__15260),
            .I(N__15257));
    Odrv4 I__1718 (
            .O(N__15257),
            .I(\POWERLED.un85_clk_100khz_3 ));
    InMux I__1717 (
            .O(N__15254),
            .I(N__15251));
    LocalMux I__1716 (
            .O(N__15251),
            .I(\POWERLED.N_4529_i ));
    CascadeMux I__1715 (
            .O(N__15248),
            .I(N__15245));
    InMux I__1714 (
            .O(N__15245),
            .I(N__15242));
    LocalMux I__1713 (
            .O(N__15242),
            .I(N__15239));
    Span12Mux_s10_v I__1712 (
            .O(N__15239),
            .I(N__15236));
    Odrv12 I__1711 (
            .O(N__15236),
            .I(\POWERLED.un85_clk_100khz_4 ));
    InMux I__1710 (
            .O(N__15233),
            .I(N__15230));
    LocalMux I__1709 (
            .O(N__15230),
            .I(\POWERLED.N_4530_i ));
    InMux I__1708 (
            .O(N__15227),
            .I(N__15224));
    LocalMux I__1707 (
            .O(N__15224),
            .I(\POWERLED.N_4531_i ));
    CascadeMux I__1706 (
            .O(N__15221),
            .I(N__15218));
    InMux I__1705 (
            .O(N__15218),
            .I(N__15215));
    LocalMux I__1704 (
            .O(N__15215),
            .I(N__15212));
    Odrv4 I__1703 (
            .O(N__15212),
            .I(\POWERLED.un85_clk_100khz_6 ));
    InMux I__1702 (
            .O(N__15209),
            .I(N__15206));
    LocalMux I__1701 (
            .O(N__15206),
            .I(\POWERLED.N_4532_i ));
    InMux I__1700 (
            .O(N__15203),
            .I(N__15200));
    LocalMux I__1699 (
            .O(N__15200),
            .I(\POWERLED.N_4533_i ));
    InMux I__1698 (
            .O(N__15197),
            .I(N__15194));
    LocalMux I__1697 (
            .O(N__15194),
            .I(\POWERLED.N_4534_i ));
    InMux I__1696 (
            .O(N__15191),
            .I(N__15187));
    InMux I__1695 (
            .O(N__15190),
            .I(N__15184));
    LocalMux I__1694 (
            .O(N__15187),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__1693 (
            .O(N__15184),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__1692 (
            .O(N__15179),
            .I(\COUNTER.counter_1_cry_25 ));
    CascadeMux I__1691 (
            .O(N__15176),
            .I(N__15172));
    InMux I__1690 (
            .O(N__15175),
            .I(N__15169));
    InMux I__1689 (
            .O(N__15172),
            .I(N__15166));
    LocalMux I__1688 (
            .O(N__15169),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__1687 (
            .O(N__15166),
            .I(\COUNTER.counterZ0Z_27 ));
    InMux I__1686 (
            .O(N__15161),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__1685 (
            .O(N__15158),
            .I(N__15154));
    InMux I__1684 (
            .O(N__15157),
            .I(N__15151));
    LocalMux I__1683 (
            .O(N__15154),
            .I(\COUNTER.counterZ0Z_28 ));
    LocalMux I__1682 (
            .O(N__15151),
            .I(\COUNTER.counterZ0Z_28 ));
    InMux I__1681 (
            .O(N__15146),
            .I(\COUNTER.counter_1_cry_27 ));
    CascadeMux I__1680 (
            .O(N__15143),
            .I(N__15139));
    InMux I__1679 (
            .O(N__15142),
            .I(N__15136));
    InMux I__1678 (
            .O(N__15139),
            .I(N__15133));
    LocalMux I__1677 (
            .O(N__15136),
            .I(\COUNTER.counterZ0Z_29 ));
    LocalMux I__1676 (
            .O(N__15133),
            .I(\COUNTER.counterZ0Z_29 ));
    InMux I__1675 (
            .O(N__15128),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__1674 (
            .O(N__15125),
            .I(N__15121));
    InMux I__1673 (
            .O(N__15124),
            .I(N__15118));
    LocalMux I__1672 (
            .O(N__15121),
            .I(\COUNTER.counterZ0Z_30 ));
    LocalMux I__1671 (
            .O(N__15118),
            .I(\COUNTER.counterZ0Z_30 ));
    InMux I__1670 (
            .O(N__15113),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__1669 (
            .O(N__15110),
            .I(\COUNTER.counter_1_cry_30 ));
    InMux I__1668 (
            .O(N__15107),
            .I(N__15103));
    InMux I__1667 (
            .O(N__15106),
            .I(N__15100));
    LocalMux I__1666 (
            .O(N__15103),
            .I(\COUNTER.counterZ0Z_31 ));
    LocalMux I__1665 (
            .O(N__15100),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__1664 (
            .O(N__15095),
            .I(N__15092));
    LocalMux I__1663 (
            .O(N__15092),
            .I(N__15088));
    InMux I__1662 (
            .O(N__15091),
            .I(N__15084));
    Span4Mux_h I__1661 (
            .O(N__15088),
            .I(N__15081));
    InMux I__1660 (
            .O(N__15087),
            .I(N__15078));
    LocalMux I__1659 (
            .O(N__15084),
            .I(\COUNTER.counterZ0Z_6 ));
    Odrv4 I__1658 (
            .O(N__15081),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__1657 (
            .O(N__15078),
            .I(\COUNTER.counterZ0Z_6 ));
    InMux I__1656 (
            .O(N__15071),
            .I(N__15068));
    LocalMux I__1655 (
            .O(N__15068),
            .I(N__15064));
    InMux I__1654 (
            .O(N__15067),
            .I(N__15060));
    Span4Mux_h I__1653 (
            .O(N__15064),
            .I(N__15057));
    InMux I__1652 (
            .O(N__15063),
            .I(N__15054));
    LocalMux I__1651 (
            .O(N__15060),
            .I(\COUNTER.counterZ0Z_5 ));
    Odrv4 I__1650 (
            .O(N__15057),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__1649 (
            .O(N__15054),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__1648 (
            .O(N__15047),
            .I(N__15044));
    LocalMux I__1647 (
            .O(N__15044),
            .I(N__15039));
    CascadeMux I__1646 (
            .O(N__15043),
            .I(N__15036));
    InMux I__1645 (
            .O(N__15042),
            .I(N__15033));
    Span4Mux_v I__1644 (
            .O(N__15039),
            .I(N__15030));
    InMux I__1643 (
            .O(N__15036),
            .I(N__15027));
    LocalMux I__1642 (
            .O(N__15033),
            .I(\COUNTER.counterZ0Z_1 ));
    Odrv4 I__1641 (
            .O(N__15030),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__1640 (
            .O(N__15027),
            .I(\COUNTER.counterZ0Z_1 ));
    InMux I__1639 (
            .O(N__15020),
            .I(N__15016));
    InMux I__1638 (
            .O(N__15019),
            .I(N__15013));
    LocalMux I__1637 (
            .O(N__15016),
            .I(N__15010));
    LocalMux I__1636 (
            .O(N__15013),
            .I(\COUNTER.counterZ0Z_7 ));
    Odrv4 I__1635 (
            .O(N__15010),
            .I(\COUNTER.counterZ0Z_7 ));
    InMux I__1634 (
            .O(N__15005),
            .I(N__15002));
    LocalMux I__1633 (
            .O(N__15002),
            .I(\POWERLED.un1_count_cry_0_i ));
    CascadeMux I__1632 (
            .O(N__14999),
            .I(N__14995));
    InMux I__1631 (
            .O(N__14998),
            .I(N__14992));
    InMux I__1630 (
            .O(N__14995),
            .I(N__14989));
    LocalMux I__1629 (
            .O(N__14992),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__1628 (
            .O(N__14989),
            .I(\COUNTER.counterZ0Z_17 ));
    InMux I__1627 (
            .O(N__14984),
            .I(bfn_2_7_0_));
    InMux I__1626 (
            .O(N__14981),
            .I(N__14977));
    InMux I__1625 (
            .O(N__14980),
            .I(N__14974));
    LocalMux I__1624 (
            .O(N__14977),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__1623 (
            .O(N__14974),
            .I(\COUNTER.counterZ0Z_18 ));
    InMux I__1622 (
            .O(N__14969),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__1621 (
            .O(N__14966),
            .I(N__14962));
    InMux I__1620 (
            .O(N__14965),
            .I(N__14959));
    LocalMux I__1619 (
            .O(N__14962),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__1618 (
            .O(N__14959),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__1617 (
            .O(N__14954),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__1616 (
            .O(N__14951),
            .I(N__14947));
    InMux I__1615 (
            .O(N__14950),
            .I(N__14944));
    LocalMux I__1614 (
            .O(N__14947),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__1613 (
            .O(N__14944),
            .I(\COUNTER.counterZ0Z_20 ));
    InMux I__1612 (
            .O(N__14939),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__1611 (
            .O(N__14936),
            .I(N__14932));
    InMux I__1610 (
            .O(N__14935),
            .I(N__14929));
    LocalMux I__1609 (
            .O(N__14932),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__1608 (
            .O(N__14929),
            .I(\COUNTER.counterZ0Z_21 ));
    InMux I__1607 (
            .O(N__14924),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__1606 (
            .O(N__14921),
            .I(N__14917));
    InMux I__1605 (
            .O(N__14920),
            .I(N__14914));
    LocalMux I__1604 (
            .O(N__14917),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__1603 (
            .O(N__14914),
            .I(\COUNTER.counterZ0Z_22 ));
    InMux I__1602 (
            .O(N__14909),
            .I(\COUNTER.counter_1_cry_21 ));
    CascadeMux I__1601 (
            .O(N__14906),
            .I(N__14902));
    InMux I__1600 (
            .O(N__14905),
            .I(N__14899));
    InMux I__1599 (
            .O(N__14902),
            .I(N__14896));
    LocalMux I__1598 (
            .O(N__14899),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__1597 (
            .O(N__14896),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__1596 (
            .O(N__14891),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__1595 (
            .O(N__14888),
            .I(N__14884));
    InMux I__1594 (
            .O(N__14887),
            .I(N__14881));
    LocalMux I__1593 (
            .O(N__14884),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__1592 (
            .O(N__14881),
            .I(\COUNTER.counterZ0Z_24 ));
    InMux I__1591 (
            .O(N__14876),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__1590 (
            .O(N__14873),
            .I(N__14869));
    InMux I__1589 (
            .O(N__14872),
            .I(N__14866));
    LocalMux I__1588 (
            .O(N__14869),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__1587 (
            .O(N__14866),
            .I(\COUNTER.counterZ0Z_25 ));
    InMux I__1586 (
            .O(N__14861),
            .I(bfn_2_8_0_));
    CascadeMux I__1585 (
            .O(N__14858),
            .I(N__14854));
    InMux I__1584 (
            .O(N__14857),
            .I(N__14851));
    InMux I__1583 (
            .O(N__14854),
            .I(N__14848));
    LocalMux I__1582 (
            .O(N__14851),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__1581 (
            .O(N__14848),
            .I(\COUNTER.counterZ0Z_9 ));
    InMux I__1580 (
            .O(N__14843),
            .I(bfn_2_6_0_));
    InMux I__1579 (
            .O(N__14840),
            .I(N__14836));
    InMux I__1578 (
            .O(N__14839),
            .I(N__14833));
    LocalMux I__1577 (
            .O(N__14836),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__1576 (
            .O(N__14833),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__1575 (
            .O(N__14828),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__1574 (
            .O(N__14825),
            .I(N__14821));
    InMux I__1573 (
            .O(N__14824),
            .I(N__14818));
    LocalMux I__1572 (
            .O(N__14821),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__1571 (
            .O(N__14818),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__1570 (
            .O(N__14813),
            .I(\COUNTER.counter_1_cry_10 ));
    CascadeMux I__1569 (
            .O(N__14810),
            .I(N__14806));
    InMux I__1568 (
            .O(N__14809),
            .I(N__14803));
    InMux I__1567 (
            .O(N__14806),
            .I(N__14800));
    LocalMux I__1566 (
            .O(N__14803),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__1565 (
            .O(N__14800),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__1564 (
            .O(N__14795),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__1563 (
            .O(N__14792),
            .I(N__14788));
    InMux I__1562 (
            .O(N__14791),
            .I(N__14785));
    LocalMux I__1561 (
            .O(N__14788),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__1560 (
            .O(N__14785),
            .I(\COUNTER.counterZ0Z_13 ));
    InMux I__1559 (
            .O(N__14780),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__1558 (
            .O(N__14777),
            .I(N__14773));
    InMux I__1557 (
            .O(N__14776),
            .I(N__14770));
    LocalMux I__1556 (
            .O(N__14773),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__1555 (
            .O(N__14770),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__1554 (
            .O(N__14765),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__1553 (
            .O(N__14762),
            .I(N__14758));
    InMux I__1552 (
            .O(N__14761),
            .I(N__14755));
    LocalMux I__1551 (
            .O(N__14758),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__1550 (
            .O(N__14755),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__1549 (
            .O(N__14750),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__1548 (
            .O(N__14747),
            .I(N__14743));
    InMux I__1547 (
            .O(N__14746),
            .I(N__14740));
    LocalMux I__1546 (
            .O(N__14743),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__1545 (
            .O(N__14740),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__1544 (
            .O(N__14735),
            .I(\COUNTER.counter_1_cry_15 ));
    CascadeMux I__1543 (
            .O(N__14732),
            .I(N__14729));
    InMux I__1542 (
            .O(N__14729),
            .I(N__14726));
    LocalMux I__1541 (
            .O(N__14726),
            .I(N__14720));
    InMux I__1540 (
            .O(N__14725),
            .I(N__14713));
    InMux I__1539 (
            .O(N__14724),
            .I(N__14713));
    InMux I__1538 (
            .O(N__14723),
            .I(N__14713));
    Odrv4 I__1537 (
            .O(N__14720),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__1536 (
            .O(N__14713),
            .I(\COUNTER.counterZ0Z_0 ));
    InMux I__1535 (
            .O(N__14708),
            .I(N__14705));
    LocalMux I__1534 (
            .O(N__14705),
            .I(N__14700));
    InMux I__1533 (
            .O(N__14704),
            .I(N__14695));
    InMux I__1532 (
            .O(N__14703),
            .I(N__14695));
    Odrv4 I__1531 (
            .O(N__14700),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__1530 (
            .O(N__14695),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__1529 (
            .O(N__14690),
            .I(N__14687));
    LocalMux I__1528 (
            .O(N__14687),
            .I(N__14684));
    Span4Mux_v I__1527 (
            .O(N__14684),
            .I(N__14681));
    Odrv4 I__1526 (
            .O(N__14681),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__1525 (
            .O(N__14678),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__1524 (
            .O(N__14675),
            .I(N__14671));
    CascadeMux I__1523 (
            .O(N__14674),
            .I(N__14667));
    LocalMux I__1522 (
            .O(N__14671),
            .I(N__14664));
    InMux I__1521 (
            .O(N__14670),
            .I(N__14659));
    InMux I__1520 (
            .O(N__14667),
            .I(N__14659));
    Odrv4 I__1519 (
            .O(N__14664),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__1518 (
            .O(N__14659),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__1517 (
            .O(N__14654),
            .I(N__14651));
    LocalMux I__1516 (
            .O(N__14651),
            .I(N__14648));
    Odrv4 I__1515 (
            .O(N__14648),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__1514 (
            .O(N__14645),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__1513 (
            .O(N__14642),
            .I(N__14639));
    LocalMux I__1512 (
            .O(N__14639),
            .I(N__14635));
    InMux I__1511 (
            .O(N__14638),
            .I(N__14631));
    Span4Mux_h I__1510 (
            .O(N__14635),
            .I(N__14628));
    InMux I__1509 (
            .O(N__14634),
            .I(N__14625));
    LocalMux I__1508 (
            .O(N__14631),
            .I(\COUNTER.counterZ0Z_4 ));
    Odrv4 I__1507 (
            .O(N__14628),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__1506 (
            .O(N__14625),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__1505 (
            .O(N__14618),
            .I(N__14615));
    LocalMux I__1504 (
            .O(N__14615),
            .I(N__14612));
    Span4Mux_v I__1503 (
            .O(N__14612),
            .I(N__14609));
    Odrv4 I__1502 (
            .O(N__14609),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__1501 (
            .O(N__14606),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__1500 (
            .O(N__14603),
            .I(N__14600));
    LocalMux I__1499 (
            .O(N__14600),
            .I(N__14597));
    Odrv4 I__1498 (
            .O(N__14597),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__1497 (
            .O(N__14594),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__1496 (
            .O(N__14591),
            .I(N__14588));
    LocalMux I__1495 (
            .O(N__14588),
            .I(N__14585));
    Span4Mux_v I__1494 (
            .O(N__14585),
            .I(N__14582));
    Odrv4 I__1493 (
            .O(N__14582),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__1492 (
            .O(N__14579),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__1491 (
            .O(N__14576),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__1490 (
            .O(N__14573),
            .I(N__14569));
    InMux I__1489 (
            .O(N__14572),
            .I(N__14566));
    LocalMux I__1488 (
            .O(N__14569),
            .I(N__14563));
    LocalMux I__1487 (
            .O(N__14566),
            .I(\COUNTER.counterZ0Z_8 ));
    Odrv4 I__1486 (
            .O(N__14563),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__1485 (
            .O(N__14558),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__1484 (
            .O(N__14555),
            .I(N__14551));
    InMux I__1483 (
            .O(N__14554),
            .I(N__14548));
    LocalMux I__1482 (
            .O(N__14551),
            .I(\DSW_PWRGD.countZ0Z_9 ));
    LocalMux I__1481 (
            .O(N__14548),
            .I(\DSW_PWRGD.countZ0Z_9 ));
    InMux I__1480 (
            .O(N__14543),
            .I(N__14539));
    InMux I__1479 (
            .O(N__14542),
            .I(N__14536));
    LocalMux I__1478 (
            .O(N__14539),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    LocalMux I__1477 (
            .O(N__14536),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    CascadeMux I__1476 (
            .O(N__14531),
            .I(N__14528));
    InMux I__1475 (
            .O(N__14528),
            .I(N__14524));
    InMux I__1474 (
            .O(N__14527),
            .I(N__14521));
    LocalMux I__1473 (
            .O(N__14524),
            .I(N__14518));
    LocalMux I__1472 (
            .O(N__14521),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    Odrv4 I__1471 (
            .O(N__14518),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    InMux I__1470 (
            .O(N__14513),
            .I(N__14509));
    InMux I__1469 (
            .O(N__14512),
            .I(N__14506));
    LocalMux I__1468 (
            .O(N__14509),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    LocalMux I__1467 (
            .O(N__14506),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    CascadeMux I__1466 (
            .O(N__14501),
            .I(\PCH_PWRGD.N_2126_i_cascade_ ));
    CascadeMux I__1465 (
            .O(N__14498),
            .I(\PCH_PWRGD.N_381_cascade_ ));
    InMux I__1464 (
            .O(N__14495),
            .I(N__14489));
    InMux I__1463 (
            .O(N__14494),
            .I(N__14489));
    LocalMux I__1462 (
            .O(N__14489),
            .I(\PCH_PWRGD.N_254_0 ));
    InMux I__1461 (
            .O(N__14486),
            .I(N__14482));
    InMux I__1460 (
            .O(N__14485),
            .I(N__14479));
    LocalMux I__1459 (
            .O(N__14482),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    LocalMux I__1458 (
            .O(N__14479),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    InMux I__1457 (
            .O(N__14474),
            .I(N__14470));
    InMux I__1456 (
            .O(N__14473),
            .I(N__14467));
    LocalMux I__1455 (
            .O(N__14470),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    LocalMux I__1454 (
            .O(N__14467),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    CascadeMux I__1453 (
            .O(N__14462),
            .I(N__14458));
    InMux I__1452 (
            .O(N__14461),
            .I(N__14455));
    InMux I__1451 (
            .O(N__14458),
            .I(N__14452));
    LocalMux I__1450 (
            .O(N__14455),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    LocalMux I__1449 (
            .O(N__14452),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    InMux I__1448 (
            .O(N__14447),
            .I(N__14443));
    InMux I__1447 (
            .O(N__14446),
            .I(N__14440));
    LocalMux I__1446 (
            .O(N__14443),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    LocalMux I__1445 (
            .O(N__14440),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    InMux I__1444 (
            .O(N__14435),
            .I(N__14432));
    LocalMux I__1443 (
            .O(N__14432),
            .I(\DSW_PWRGD.un4_count_11 ));
    InMux I__1442 (
            .O(N__14429),
            .I(N__14426));
    LocalMux I__1441 (
            .O(N__14426),
            .I(\DSW_PWRGD.un4_count_10 ));
    CascadeMux I__1440 (
            .O(N__14423),
            .I(\DSW_PWRGD.un4_count_8_cascade_ ));
    InMux I__1439 (
            .O(N__14420),
            .I(N__14417));
    LocalMux I__1438 (
            .O(N__14417),
            .I(\DSW_PWRGD.un4_count_9 ));
    CascadeMux I__1437 (
            .O(N__14414),
            .I(N__14409));
    CascadeMux I__1436 (
            .O(N__14413),
            .I(N__14406));
    InMux I__1435 (
            .O(N__14412),
            .I(N__14399));
    InMux I__1434 (
            .O(N__14409),
            .I(N__14399));
    InMux I__1433 (
            .O(N__14406),
            .I(N__14399));
    LocalMux I__1432 (
            .O(N__14399),
            .I(N__14396));
    Odrv4 I__1431 (
            .O(N__14396),
            .I(\DSW_PWRGD.N_1_i ));
    InMux I__1430 (
            .O(N__14393),
            .I(N__14390));
    LocalMux I__1429 (
            .O(N__14390),
            .I(\PCH_PWRGD.N_381 ));
    InMux I__1428 (
            .O(N__14387),
            .I(N__14383));
    InMux I__1427 (
            .O(N__14386),
            .I(N__14380));
    LocalMux I__1426 (
            .O(N__14383),
            .I(\PCH_PWRGD.N_2126_i ));
    LocalMux I__1425 (
            .O(N__14380),
            .I(\PCH_PWRGD.N_2126_i ));
    CascadeMux I__1424 (
            .O(N__14375),
            .I(N__14372));
    InMux I__1423 (
            .O(N__14372),
            .I(N__14366));
    InMux I__1422 (
            .O(N__14371),
            .I(N__14361));
    InMux I__1421 (
            .O(N__14370),
            .I(N__14361));
    InMux I__1420 (
            .O(N__14369),
            .I(N__14358));
    LocalMux I__1419 (
            .O(N__14366),
            .I(N__14351));
    LocalMux I__1418 (
            .O(N__14361),
            .I(N__14351));
    LocalMux I__1417 (
            .O(N__14358),
            .I(N__14351));
    Span12Mux_s8_v I__1416 (
            .O(N__14351),
            .I(N__14348));
    Odrv12 I__1415 (
            .O(N__14348),
            .I(vr_ready_vccin));
    CascadeMux I__1414 (
            .O(N__14345),
            .I(\PCH_PWRGD.N_255_0_cascade_ ));
    CascadeMux I__1413 (
            .O(N__14342),
            .I(\PCH_PWRGD.count_RNIZ0Z_1_cascade_ ));
    CascadeMux I__1412 (
            .O(N__14339),
            .I(N__14336));
    InMux I__1411 (
            .O(N__14336),
            .I(N__14333));
    LocalMux I__1410 (
            .O(N__14333),
            .I(\PCH_PWRGD.count_0_1 ));
    InMux I__1409 (
            .O(N__14330),
            .I(N__14326));
    InMux I__1408 (
            .O(N__14329),
            .I(N__14323));
    LocalMux I__1407 (
            .O(N__14326),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    LocalMux I__1406 (
            .O(N__14323),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    InMux I__1405 (
            .O(N__14318),
            .I(N__14314));
    InMux I__1404 (
            .O(N__14317),
            .I(N__14311));
    LocalMux I__1403 (
            .O(N__14314),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    LocalMux I__1402 (
            .O(N__14311),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    CascadeMux I__1401 (
            .O(N__14306),
            .I(N__14302));
    InMux I__1400 (
            .O(N__14305),
            .I(N__14299));
    InMux I__1399 (
            .O(N__14302),
            .I(N__14296));
    LocalMux I__1398 (
            .O(N__14299),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    LocalMux I__1397 (
            .O(N__14296),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    InMux I__1396 (
            .O(N__14291),
            .I(N__14287));
    InMux I__1395 (
            .O(N__14290),
            .I(N__14284));
    LocalMux I__1394 (
            .O(N__14287),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    LocalMux I__1393 (
            .O(N__14284),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    InMux I__1392 (
            .O(N__14279),
            .I(N__14273));
    InMux I__1391 (
            .O(N__14278),
            .I(N__14273));
    LocalMux I__1390 (
            .O(N__14273),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    CascadeMux I__1389 (
            .O(N__14270),
            .I(\PCH_PWRGD.curr_state_RNI3DJUZ0Z_0_cascade_ ));
    InMux I__1388 (
            .O(N__14267),
            .I(N__14263));
    InMux I__1387 (
            .O(N__14266),
            .I(N__14260));
    LocalMux I__1386 (
            .O(N__14263),
            .I(N__14257));
    LocalMux I__1385 (
            .O(N__14260),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    Odrv4 I__1384 (
            .O(N__14257),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    InMux I__1383 (
            .O(N__14252),
            .I(N__14248));
    InMux I__1382 (
            .O(N__14251),
            .I(N__14245));
    LocalMux I__1381 (
            .O(N__14248),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    LocalMux I__1380 (
            .O(N__14245),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    CascadeMux I__1379 (
            .O(N__14240),
            .I(N__14236));
    InMux I__1378 (
            .O(N__14239),
            .I(N__14233));
    InMux I__1377 (
            .O(N__14236),
            .I(N__14230));
    LocalMux I__1376 (
            .O(N__14233),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    LocalMux I__1375 (
            .O(N__14230),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    InMux I__1374 (
            .O(N__14225),
            .I(N__14221));
    InMux I__1373 (
            .O(N__14224),
            .I(N__14218));
    LocalMux I__1372 (
            .O(N__14221),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    LocalMux I__1371 (
            .O(N__14218),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    InMux I__1370 (
            .O(N__14213),
            .I(N__14210));
    LocalMux I__1369 (
            .O(N__14210),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__1368 (
            .O(N__14207),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    InMux I__1367 (
            .O(N__14204),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    CascadeMux I__1366 (
            .O(N__14201),
            .I(\POWERLED.mult1_un103_sum_s_8_cascade_ ));
    CascadeMux I__1365 (
            .O(N__14198),
            .I(N__14193));
    CascadeMux I__1364 (
            .O(N__14197),
            .I(N__14190));
    CascadeMux I__1363 (
            .O(N__14196),
            .I(N__14187));
    InMux I__1362 (
            .O(N__14193),
            .I(N__14184));
    InMux I__1361 (
            .O(N__14190),
            .I(N__14179));
    InMux I__1360 (
            .O(N__14187),
            .I(N__14179));
    LocalMux I__1359 (
            .O(N__14184),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    LocalMux I__1358 (
            .O(N__14179),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    CascadeMux I__1357 (
            .O(N__14174),
            .I(\PCH_PWRGD.count_rst_6_cascade_ ));
    CascadeMux I__1356 (
            .O(N__14171),
            .I(\PCH_PWRGD.count_rst_14_cascade_ ));
    CascadeMux I__1355 (
            .O(N__14168),
            .I(\PCH_PWRGD.countZ0Z_0_cascade_ ));
    InMux I__1354 (
            .O(N__14165),
            .I(N__14162));
    LocalMux I__1353 (
            .O(N__14162),
            .I(\PCH_PWRGD.count_RNIZ0Z_1 ));
    InMux I__1352 (
            .O(N__14159),
            .I(N__14156));
    LocalMux I__1351 (
            .O(N__14156),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__1350 (
            .O(N__14153),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    InMux I__1349 (
            .O(N__14150),
            .I(N__14147));
    LocalMux I__1348 (
            .O(N__14147),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__1347 (
            .O(N__14144),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__1346 (
            .O(N__14141),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    InMux I__1345 (
            .O(N__14138),
            .I(N__14135));
    LocalMux I__1344 (
            .O(N__14135),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__1343 (
            .O(N__14132),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    InMux I__1342 (
            .O(N__14129),
            .I(N__14126));
    LocalMux I__1341 (
            .O(N__14126),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__1340 (
            .O(N__14123),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    InMux I__1339 (
            .O(N__14120),
            .I(N__14117));
    LocalMux I__1338 (
            .O(N__14117),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__1337 (
            .O(N__14114),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    InMux I__1336 (
            .O(N__14111),
            .I(N__14108));
    LocalMux I__1335 (
            .O(N__14108),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__1334 (
            .O(N__14105),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__1333 (
            .O(N__14102),
            .I(N__14099));
    LocalMux I__1332 (
            .O(N__14099),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__1331 (
            .O(N__14096),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    InMux I__1330 (
            .O(N__14093),
            .I(N__14090));
    LocalMux I__1329 (
            .O(N__14090),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__1328 (
            .O(N__14087),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    InMux I__1327 (
            .O(N__14084),
            .I(N__14081));
    LocalMux I__1326 (
            .O(N__14081),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__1325 (
            .O(N__14078),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__1324 (
            .O(N__14075),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    CascadeMux I__1323 (
            .O(N__14072),
            .I(\POWERLED.mult1_un117_sum_s_8_cascade_ ));
    CascadeMux I__1322 (
            .O(N__14069),
            .I(N__14064));
    CascadeMux I__1321 (
            .O(N__14068),
            .I(N__14061));
    CascadeMux I__1320 (
            .O(N__14067),
            .I(N__14058));
    InMux I__1319 (
            .O(N__14064),
            .I(N__14055));
    InMux I__1318 (
            .O(N__14061),
            .I(N__14050));
    InMux I__1317 (
            .O(N__14058),
            .I(N__14050));
    LocalMux I__1316 (
            .O(N__14055),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    LocalMux I__1315 (
            .O(N__14050),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    InMux I__1314 (
            .O(N__14045),
            .I(N__14042));
    LocalMux I__1313 (
            .O(N__14042),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__1312 (
            .O(N__14039),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    InMux I__1311 (
            .O(N__14036),
            .I(N__14033));
    LocalMux I__1310 (
            .O(N__14033),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__1309 (
            .O(N__14030),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    InMux I__1308 (
            .O(N__14027),
            .I(N__14024));
    LocalMux I__1307 (
            .O(N__14024),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__1306 (
            .O(N__14021),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__1305 (
            .O(N__14018),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__1304 (
            .O(N__14015),
            .I(N__14012));
    LocalMux I__1303 (
            .O(N__14012),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__1302 (
            .O(N__14009),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    InMux I__1301 (
            .O(N__14006),
            .I(N__14003));
    LocalMux I__1300 (
            .O(N__14003),
            .I(N__13999));
    InMux I__1299 (
            .O(N__14002),
            .I(N__13996));
    Odrv12 I__1298 (
            .O(N__13999),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    LocalMux I__1297 (
            .O(N__13996),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__1296 (
            .O(N__13991),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    InMux I__1295 (
            .O(N__13988),
            .I(N__13985));
    LocalMux I__1294 (
            .O(N__13985),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__1293 (
            .O(N__13982),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__1292 (
            .O(N__13979),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    InMux I__1291 (
            .O(N__13976),
            .I(N__13968));
    InMux I__1290 (
            .O(N__13975),
            .I(N__13968));
    CascadeMux I__1289 (
            .O(N__13974),
            .I(N__13965));
    CascadeMux I__1288 (
            .O(N__13973),
            .I(N__13962));
    LocalMux I__1287 (
            .O(N__13968),
            .I(N__13957));
    InMux I__1286 (
            .O(N__13965),
            .I(N__13954));
    InMux I__1285 (
            .O(N__13962),
            .I(N__13949));
    InMux I__1284 (
            .O(N__13961),
            .I(N__13949));
    InMux I__1283 (
            .O(N__13960),
            .I(N__13946));
    Odrv12 I__1282 (
            .O(N__13957),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__1281 (
            .O(N__13954),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__1280 (
            .O(N__13949),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__1279 (
            .O(N__13946),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    CascadeMux I__1278 (
            .O(N__13937),
            .I(\POWERLED.mult1_un124_sum_s_8_cascade_ ));
    InMux I__1277 (
            .O(N__13934),
            .I(N__13931));
    LocalMux I__1276 (
            .O(N__13931),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__1275 (
            .O(N__13928),
            .I(N__13925));
    LocalMux I__1274 (
            .O(N__13925),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__1273 (
            .O(N__13922),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    InMux I__1272 (
            .O(N__13919),
            .I(N__13916));
    LocalMux I__1271 (
            .O(N__13916),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__1270 (
            .O(N__13913),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__1269 (
            .O(N__13910),
            .I(N__13907));
    LocalMux I__1268 (
            .O(N__13907),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__1267 (
            .O(N__13904),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    InMux I__1266 (
            .O(N__13901),
            .I(N__13898));
    LocalMux I__1265 (
            .O(N__13898),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__1264 (
            .O(N__13895),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    InMux I__1263 (
            .O(N__13892),
            .I(N__13889));
    LocalMux I__1262 (
            .O(N__13889),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    InMux I__1261 (
            .O(N__13886),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    CascadeMux I__1260 (
            .O(N__13883),
            .I(N__13880));
    InMux I__1259 (
            .O(N__13880),
            .I(N__13877));
    LocalMux I__1258 (
            .O(N__13877),
            .I(N__13874));
    Odrv4 I__1257 (
            .O(N__13874),
            .I(\POWERLED.mult1_un131_sum_axb_7_l_fx ));
    InMux I__1256 (
            .O(N__13871),
            .I(N__13868));
    LocalMux I__1255 (
            .O(N__13868),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__1254 (
            .O(N__13865),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__1253 (
            .O(N__13862),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__1252 (
            .O(N__13859),
            .I(N__13856));
    InMux I__1251 (
            .O(N__13856),
            .I(N__13853));
    LocalMux I__1250 (
            .O(N__13853),
            .I(\POWERLED.mult1_un131_sum_axb_4_l_fx ));
    InMux I__1249 (
            .O(N__13850),
            .I(N__13844));
    InMux I__1248 (
            .O(N__13849),
            .I(N__13844));
    LocalMux I__1247 (
            .O(N__13844),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__1246 (
            .O(N__13841),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    InMux I__1245 (
            .O(N__13838),
            .I(N__13835));
    LocalMux I__1244 (
            .O(N__13835),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__1243 (
            .O(N__13832),
            .I(N__13829));
    LocalMux I__1242 (
            .O(N__13829),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__1241 (
            .O(N__13826),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    InMux I__1240 (
            .O(N__13823),
            .I(N__13820));
    LocalMux I__1239 (
            .O(N__13820),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__1238 (
            .O(N__13817),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    InMux I__1237 (
            .O(N__13814),
            .I(N__13811));
    LocalMux I__1236 (
            .O(N__13811),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__1235 (
            .O(N__13808),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    CascadeMux I__1234 (
            .O(N__13805),
            .I(N__13802));
    InMux I__1233 (
            .O(N__13802),
            .I(N__13799));
    LocalMux I__1232 (
            .O(N__13799),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    InMux I__1231 (
            .O(N__13796),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    InMux I__1230 (
            .O(N__13793),
            .I(N__13790));
    LocalMux I__1229 (
            .O(N__13790),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__1228 (
            .O(N__13787),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    InMux I__1227 (
            .O(N__13784),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    CascadeMux I__1226 (
            .O(N__13781),
            .I(N__13777));
    CascadeMux I__1225 (
            .O(N__13780),
            .I(N__13774));
    InMux I__1224 (
            .O(N__13777),
            .I(N__13769));
    InMux I__1223 (
            .O(N__13774),
            .I(N__13764));
    InMux I__1222 (
            .O(N__13773),
            .I(N__13764));
    InMux I__1221 (
            .O(N__13772),
            .I(N__13761));
    LocalMux I__1220 (
            .O(N__13769),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__1219 (
            .O(N__13764),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__1218 (
            .O(N__13761),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__1217 (
            .O(N__13754),
            .I(\POWERLED.mult1_un138_sum_s_8_cascade_ ));
    InMux I__1216 (
            .O(N__13751),
            .I(N__13748));
    LocalMux I__1215 (
            .O(N__13748),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__1214 (
            .O(N__13745),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__1213 (
            .O(N__13742),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    InMux I__1212 (
            .O(N__13739),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    InMux I__1211 (
            .O(N__13736),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    InMux I__1210 (
            .O(N__13733),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    InMux I__1209 (
            .O(N__13730),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    InMux I__1208 (
            .O(N__13727),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    CascadeMux I__1207 (
            .O(N__13724),
            .I(N__13720));
    InMux I__1206 (
            .O(N__13723),
            .I(N__13712));
    InMux I__1205 (
            .O(N__13720),
            .I(N__13712));
    InMux I__1204 (
            .O(N__13719),
            .I(N__13712));
    LocalMux I__1203 (
            .O(N__13712),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    InMux I__1202 (
            .O(N__13709),
            .I(bfn_1_4_0_));
    CascadeMux I__1201 (
            .O(N__13706),
            .I(N__13702));
    InMux I__1200 (
            .O(N__13705),
            .I(N__13699));
    InMux I__1199 (
            .O(N__13702),
            .I(N__13696));
    LocalMux I__1198 (
            .O(N__13699),
            .I(N__13691));
    LocalMux I__1197 (
            .O(N__13696),
            .I(N__13691));
    Odrv12 I__1196 (
            .O(N__13691),
            .I(\DSW_PWRGD.un1_curr_state10_0 ));
    InMux I__1195 (
            .O(N__13688),
            .I(N__13673));
    InMux I__1194 (
            .O(N__13687),
            .I(N__13673));
    InMux I__1193 (
            .O(N__13686),
            .I(N__13673));
    InMux I__1192 (
            .O(N__13685),
            .I(N__13673));
    InMux I__1191 (
            .O(N__13684),
            .I(N__13673));
    LocalMux I__1190 (
            .O(N__13673),
            .I(N__13670));
    IoSpan4Mux I__1189 (
            .O(N__13670),
            .I(N__13667));
    IoSpan4Mux I__1188 (
            .O(N__13667),
            .I(N__13664));
    Odrv4 I__1187 (
            .O(N__13664),
            .I(v33dsw_ok));
    InMux I__1186 (
            .O(N__13661),
            .I(N__13646));
    InMux I__1185 (
            .O(N__13660),
            .I(N__13646));
    InMux I__1184 (
            .O(N__13659),
            .I(N__13646));
    InMux I__1183 (
            .O(N__13658),
            .I(N__13646));
    InMux I__1182 (
            .O(N__13657),
            .I(N__13646));
    LocalMux I__1181 (
            .O(N__13646),
            .I(\DSW_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__1180 (
            .O(N__13643),
            .I(N__13638));
    InMux I__1179 (
            .O(N__13642),
            .I(N__13627));
    InMux I__1178 (
            .O(N__13641),
            .I(N__13627));
    InMux I__1177 (
            .O(N__13638),
            .I(N__13627));
    InMux I__1176 (
            .O(N__13637),
            .I(N__13627));
    InMux I__1175 (
            .O(N__13636),
            .I(N__13624));
    LocalMux I__1174 (
            .O(N__13627),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__1173 (
            .O(N__13624),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__1172 (
            .O(N__13619),
            .I(DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_));
    SRMux I__1171 (
            .O(N__13616),
            .I(N__13611));
    SRMux I__1170 (
            .O(N__13615),
            .I(N__13608));
    SRMux I__1169 (
            .O(N__13614),
            .I(N__13605));
    LocalMux I__1168 (
            .O(N__13611),
            .I(N__13602));
    LocalMux I__1167 (
            .O(N__13608),
            .I(N__13599));
    LocalMux I__1166 (
            .O(N__13605),
            .I(N__13596));
    Span4Mux_s3_v I__1165 (
            .O(N__13602),
            .I(N__13591));
    Span4Mux_s1_h I__1164 (
            .O(N__13599),
            .I(N__13591));
    Odrv4 I__1163 (
            .O(N__13596),
            .I(G_27));
    Odrv4 I__1162 (
            .O(N__13591),
            .I(G_27));
    CascadeMux I__1161 (
            .O(N__13586),
            .I(G_27_cascade_));
    CEMux I__1160 (
            .O(N__13583),
            .I(N__13580));
    LocalMux I__1159 (
            .O(N__13580),
            .I(N__13577));
    Odrv4 I__1158 (
            .O(N__13577),
            .I(\DSW_PWRGD.N_27_1 ));
    InMux I__1157 (
            .O(N__13574),
            .I(\DSW_PWRGD.un1_count_1_cry_5 ));
    InMux I__1156 (
            .O(N__13571),
            .I(\DSW_PWRGD.un1_count_1_cry_6 ));
    InMux I__1155 (
            .O(N__13568),
            .I(bfn_1_3_0_));
    InMux I__1154 (
            .O(N__13565),
            .I(\DSW_PWRGD.un1_count_1_cry_8 ));
    InMux I__1153 (
            .O(N__13562),
            .I(\DSW_PWRGD.un1_count_1_cry_9 ));
    InMux I__1152 (
            .O(N__13559),
            .I(\DSW_PWRGD.un1_count_1_cry_10 ));
    InMux I__1151 (
            .O(N__13556),
            .I(\DSW_PWRGD.un1_count_1_cry_11 ));
    InMux I__1150 (
            .O(N__13553),
            .I(\DSW_PWRGD.un1_count_1_cry_12 ));
    InMux I__1149 (
            .O(N__13550),
            .I(\DSW_PWRGD.un1_count_1_cry_13 ));
    InMux I__1148 (
            .O(N__13547),
            .I(\DSW_PWRGD.un1_count_1_cry_0 ));
    InMux I__1147 (
            .O(N__13544),
            .I(\DSW_PWRGD.un1_count_1_cry_1 ));
    InMux I__1146 (
            .O(N__13541),
            .I(\DSW_PWRGD.un1_count_1_cry_2 ));
    InMux I__1145 (
            .O(N__13538),
            .I(\DSW_PWRGD.un1_count_1_cry_3 ));
    InMux I__1144 (
            .O(N__13535),
            .I(\DSW_PWRGD.un1_count_1_cry_4 ));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(\POWERLED.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(\POWERLED.un1_count_cry_8 ),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\PCH_PWRGD.un2_count_1_cry_8 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(COUNTER_un4_counter_7),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_2_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_5_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_7_cZ0 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_7 ),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_15 ),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_1_4_0_));
    ICE_GB N_579_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__23806),
            .GLOBALBUFFEROUTPUT(N_579_g));
    ICE_GB N_27_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__25922),
            .GLOBALBUFFEROUTPUT(N_27_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \DSW_PWRGD.count_0_LC_1_2_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_0_LC_1_2_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_0_LC_1_2_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_0_LC_1_2_0  (
            .in0(N__29557),
            .in1(N__14305),
            .in2(N__13706),
            .in3(N__13705),
            .lcout(\DSW_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_0 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_1_LC_1_2_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_1_LC_1_2_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_1_LC_1_2_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_1_LC_1_2_1  (
            .in0(N__29553),
            .in1(N__14291),
            .in2(_gnd_net_),
            .in3(N__13547),
            .lcout(\DSW_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_0 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_1 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_2_LC_1_2_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_2_LC_1_2_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_2_LC_1_2_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_2_LC_1_2_2  (
            .in0(N__29558),
            .in1(N__14513),
            .in2(_gnd_net_),
            .in3(N__13544),
            .lcout(\DSW_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_1 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_2 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_3_LC_1_2_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_3_LC_1_2_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_3_LC_1_2_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_3_LC_1_2_3  (
            .in0(N__29554),
            .in1(N__14330),
            .in2(_gnd_net_),
            .in3(N__13541),
            .lcout(\DSW_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_2 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_3 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_4_LC_1_2_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_4_LC_1_2_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_4_LC_1_2_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_4_LC_1_2_4  (
            .in0(N__29559),
            .in1(N__14318),
            .in2(_gnd_net_),
            .in3(N__13538),
            .lcout(\DSW_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_3 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_4 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_5_LC_1_2_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_5_LC_1_2_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_5_LC_1_2_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_5_LC_1_2_5  (
            .in0(N__29555),
            .in1(N__14225),
            .in2(_gnd_net_),
            .in3(N__13535),
            .lcout(\DSW_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_4 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_5 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_6_LC_1_2_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_6_LC_1_2_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_6_LC_1_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_6_LC_1_2_6  (
            .in0(N__29560),
            .in1(N__14239),
            .in2(_gnd_net_),
            .in3(N__13574),
            .lcout(\DSW_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_5 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_6 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_7_LC_1_2_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_7_LC_1_2_7 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_7_LC_1_2_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_7_LC_1_2_7  (
            .in0(N__29556),
            .in1(N__14543),
            .in2(_gnd_net_),
            .in3(N__13571),
            .lcout(\DSW_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_6 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_7 ),
            .clk(N__32928),
            .ce(),
            .sr(N__13616));
    defparam \DSW_PWRGD.count_8_LC_1_3_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_8_LC_1_3_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_8_LC_1_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_8_LC_1_3_0  (
            .in0(N__29574),
            .in1(N__14527),
            .in2(_gnd_net_),
            .in3(N__13568),
            .lcout(\DSW_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_8 ),
            .clk(N__32973),
            .ce(),
            .sr(N__13614));
    defparam \DSW_PWRGD.count_9_LC_1_3_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_9_LC_1_3_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_9_LC_1_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_9_LC_1_3_1  (
            .in0(N__29570),
            .in1(N__14555),
            .in2(_gnd_net_),
            .in3(N__13565),
            .lcout(\DSW_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_8 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_9 ),
            .clk(N__32973),
            .ce(),
            .sr(N__13614));
    defparam \DSW_PWRGD.count_10_LC_1_3_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_10_LC_1_3_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_10_LC_1_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_10_LC_1_3_2  (
            .in0(N__29571),
            .in1(N__14252),
            .in2(_gnd_net_),
            .in3(N__13562),
            .lcout(\DSW_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_9 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_10 ),
            .clk(N__32973),
            .ce(),
            .sr(N__13614));
    defparam \DSW_PWRGD.count_11_LC_1_3_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_11_LC_1_3_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_11_LC_1_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_11_LC_1_3_3  (
            .in0(N__29568),
            .in1(N__14266),
            .in2(_gnd_net_),
            .in3(N__13559),
            .lcout(\DSW_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_10 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_11 ),
            .clk(N__32973),
            .ce(),
            .sr(N__13614));
    defparam \DSW_PWRGD.count_12_LC_1_3_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_12_LC_1_3_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_12_LC_1_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_12_LC_1_3_4  (
            .in0(N__29572),
            .in1(N__14486),
            .in2(_gnd_net_),
            .in3(N__13556),
            .lcout(\DSW_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_11 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_12 ),
            .clk(N__32973),
            .ce(),
            .sr(N__13614));
    defparam \DSW_PWRGD.count_13_LC_1_3_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_13_LC_1_3_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_13_LC_1_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_13_LC_1_3_5  (
            .in0(N__29569),
            .in1(N__14474),
            .in2(_gnd_net_),
            .in3(N__13553),
            .lcout(\DSW_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_12 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_13 ),
            .clk(N__32973),
            .ce(),
            .sr(N__13614));
    defparam \DSW_PWRGD.count_14_LC_1_3_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_14_LC_1_3_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_14_LC_1_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_14_LC_1_3_6  (
            .in0(N__29573),
            .in1(N__14461),
            .in2(_gnd_net_),
            .in3(N__13550),
            .lcout(\DSW_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_13 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14 ),
            .clk(N__32973),
            .ce(),
            .sr(N__13614));
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_3_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_3_7  (
            .in0(_gnd_net_),
            .in1(N__27470),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_14 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_15_LC_1_4_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_15_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_esr_15_LC_1_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DSW_PWRGD.count_esr_15_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(N__14447),
            .in2(_gnd_net_),
            .in3(N__13709),
            .lcout(\DSW_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32959),
            .ce(N__13583),
            .sr(N__13615));
    defparam \DSW_PWRGD.DSW_PWROK_LC_1_5_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.DSW_PWROK_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.DSW_PWROK_LC_1_5_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \DSW_PWRGD.DSW_PWROK_LC_1_5_1  (
            .in0(N__13684),
            .in1(N__13659),
            .in2(_gnd_net_),
            .in3(N__13641),
            .lcout(dsw_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32974),
            .ce(N__29408),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_1_5_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_1_5_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \DSW_PWRGD.curr_state_RNIADII_0_LC_1_5_2  (
            .in0(N__13658),
            .in1(N__13636),
            .in2(_gnd_net_),
            .in3(N__13687),
            .lcout(\DSW_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_0_LC_1_5_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_0_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_0_LC_1_5_3 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \DSW_PWRGD.curr_state_0_LC_1_5_3  (
            .in0(N__13685),
            .in1(N__13660),
            .in2(N__14414),
            .in3(N__13642),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32974),
            .ce(N__29408),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_1_LC_1_5_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_1_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_1_LC_1_5_4 .LUT_INIT=16'b0000010000001110;
    LogicCell40 \DSW_PWRGD.curr_state_1_LC_1_5_4  (
            .in0(N__13661),
            .in1(N__13686),
            .in2(N__13643),
            .in3(N__14412),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32974),
            .ce(N__29408),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_1_5_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_1_5_5 .LUT_INIT=16'b1111111100011101;
    LogicCell40 \DSW_PWRGD.curr_state_RNILLF15_0_LC_1_5_5  (
            .in0(N__13688),
            .in1(N__13657),
            .in2(N__14413),
            .in3(N__13637),
            .lcout(),
            .ltout(DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.G_27_LC_1_5_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.G_27_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.G_27_LC_1_5_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \VPP_VDDQ.G_27_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13619),
            .in3(N__29541),
            .lcout(G_27),
            .ltout(G_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_1_5_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_1_5_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \DSW_PWRGD.count_esr_RNO_0_15_LC_1_5_7  (
            .in0(N__29542),
            .in1(_gnd_net_),
            .in2(N__13586),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.N_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_1_7_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_1_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_1_7_0  (
            .in0(N__14824),
            .in1(N__14839),
            .in2(N__14858),
            .in3(N__14573),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_1_7_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_1_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_1_7_1  (
            .in0(N__14791),
            .in1(N__14776),
            .in2(N__14810),
            .in3(N__14761),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_1_7_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_1_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_1_7_2  (
            .in0(N__14746),
            .in1(N__14965),
            .in2(N__14999),
            .in3(N__14980),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_1_7_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_1_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_1_7_3  (
            .in0(N__14935),
            .in1(N__14950),
            .in2(N__14906),
            .in3(N__14920),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_1_7_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_1_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_1_7_4  (
            .in0(N__15190),
            .in1(N__14872),
            .in2(N__15176),
            .in3(N__14887),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_1_8_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_1_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_1_8_0  (
            .in0(N__14703),
            .in1(N__14634),
            .in2(N__14674),
            .in3(N__14723),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_1_8_1 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_1_8_1 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \COUNTER.counter_0_LC_1_8_1  (
            .in0(N__14724),
            .in1(_gnd_net_),
            .in2(N__26030),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33066),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_1_8_2 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_1_8_2 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_1_LC_1_8_2  (
            .in0(N__15042),
            .in1(N__26003),
            .in2(_gnd_net_),
            .in3(N__14725),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33066),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_1_8_3 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_1_8_3 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \COUNTER.counter_2_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__14690),
            .in2(N__26027),
            .in3(N__14704),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33066),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_1_8_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_1_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_1_8_4  (
            .in0(N__15157),
            .in1(N__15124),
            .in2(N__15143),
            .in3(N__15106),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_1_8_5 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_1_8_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_1_8_5 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \COUNTER.counter_3_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__14654),
            .in2(N__26028),
            .in3(N__14670),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33066),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_1_8_6 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_1_8_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_5_LC_1_8_6  (
            .in0(N__14603),
            .in1(N__26002),
            .in2(_gnd_net_),
            .in3(N__15067),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33066),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_1_8_7 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_1_8_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_1_8_7 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \COUNTER.counter_6_LC_1_8_7  (
            .in0(N__14591),
            .in1(_gnd_net_),
            .in2(N__26029),
            .in3(N__15091),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33066),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_1_9_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_1_9_0 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \POWERLED.func_state_1_LC_1_9_0  (
            .in0(N__23807),
            .in1(N__20545),
            .in2(N__21794),
            .in3(N__20531),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33067),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_1_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_1_9_1 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \POWERLED.func_state_0_LC_1_9_1  (
            .in0(N__21721),
            .in1(N__23808),
            .in2(N__21793),
            .in3(N__21707),
            .lcout(\POWERLED.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33067),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_1_9_2 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_1_9_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_1_9_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_4_LC_1_9_2  (
            .in0(N__14618),
            .in1(N__14638),
            .in2(_gnd_net_),
            .in3(N__26026),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33067),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_9_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_9_3  (
            .in0(N__17779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_1_9_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_1_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__14006),
            .in2(_gnd_net_),
            .in3(N__13976),
            .lcout(\POWERLED.mult1_un131_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17778),
            .lcout(\POWERLED.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_7  (
            .in0(N__13975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__18002),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__13719),
            .in2(N__15371),
            .in3(N__13742),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__13832),
            .in2(N__13724),
            .in3(N__13739),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__13823),
            .in2(N__13781),
            .in3(N__13736),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__13814),
            .in2(N__13780),
            .in3(N__13733),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_10_5  (
            .in0(N__17777),
            .in1(N__13723),
            .in2(N__13805),
            .in3(N__13730),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_10_6  (
            .in0(N__13793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13727),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13773),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__17977),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__15482),
            .in2(N__15402),
            .in3(N__13826),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__13751),
            .in2(N__15404),
            .in3(N__13817),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__13910),
            .in2(N__15439),
            .in3(N__13808),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__13901),
            .in2(N__15440),
            .in3(N__13796),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5  (
            .in0(N__13772),
            .in1(N__13892),
            .in2(N__15403),
            .in3(N__13787),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6  (
            .in0(N__13871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13784),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(\POWERLED.mult1_un138_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13754),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__17957),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__13934),
            .in2(N__15380),
            .in3(N__13745),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__13850),
            .in2(N__13859),
            .in3(N__13904),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__13838),
            .in2(N__13974),
            .in3(N__13895),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__14015),
            .in2(N__13973),
            .in3(N__13886),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_12_5  (
            .in0(N__15430),
            .in1(N__14002),
            .in2(N__13883),
            .in3(N__13865),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_12_6  (
            .in0(N__13988),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13862),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_1_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_1_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_1_12_7  (
            .in0(N__13849),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13961),
            .lcout(\POWERLED.mult1_un131_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__17936),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__15677),
            .in2(N__14067),
            .in3(N__13841),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__13928),
            .in2(N__14069),
            .in3(N__14018),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__13919),
            .in2(N__15670),
            .in3(N__14009),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__14102),
            .in2(N__15671),
            .in3(N__13991),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_13_5  (
            .in0(N__13960),
            .in1(N__14093),
            .in2(N__14068),
            .in3(N__13982),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_13_6  (
            .in0(N__14084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13979),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(\POWERLED.mult1_un124_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13937),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_1_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_1_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__17915),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_1_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__15602),
            .in2(N__15555),
            .in3(N__13922),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_1_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__14045),
            .in2(N__15557),
            .in3(N__13913),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_1_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__14036),
            .in2(N__15594),
            .in3(N__14096),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_1_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__14027),
            .in2(N__15595),
            .in3(N__14087),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_1_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_1_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_1_14_5  (
            .in0(N__15662),
            .in1(N__14159),
            .in2(N__15556),
            .in3(N__14078),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_1_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_1_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_1_14_6  (
            .in0(N__14150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14075),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(\POWERLED.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_1_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_1_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14072),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__17888),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__15827),
            .in2(N__14196),
            .in3(N__14039),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__14138),
            .in2(N__14198),
            .in3(N__14030),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__14129),
            .in2(N__15528),
            .in3(N__14021),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__14120),
            .in2(N__15529),
            .in3(N__14153),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_15_5  (
            .in0(N__15583),
            .in1(N__14111),
            .in2(N__14197),
            .in3(N__14144),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_15_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_15_6  (
            .in0(N__14213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14141),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_16_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__18161),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_16_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__15803),
            .in2(N__15820),
            .in3(N__14132),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_16_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__15816),
            .in2(N__15740),
            .in3(N__14123),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_16_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__15728),
            .in2(N__21891),
            .in3(N__14114),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_16_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__15719),
            .in2(N__21892),
            .in3(N__14105),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_16_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_16_5  (
            .in0(N__15527),
            .in1(N__15710),
            .in2(N__15821),
            .in3(N__14207),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_16_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_16_6  (
            .in0(N__15701),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14204),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(\POWERLED.mult1_un103_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_16_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_16_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14201),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI8CTK3_1_LC_2_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI8CTK3_1_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI8CTK3_1_LC_2_1_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \PCH_PWRGD.count_RNI8CTK3_1_LC_2_1_0  (
            .in0(N__17332),
            .in1(N__18635),
            .in2(N__14339),
            .in3(N__14165),
            .lcout(\PCH_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNI16MB1_LC_2_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNI16MB1_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNI16MB1_LC_2_1_1 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_c_RNI16MB1_LC_2_1_1  (
            .in0(N__17116),
            .in1(N__17333),
            .in2(N__17142),
            .in3(N__17483),
            .lcout(\PCH_PWRGD.count_rst_6 ),
            .ltout(\PCH_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIDC024_8_LC_2_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIDC024_8_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIDC024_8_LC_2_1_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNIDC024_8_LC_2_1_2  (
            .in0(_gnd_net_),
            .in1(N__15934),
            .in2(N__14174),
            .in3(N__18636),
            .lcout(\PCH_PWRGD.un2_count_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI3DJU_0_LC_2_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI3DJU_0_LC_2_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI3DJU_0_LC_2_1_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PCH_PWRGD.count_RNI3DJU_0_LC_2_1_3  (
            .in0(N__16976),
            .in1(N__17482),
            .in2(_gnd_net_),
            .in3(N__17331),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI7BTK3_0_LC_2_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI7BTK3_0_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI7BTK3_0_LC_2_1_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNI7BTK3_0_LC_2_1_4  (
            .in0(_gnd_net_),
            .in1(N__16010),
            .in2(N__14171),
            .in3(N__18634),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(\PCH_PWRGD.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI_1_LC_2_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI_1_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI_1_LC_2_1_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PCH_PWRGD.count_RNI_1_LC_2_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14168),
            .in3(N__17013),
            .lcout(\PCH_PWRGD.count_RNIZ0Z_1 ),
            .ltout(\PCH_PWRGD.count_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_1_LC_2_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_1_LC_2_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_1_LC_2_1_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \PCH_PWRGD.count_1_LC_2_1_6  (
            .in0(N__17334),
            .in1(_gnd_net_),
            .in2(N__14342),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32844),
            .ce(N__18701),
            .sr(N__18879));
    defparam \PCH_PWRGD.count_8_LC_2_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_8_LC_2_1_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_8_LC_2_1_7 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \PCH_PWRGD.count_8_LC_2_1_7  (
            .in0(N__17117),
            .in1(N__17335),
            .in2(N__17143),
            .in3(N__17484),
            .lcout(\PCH_PWRGD.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32844),
            .ce(N__18701),
            .sr(N__18879));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIB2J23_LC_2_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIB2J23_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIB2J23_LC_2_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIB2J23_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__20326),
            .in2(_gnd_net_),
            .in3(N__30585),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNI8U0P_0_LC_2_2_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNI8U0P_0_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNI8U0P_0_LC_2_2_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_RNI8U0P_0_LC_2_2_3  (
            .in0(N__14329),
            .in1(N__14317),
            .in2(N__14306),
            .in3(N__14290),
            .lcout(\DSW_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_2_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_2_2_4 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_LC_2_2_4  (
            .in0(N__14279),
            .in1(N__15898),
            .in2(N__31802),
            .in3(N__14495),
            .lcout(\PCH_PWRGD.delayed_vccin_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32927),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_2_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_2_2_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_2_2_5  (
            .in0(_gnd_net_),
            .in1(N__17306),
            .in2(_gnd_net_),
            .in3(N__32004),
            .lcout(\PCH_PWRGD.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_LC_2_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_LC_2_2_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI3DJU_0_LC_2_2_6  (
            .in0(N__14386),
            .in1(N__16120),
            .in2(N__14375),
            .in3(N__30584),
            .lcout(\PCH_PWRGD.curr_state_RNI3DJUZ0Z_0 ),
            .ltout(\PCH_PWRGD.curr_state_RNI3DJUZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIM8IJ2_LC_2_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIM8IJ2_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIM8IJ2_LC_2_2_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIM8IJ2_LC_2_2_7  (
            .in0(N__14494),
            .in1(N__14278),
            .in2(N__14270),
            .in3(N__31795),
            .lcout(PCH_PWRGD_delayed_vccin_ok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIEFB91_5_LC_2_3_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIEFB91_5_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIEFB91_5_LC_2_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_RNIEFB91_5_LC_2_3_0  (
            .in0(N__14267),
            .in1(N__14251),
            .in2(N__14240),
            .in3(N__14224),
            .lcout(\DSW_PWRGD.un4_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIQG1P_2_LC_2_3_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIQG1P_2_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIQG1P_2_LC_2_3_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIQG1P_2_LC_2_3_1  (
            .in0(N__14554),
            .in1(N__14542),
            .in2(N__14531),
            .in3(N__14512),
            .lcout(\DSW_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_LC_2_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16075),
            .lcout(\PCH_PWRGD.N_2126_i ),
            .ltout(\PCH_PWRGD.N_2126_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_3_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_LC_2_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14501),
            .in3(N__16119),
            .lcout(\PCH_PWRGD.N_381 ),
            .ltout(\PCH_PWRGD.N_381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_0_LC_2_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_0_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_0_LC_2_3_4 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI3DJU_0_0_LC_2_3_4  (
            .in0(N__30549),
            .in1(_gnd_net_),
            .in2(N__14498),
            .in3(N__14371),
            .lcout(\PCH_PWRGD.N_254_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_3_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_3_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_3_5  (
            .in0(N__14485),
            .in1(N__14473),
            .in2(N__14462),
            .in3(N__14446),
            .lcout(),
            .ltout(\DSW_PWRGD.un4_count_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_3_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_3_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIB8TE4_0_LC_2_3_6  (
            .in0(N__14435),
            .in1(N__14429),
            .in2(N__14423),
            .in3(N__14420),
            .lcout(\DSW_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_3_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_3_7  (
            .in0(N__14370),
            .in1(N__14393),
            .in2(_gnd_net_),
            .in3(N__30548),
            .lcout(\PCH_PWRGD.N_386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_4_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_4_0  (
            .in0(N__14387),
            .in1(N__14369),
            .in2(_gnd_net_),
            .in3(N__30583),
            .lcout(),
            .ltout(\PCH_PWRGD.N_255_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI7EHJ2_0_LC_2_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI7EHJ2_0_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI7EHJ2_0_LC_2_4_1 .LUT_INIT=16'b1100110100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI7EHJ2_0_LC_2_4_1  (
            .in0(N__16121),
            .in1(N__17330),
            .in2(N__14345),
            .in3(N__31793),
            .lcout(\PCH_PWRGD.curr_state_RNI7EHJ2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_2_5_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_2_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(N__15047),
            .in2(N__14732),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_5_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_2_5_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_2_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(N__14708),
            .in2(_gnd_net_),
            .in3(N__14678),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_2_5_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_2_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(N__14675),
            .in2(_gnd_net_),
            .in3(N__14645),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_2_5_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_2_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__14642),
            .in2(_gnd_net_),
            .in3(N__14606),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_2_5_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_2_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(N__15071),
            .in2(_gnd_net_),
            .in3(N__14594),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_2_5_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_2_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(N__15095),
            .in2(_gnd_net_),
            .in3(N__14579),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_2_5_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_2_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_2_5_6  (
            .in0(_gnd_net_),
            .in1(N__15019),
            .in2(_gnd_net_),
            .in3(N__14576),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__33086),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_2_5_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_2_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(N__14572),
            .in2(_gnd_net_),
            .in3(N__14558),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__33086),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_2_6_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_2_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__14857),
            .in2(_gnd_net_),
            .in3(N__14843),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_2_6_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_2_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__14840),
            .in2(_gnd_net_),
            .in3(N__14828),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_2_6_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_2_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(N__14825),
            .in2(_gnd_net_),
            .in3(N__14813),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_2_6_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_2_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__14809),
            .in2(_gnd_net_),
            .in3(N__14795),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_2_6_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_2_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__14792),
            .in2(_gnd_net_),
            .in3(N__14780),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_2_6_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_2_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_2_6_5  (
            .in0(_gnd_net_),
            .in1(N__14777),
            .in2(_gnd_net_),
            .in3(N__14765),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_2_6_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_2_6_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_2_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(N__14762),
            .in2(_gnd_net_),
            .in3(N__14750),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_2_6_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_2_6_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_2_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__14747),
            .in2(_gnd_net_),
            .in3(N__14735),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__32963),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_2_7_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_2_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__14998),
            .in2(_gnd_net_),
            .in3(N__14984),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_2_7_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_2_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__14981),
            .in2(_gnd_net_),
            .in3(N__14969),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_2_7_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_2_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__14966),
            .in2(_gnd_net_),
            .in3(N__14954),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_2_7_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_2_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__14951),
            .in2(_gnd_net_),
            .in3(N__14939),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_2_7_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_2_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__14936),
            .in2(_gnd_net_),
            .in3(N__14924),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_2_7_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_2_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__14921),
            .in2(_gnd_net_),
            .in3(N__14909),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_2_7_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_2_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__14905),
            .in2(_gnd_net_),
            .in3(N__14891),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_2_7_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_2_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__14888),
            .in2(_gnd_net_),
            .in3(N__14876),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__33069),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_2_8_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_2_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__14873),
            .in2(_gnd_net_),
            .in3(N__14861),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__33059),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_2_8_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_2_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__15191),
            .in2(_gnd_net_),
            .in3(N__15179),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__33059),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_2_8_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_2_8_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_2_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__15175),
            .in2(_gnd_net_),
            .in3(N__15161),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__33059),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_2_8_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_2_8_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_2_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(N__15158),
            .in2(_gnd_net_),
            .in3(N__15146),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__33059),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_2_8_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_2_8_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_2_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_29_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__15142),
            .in2(_gnd_net_),
            .in3(N__15128),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__33059),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_2_8_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_2_8_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_2_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_30_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__15125),
            .in2(_gnd_net_),
            .in3(N__15113),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__33059),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_2_8_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_2_8_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_2_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__15107),
            .in2(_gnd_net_),
            .in3(N__15110),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33059),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_2_8_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_2_8_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_2_8_7  (
            .in0(N__15087),
            .in1(N__15063),
            .in2(N__15043),
            .in3(N__15020),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_2_9_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_2_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__15005),
            .in2(N__16430),
            .in3(N__25100),
            .lcout(\POWERLED.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_2_9_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__15290),
            .in2(N__15281),
            .in3(N__25148),
            .lcout(\POWERLED.N_4527_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_0 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_2_9_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_2_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__15272),
            .in2(N__16469),
            .in3(N__19334),
            .lcout(\POWERLED.N_4528_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_1 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_2_9_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_2_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__15254),
            .in2(N__15266),
            .in3(N__19295),
            .lcout(\POWERLED.N_4529_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_2 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_2_9_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_2_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__15233),
            .in2(N__15248),
            .in3(N__19256),
            .lcout(\POWERLED.N_4530_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_3 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_2_9_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_2_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_2_9_5  (
            .in0(N__20741),
            .in1(N__15227),
            .in2(N__15476),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4531_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_4 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_2_9_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_2_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_2_9_6  (
            .in0(N__20651),
            .in1(N__15209),
            .in2(N__15221),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4532_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_5 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_2_9_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_2_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__15203),
            .in2(N__15641),
            .in3(N__19553),
            .lcout(\POWERLED.N_4533_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_6 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_2_10_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_2_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_2_10_0  (
            .in0(N__19514),
            .in1(N__15197),
            .in2(N__15692),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4534_i ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_2_10_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_2_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_2_10_1  (
            .in0(N__19595),
            .in1(N__15347),
            .in2(N__15494),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4535_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_8 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_2_10_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_2_10_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_2_10_2  (
            .in0(N__19469),
            .in1(N__15341),
            .in2(N__21851),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4536_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_9 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_2_10_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_2_10_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_2_10_3  (
            .in0(N__19418),
            .in1(N__15335),
            .in2(N__15461),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4537_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_10 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_2_10_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_2_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_2_10_4  (
            .in0(N__21998),
            .in1(N__15329),
            .in2(N__15626),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4538_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_11 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_2_10_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_2_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__15356),
            .in2(N__15323),
            .in3(N__20486),
            .lcout(\POWERLED.N_4539_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_12 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_2_10_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_2_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_2_10_6  (
            .in0(N__20696),
            .in1(N__15782),
            .in2(N__15314),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4540_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_13 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_2_10_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_2_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_2_10_7  (
            .in0(N__19655),
            .in1(N__15614),
            .in2(N__15305),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4541_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_14 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_2_11_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_2_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15293),
            .lcout(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_11_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_11_1  (
            .in0(N__16526),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15533),
            .lcout(\POWERLED.un85_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_11_5  (
            .in0(N__17953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15438),
            .lcout(\POWERLED.un85_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16826),
            .lcout(\POWERLED.un85_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_SUSn_RNIN4K9_LC_2_12_1.C_ON=1'b0;
    defparam SLP_SUSn_RNIN4K9_LC_2_12_1.SEQ_MODE=4'b0000;
    defparam SLP_SUSn_RNIN4K9_LC_2_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 SLP_SUSn_RNIN4K9_LC_2_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16256),
            .lcout(v33a_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_2_12_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_2_12_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_2_12_2  (
            .in0(N__15431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_12_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_12_3  (
            .in0(N__17935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_12_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_12_4  (
            .in0(N__17981),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20111),
            .lcout(\POWERLED.un85_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_13_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15596),
            .lcout(\POWERLED.un85_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17914),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_LC_2_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_LC_2_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_15_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23379),
            .lcout(\POWERLED.N_2215_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15669),
            .lcout(\POWERLED.un85_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18395),
            .lcout(\POWERLED.un85_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_14_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18314),
            .lcout(\POWERLED.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_14_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18104),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_2_14_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_2_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17884),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15590),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_14_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__20204),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_14_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_14_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_2_14_7  (
            .in0(N__15773),
            .in1(N__29276),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__18124),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__15749),
            .in2(N__15844),
            .in3(N__15731),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__15840),
            .in2(N__16658),
            .in3(N__15722),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__16815),
            .in2(N__16643),
            .in3(N__15713),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__16865),
            .in2(N__16822),
            .in3(N__15704),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_15_5  (
            .in0(N__21880),
            .in1(N__16853),
            .in2(N__15845),
            .in3(N__15695),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__16841),
            .in2(_gnd_net_),
            .in3(N__15848),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16814),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_16_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18160),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_6  (
            .in0(N__21881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_2_16_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_2_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18128),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_4_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_4_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_4_1_0  (
            .in0(N__15788),
            .in1(N__16046),
            .in2(_gnd_net_),
            .in3(N__31959),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_1 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_1  (
            .in0(N__15910),
            .in1(N__16117),
            .in2(N__15797),
            .in3(N__15953),
            .lcout(),
            .ltout(\PCH_PWRGD.m4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI09KEQ_0_LC_4_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI09KEQ_0_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI09KEQ_0_LC_4_1_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNI09KEQ_0_LC_4_1_2  (
            .in0(_gnd_net_),
            .in1(N__15887),
            .in2(N__15794),
            .in3(N__31960),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_3 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_4_1_3  (
            .in0(N__16068),
            .in1(N__17481),
            .in2(N__15791),
            .in3(N__17393),
            .lcout(\PCH_PWRGD.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32843),
            .ce(N__31764),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIFF124_9_LC_4_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIFF124_9_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIFF124_9_LC_4_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNIFF124_9_LC_4_1_5  (
            .in0(N__17030),
            .in1(N__17234),
            .in2(_gnd_net_),
            .in3(N__18692),
            .lcout(\PCH_PWRGD.countZ0Z_9 ),
            .ltout(\PCH_PWRGD.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIDC024_0_8_LC_4_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIDC024_0_8_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIDC024_0_8_LC_4_1_6 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \PCH_PWRGD.count_RNIDC024_0_8_LC_4_1_6  (
            .in0(N__18693),
            .in1(N__15938),
            .in2(N__15923),
            .in3(N__15920),
            .lcout(\PCH_PWRGD.un12_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_7 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_7 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_4_1_7  (
            .in0(N__16067),
            .in1(N__16116),
            .in2(N__15911),
            .in3(N__15952),
            .lcout(\PCH_PWRGD.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32843),
            .ce(N__31764),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI3TQ14_0_3_LC_4_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI3TQ14_0_3_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI3TQ14_0_3_LC_4_2_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \PCH_PWRGD.count_RNI3TQ14_0_3_LC_4_2_0  (
            .in0(N__15881),
            .in1(N__15869),
            .in2(N__18713),
            .in3(N__16909),
            .lcout(\PCH_PWRGD.un12_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNISRGB1_LC_4_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNISRGB1_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNISRGB1_LC_4_2_1 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_c_RNISRGB1_LC_4_2_1  (
            .in0(N__16927),
            .in1(N__16943),
            .in2(N__17478),
            .in3(N__17380),
            .lcout(\PCH_PWRGD.count_rst_11 ),
            .ltout(\PCH_PWRGD.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI3TQ14_3_LC_4_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI3TQ14_3_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI3TQ14_3_LC_4_2_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \PCH_PWRGD.count_RNI3TQ14_3_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(N__18680),
            .in2(N__15875),
            .in3(N__15868),
            .lcout(\PCH_PWRGD.un2_count_1_axb_3 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_3_LC_4_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_3_LC_4_2_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_3_LC_4_2_3 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \PCH_PWRGD.count_3_LC_4_2_3  (
            .in0(N__17448),
            .in1(N__16931),
            .in2(N__15872),
            .in3(N__17384),
            .lcout(\PCH_PWRGD.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32769),
            .ce(N__18717),
            .sr(N__18913));
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNITTHB1_LC_4_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNITTHB1_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNITTHB1_LC_4_2_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_c_RNITTHB1_LC_4_2_4  (
            .in0(N__17381),
            .in1(N__17446),
            .in2(N__16913),
            .in3(N__16891),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI50S14_4_LC_4_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI50S14_4_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI50S14_4_LC_4_2_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNI50S14_4_LC_4_2_5  (
            .in0(N__18681),
            .in1(_gnd_net_),
            .in2(N__15860),
            .in3(N__15854),
            .lcout(\PCH_PWRGD.countZ0Z_4 ),
            .ltout(\PCH_PWRGD.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_4_LC_4_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_4_LC_4_2_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_4_LC_4_2_6 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.count_4_LC_4_2_6  (
            .in0(N__17382),
            .in1(N__17449),
            .in2(N__15857),
            .in3(N__16892),
            .lcout(\PCH_PWRGD.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32769),
            .ce(N__18717),
            .sr(N__18913));
    defparam \PCH_PWRGD.count_0_LC_4_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_LC_4_2_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_0_LC_4_2_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \PCH_PWRGD.count_0_LC_4_2_7  (
            .in0(N__17447),
            .in1(N__16990),
            .in2(_gnd_net_),
            .in3(N__17383),
            .lcout(\PCH_PWRGD.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32769),
            .ce(N__18717),
            .sr(N__18913));
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIBHA61_LC_4_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIBHA61_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIBHA61_LC_4_3_0 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_c_RNIBHA61_LC_4_3_0  (
            .in0(N__17377),
            .in1(N__17080),
            .in2(N__17480),
            .in3(N__17093),
            .lcout(\PCH_PWRGD.count_rst_3 ),
            .ltout(\PCH_PWRGD.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI14454_11_LC_4_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI14454_11_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI14454_11_LC_4_3_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \PCH_PWRGD.count_RNI14454_11_LC_4_3_1  (
            .in0(N__15982),
            .in1(_gnd_net_),
            .in2(N__15998),
            .in3(N__18702),
            .lcout(\PCH_PWRGD.un2_count_1_axb_11 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_11_LC_4_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_11_LC_4_3_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_11_LC_4_3_2 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.count_11_LC_4_3_2  (
            .in0(N__17378),
            .in1(N__17459),
            .in2(N__15995),
            .in3(N__17081),
            .lcout(\PCH_PWRGD.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32985),
            .ce(N__18719),
            .sr(N__18937));
    defparam \PCH_PWRGD.count_RNI14454_0_11_LC_4_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI14454_0_11_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI14454_0_11_LC_4_3_3 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \PCH_PWRGD.count_RNI14454_0_11_LC_4_3_3  (
            .in0(N__15992),
            .in1(N__17021),
            .in2(N__15986),
            .in3(N__18703),
            .lcout(),
            .ltout(\PCH_PWRGD.un12_clk_100khz_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOGSAG_3_LC_4_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOGSAG_3_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOGSAG_3_LC_4_3_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIOGSAG_3_LC_4_3_4  (
            .in0(N__15974),
            .in1(N__16760),
            .in2(N__15968),
            .in3(N__15965),
            .lcout(),
            .ltout(\PCH_PWRGD.un12_clk_100khz_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIVBLSO_2_LC_4_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIVBLSO_2_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIVBLSO_2_LC_4_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIVBLSO_2_LC_4_3_5  (
            .in0(N__18797),
            .in1(N__16034),
            .in2(N__15956),
            .in3(N__18521),
            .lcout(\PCH_PWRGD.N_1_i ),
            .ltout(\PCH_PWRGD.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIVBLSO_0_2_LC_4_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIVBLSO_0_2_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIVBLSO_0_2_LC_4_3_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.count_RNIVBLSO_0_2_LC_4_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15941),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2 ),
            .ltout(\PCH_PWRGD.count_RNIVBLSO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_3_7 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_3_7  (
            .in0(N__16118),
            .in1(N__16079),
            .in2(N__16049),
            .in3(N__17379),
            .lcout(\PCH_PWRGD.curr_state_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_14_LC_4_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_14_LC_4_4_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_14_LC_4_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_14_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17527),
            .lcout(\PCH_PWRGD.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32819),
            .ce(N__18666),
            .sr(N__18927));
    defparam \PCH_PWRGD.count_RNI9G854_15_LC_4_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI9G854_15_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI9G854_15_LC_4_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNI9G854_15_LC_4_4_1  (
            .in0(N__16016),
            .in1(N__17500),
            .in2(_gnd_net_),
            .in3(N__18665),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(\PCH_PWRGD.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI_15_LC_4_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI_15_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI_15_LC_4_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_RNI_15_LC_4_4_2  (
            .in0(N__16989),
            .in1(N__17540),
            .in2(N__16037),
            .in3(N__17066),
            .lcout(\PCH_PWRGD.un12_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNILIKA4_14_LC_4_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNILIKA4_14_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNILIKA4_14_LC_4_4_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \PCH_PWRGD.count_RNILIKA4_14_LC_4_4_3  (
            .in0(N__16028),
            .in1(_gnd_net_),
            .in2(N__17528),
            .in3(N__18664),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI5A654_13_LC_4_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI5A654_13_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI5A654_13_LC_4_4_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNI5A654_13_LC_4_4_5  (
            .in0(N__16022),
            .in1(N__18663),
            .in2(_gnd_net_),
            .in3(N__17053),
            .lcout(\PCH_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_13_LC_4_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_13_LC_4_4_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_13_LC_4_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_13_LC_4_4_6  (
            .in0(N__17054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32819),
            .ce(N__18666),
            .sr(N__18927));
    defparam \PCH_PWRGD.count_15_LC_4_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_15_LC_4_4_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_15_LC_4_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_15_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17501),
            .lcout(\PCH_PWRGD.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32819),
            .ce(N__18666),
            .sr(N__18927));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_4_5_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_4_5_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_LC_4_5_0  (
            .in0(N__30415),
            .in1(N__17642),
            .in2(_gnd_net_),
            .in3(N__16185),
            .lcout(RSMRST_PWRGD_RSMRSTn_2_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33085),
            .ce(N__29415),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_LC_4_5_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_LC_4_5_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_0_LC_4_5_2  (
            .in0(N__30418),
            .in1(N__17640),
            .in2(_gnd_net_),
            .in3(N__16182),
            .lcout(\RSMRST_PWRGD.N_256_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_5_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_5_3 .LUT_INIT=16'b0000011100000010;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_4_5_3  (
            .in0(N__16184),
            .in1(N__17222),
            .in2(N__17650),
            .in3(N__30416),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33085),
            .ce(N__29415),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_o2_LC_4_5_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_o2_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_o2_LC_4_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_o2_LC_4_5_4  (
            .in0(N__30417),
            .in1(N__17221),
            .in2(_gnd_net_),
            .in3(N__16183),
            .lcout(N_187),
            .ltout(N_187_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_5_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_5_5 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_4_5_5  (
            .in0(N__17646),
            .in1(_gnd_net_),
            .in2(N__16310),
            .in3(N__16187),
            .lcout(RSMRST_PWRGD_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33085),
            .ce(N__29415),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_5_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_5_6  (
            .in0(N__16296),
            .in1(N__16265),
            .in2(N__16255),
            .in3(N__16219),
            .lcout(rsmrst_pwrgd_signal),
            .ltout(rsmrst_pwrgd_signal_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_4_5_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_4_5_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_LC_4_5_7  (
            .in0(N__17641),
            .in1(_gnd_net_),
            .in2(N__16190),
            .in3(N__16186),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33085),
            .ce(N__29415),
            .sr(_gnd_net_));
    defparam \POWERLED.count_4_LC_4_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_4_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_4_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_4_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19229),
            .lcout(\POWERLED.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32964),
            .ce(N__31765),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_4_7_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_4_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16163),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_4_7_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_4_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_4_7_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_4_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16133),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_4_7_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_4_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16400),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_4_7_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_4_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16388),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_4_7_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_4_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16376),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_4_7_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_4_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__16364),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_4_7_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_4_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16355),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(COUNTER_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_8_0.C_ON=1'b0;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_8_0.SEQ_MODE=4'b0000;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16340),
            .lcout(COUNTER_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.slp_s3n_signal_i_LC_4_8_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.slp_s3n_signal_i_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.slp_s3n_signal_i_LC_4_8_7 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \PCH_PWRGD.slp_s3n_signal_i_LC_4_8_7  (
            .in0(N__22387),
            .in1(N__22489),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__26933),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__16418),
            .in2(N__16450),
            .in3(N__16514),
            .lcout(G_2121),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__16446),
            .in2(N__16412),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__16515),
            .in2(N__16568),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__16556),
            .in2(N__16522),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__16547),
            .in2(N__16451),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_9_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_9_6  (
            .in0(N__16538),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16433),
            .lcout(\POWERLED.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26490),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_4_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_4_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__26491),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_4_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_4_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__16479),
            .in2(N__16493),
            .in3(N__16403),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_4_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_4_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__17840),
            .in2(N__16484),
            .in3(N__16559),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_4_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_4_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__18023),
            .in2(N__17822),
            .in3(N__16550),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_4_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_4_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__17798),
            .in2(N__18029),
            .in3(N__16541),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_4_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_4_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_4_10_5  (
            .in0(N__16513),
            .in1(N__16483),
            .in2(N__17747),
            .in3(N__16532),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_4_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_4_10_6  (
            .in0(N__17699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16529),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26266),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_4_11_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_4_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_4_11_0  (
            .in0(N__18028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_4_11_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_4_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18027),
            .lcout(\POWERLED.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_4_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_4_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17992),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19828),
            .lcout(\POWERLED.mult1_un47_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18061),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_4_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_4_12_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_15_LC_4_12_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.dutycycle_15_LC_4_12_0  (
            .in0(N__19903),
            .in1(N__25817),
            .in2(N__19928),
            .in3(N__21068),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33113),
            .ce(),
            .sr(N__22884));
    defparam \POWERLED.dutycycle_12_LC_4_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_12_LC_4_12_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_12_LC_4_12_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.dutycycle_12_LC_4_12_2  (
            .in0(N__23492),
            .in1(N__25816),
            .in2(N__23512),
            .in3(N__23642),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33113),
            .ce(),
            .sr(N__22884));
    defparam \POWERLED.dutycycle_RNI_2_14_LC_4_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_4_12_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \POWERLED.dutycycle_RNI_2_14_LC_4_12_4  (
            .in0(N__19753),
            .in1(N__23470),
            .in2(N__21215),
            .in3(N__23045),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_9_LC_4_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_9_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_9_LC_4_12_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_9_LC_4_12_5  (
            .in0(N__24280),
            .in1(N__23264),
            .in2(N__16586),
            .in3(N__22640),
            .lcout(\POWERLED.N_336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_11_LC_4_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_4_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_11_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(N__23469),
            .in2(_gnd_net_),
            .in3(N__24279),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_46_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_14_LC_4_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_4_12_7 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_14_LC_4_12_7  (
            .in0(N__22649),
            .in1(N__21211),
            .in2(N__16583),
            .in3(N__20264),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18062),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__16580),
            .in2(_gnd_net_),
            .in3(N__16571),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__20051),
            .in2(N__18197),
            .in3(N__16628),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__27461),
            .in2(N__20027),
            .in3(N__16625),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__27469),
            .in2(N__20003),
            .in3(N__16622),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_13_5  (
            .in0(N__16725),
            .in1(N__26108),
            .in2(N__26081),
            .in3(N__16619),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_13_6 .LUT_INIT=16'b0011000011001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__25411),
            .in2(N__25432),
            .in3(N__16616),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(\POWERLED.mult1_un54_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16613),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__18188),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__16610),
            .in2(N__16693),
            .in3(N__16601),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__16689),
            .in2(N__16598),
            .in3(N__16589),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__16739),
            .in2(N__16730),
            .in3(N__16733),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__16729),
            .in2(N__16712),
            .in3(N__16703),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_14_5  (
            .in0(N__18305),
            .in1(N__16700),
            .in2(N__16694),
            .in3(N__16676),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16673),
            .in3(N__16664),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(\POWERLED.mult1_un61_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16661),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__18100),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__18209),
            .in2(N__16789),
            .in3(N__16646),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__16785),
            .in2(N__18452),
            .in3(N__16631),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__18383),
            .in2(N__18440),
            .in3(N__16856),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__18428),
            .in2(N__18391),
            .in3(N__16844),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_15_5  (
            .in0(N__16813),
            .in1(N__18419),
            .in2(N__16790),
            .in3(N__16832),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18410),
            .in3(N__16829),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18382),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI73T14_5_LC_5_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI73T14_5_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI73T14_5_LC_5_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNI73T14_5_LC_5_1_0  (
            .in0(N__16768),
            .in1(N__16747),
            .in2(_gnd_net_),
            .in3(N__18690),
            .lcout(\PCH_PWRGD.un2_count_1_axb_5 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_5_LC_5_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_5_LC_5_1_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_5_LC_5_1_1 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \PCH_PWRGD.count_5_LC_5_1_1  (
            .in0(N__17487),
            .in1(N__17192),
            .in2(N__16772),
            .in3(N__17388),
            .lcout(\PCH_PWRGD.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32693),
            .ce(N__18697),
            .sr(N__18938));
    defparam \PCH_PWRGD.count_RNI73T14_0_5_LC_5_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI73T14_0_5_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI73T14_0_5_LC_5_1_2 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \PCH_PWRGD.count_RNI73T14_0_5_LC_5_1_2  (
            .in0(N__16769),
            .in1(N__17176),
            .in2(N__18715),
            .in3(N__16748),
            .lcout(\PCH_PWRGD.un12_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIUVIB1_LC_5_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIUVIB1_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIUVIB1_LC_5_1_3 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_c_RNIUVIB1_LC_5_1_3  (
            .in0(N__17485),
            .in1(N__17191),
            .in2(N__16880),
            .in3(N__17385),
            .lcout(\PCH_PWRGD.count_rst_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNI04LB1_LC_5_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNI04LB1_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNI04LB1_LC_5_1_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_c_RNI04LB1_LC_5_1_4  (
            .in0(N__17386),
            .in1(N__17486),
            .in2(N__17162),
            .in3(N__17177),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIB9V14_7_LC_5_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIB9V14_7_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIB9V14_7_LC_5_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIB9V14_7_LC_5_1_5  (
            .in0(N__18691),
            .in1(_gnd_net_),
            .in2(N__17042),
            .in3(N__17036),
            .lcout(\PCH_PWRGD.countZ0Z_7 ),
            .ltout(\PCH_PWRGD.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_7_LC_5_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_7_LC_5_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_7_LC_5_1_6 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.count_7_LC_5_1_6  (
            .in0(N__17387),
            .in1(N__17488),
            .in2(N__17039),
            .in3(N__17161),
            .lcout(\PCH_PWRGD.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32693),
            .ce(N__18697),
            .sr(N__18938));
    defparam \PCH_PWRGD.count_9_LC_5_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_9_LC_5_1_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_9_LC_5_1_7 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \PCH_PWRGD.count_9_LC_5_1_7  (
            .in0(N__17392),
            .in1(N__17249),
            .in2(N__17492),
            .in3(N__17265),
            .lcout(\PCH_PWRGD.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32693),
            .ce(N__18697),
            .sr(N__18938));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_5_2_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_5_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__17020),
            .in2(N__16991),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSC_LC_5_2_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSC_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSC_LC_5_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSC_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__18944),
            .in2(_gnd_net_),
            .in3(N__16946),
            .lcout(\PCH_PWRGD.un2_count_1_cry_1_c_RNIOCSCZ0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_5_2_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_5_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__16942),
            .in2(_gnd_net_),
            .in3(N__16916),
            .lcout(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_5_2_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_5_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__16908),
            .in2(_gnd_net_),
            .in3(N__16883),
            .lcout(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_5_2_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_5_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__16876),
            .in2(_gnd_net_),
            .in3(N__17183),
            .lcout(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNIV1KB1_LC_5_2_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNIV1KB1_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNIV1KB1_LC_5_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_5_c_RNIV1KB1_LC_5_2_5  (
            .in0(N__17389),
            .in1(N__18814),
            .in2(_gnd_net_),
            .in3(N__17180),
            .lcout(\PCH_PWRGD.count_rst_8 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_5_2_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_5_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__17175),
            .in2(_gnd_net_),
            .in3(N__17147),
            .lcout(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_5_2_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_5_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__17144),
            .in2(_gnd_net_),
            .in3(N__17102),
            .lcout(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_7 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_5_3_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_5_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__17266),
            .in2(_gnd_net_),
            .in3(N__17099),
            .lcout(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNI3AOB1_LC_5_3_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNI3AOB1_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNI3AOB1_LC_5_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_9_c_RNI3AOB1_LC_5_3_1  (
            .in0(N__17394),
            .in1(N__17660),
            .in2(_gnd_net_),
            .in3(N__17096),
            .lcout(\PCH_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_5_3_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_5_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(N__17092),
            .in2(_gnd_net_),
            .in3(N__17072),
            .lcout(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNICJB61_LC_5_3_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNICJB61_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNICJB61_LC_5_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_11_c_RNICJB61_LC_5_3_3  (
            .in0(N__17395),
            .in1(N__18764),
            .in2(_gnd_net_),
            .in3(N__17069),
            .lcout(\PCH_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIDLC61_LC_5_3_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIDLC61_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIDLC61_LC_5_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_12_c_RNIDLC61_LC_5_3_4  (
            .in0(N__17391),
            .in1(N__17065),
            .in2(_gnd_net_),
            .in3(N__17045),
            .lcout(\PCH_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNISSQB1_LC_5_3_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNISSQB1_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNISSQB1_LC_5_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_13_c_RNISSQB1_LC_5_3_5  (
            .in0(N__18926),
            .in1(N__17539),
            .in2(_gnd_net_),
            .in3(N__17516),
            .lcout(\PCH_PWRGD.count_rst_0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNIFPE61_LC_5_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNIFPE61_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNIFPE61_LC_5_3_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_14_c_RNIFPE61_LC_5_3_6  (
            .in0(N__17513),
            .in1(N__17396),
            .in2(_gnd_net_),
            .in3(N__17504),
            .lcout(\PCH_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNI28NB1_LC_5_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNI28NB1_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNI28NB1_LC_5_3_7 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_c_RNI28NB1_LC_5_3_7  (
            .in0(N__17479),
            .in1(N__17390),
            .in2(N__17270),
            .in3(N__17245),
            .lcout(\PCH_PWRGD.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI9RLK1_3_LC_5_4_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI9RLK1_3_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI9RLK1_3_LC_5_4_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_RNI9RLK1_3_LC_5_4_0  (
            .in0(N__19021),
            .in1(N__19036),
            .in2(N__19070),
            .in3(N__19006),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_5_4_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_5_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIR8OP4_10_LC_5_4_1  (
            .in0(N__17198),
            .in1(N__17204),
            .in2(N__17225),
            .in3(N__17210),
            .lcout(\RSMRST_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_5_4_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_5_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_5_4_2  (
            .in0(N__19156),
            .in1(N__19138),
            .in2(N__19193),
            .in3(N__19207),
            .lcout(\RSMRST_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIBFU91_13_LC_5_4_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIBFU91_13_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIBFU91_13_LC_5_4_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \RSMRST_PWRGD.count_RNIBFU91_13_LC_5_4_3  (
            .in0(N__19084),
            .in1(N__18487),
            .in2(N__19175),
            .in3(N__18475),
            .lcout(\RSMRST_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIQUU91_10_LC_5_4_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIQUU91_10_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIQUU91_10_LC_5_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIQUU91_10_LC_5_4_4  (
            .in0(N__19051),
            .in1(N__18973),
            .in2(N__18992),
            .in3(N__18958),
            .lcout(\RSMRST_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_5_5_0 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_5_5_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.curr_state_RNI1KAM_0_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(N__31800),
            .in2(_gnd_net_),
            .in3(N__25213),
            .lcout(\POWERLED.g0_i_o3_0 ),
            .ltout(\POWERLED.g0_i_o3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_5_5_1 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_5_5_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.pwm_out_LC_5_5_1 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \POWERLED.pwm_out_LC_5_5_1  (
            .in0(N__17596),
            .in1(N__25248),
            .in2(N__17600),
            .in3(N__19342),
            .lcout(\POWERLED.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32900),
            .ce(),
            .sr(N__19373));
    defparam \POWERLED.pwm_out_RNIB7P12_LC_5_5_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNIB7P12_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNIB7P12_LC_5_5_2 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \POWERLED.pwm_out_RNIB7P12_LC_5_5_2  (
            .in0(N__25249),
            .in1(N__17597),
            .in2(N__19346),
            .in3(N__17588),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_5_5_3 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_5_5_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_5_5_3  (
            .in0(N__25214),
            .in1(N__25182),
            .in2(_gnd_net_),
            .in3(N__25247),
            .lcout(),
            .ltout(\POWERLED.curr_state_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_5_5_4 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_5_5_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.curr_state_RNI2P6L_0_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__25163),
            .in2(N__17564),
            .in3(N__31967),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(\POWERLED.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_5_5_5 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_5_5_5 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \POWERLED.curr_state_RNIE5D5_0_LC_5_5_5  (
            .in0(N__31968),
            .in1(_gnd_net_),
            .in2(N__17561),
            .in3(N__25181),
            .lcout(\POWERLED.count_0_sqmuxa_i ),
            .ltout(\POWERLED.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_0_LC_5_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_0_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_0_LC_5_5_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_RNI_0_LC_5_5_6  (
            .in0(N__25084),
            .in1(_gnd_net_),
            .in2(N__17558),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.count_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIFAFE_0_LC_5_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIFAFE_0_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIFAFE_0_LC_5_5_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIFAFE_0_LC_5_5_7  (
            .in0(N__31969),
            .in1(_gnd_net_),
            .in2(N__17555),
            .in3(N__24965),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI96U14_6_LC_5_6_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI96U14_6_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI96U14_6_LC_5_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNI96U14_6_LC_5_6_0  (
            .in0(N__18688),
            .in1(N__17666),
            .in2(_gnd_net_),
            .in3(N__17551),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_6_LC_5_6_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_6_LC_5_6_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_6_LC_5_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_6_LC_5_6_1  (
            .in0(N__17552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32989),
            .ce(N__18718),
            .sr(N__18928));
    defparam \PCH_PWRGD.count_RNIORHA4_10_LC_5_6_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIORHA4_10_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIORHA4_10_LC_5_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNIORHA4_10_LC_5_6_2  (
            .in0(N__18689),
            .in1(N__18736),
            .in2(_gnd_net_),
            .in3(N__18757),
            .lcout(\PCH_PWRGD.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_10_LC_5_6_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_10_LC_5_6_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_10_LC_5_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_10_LC_5_6_3  (
            .in0(N__18758),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32989),
            .ce(N__18718),
            .sr(N__18928));
    defparam \POWERLED.G_11_LC_5_6_4 .C_ON=1'b0;
    defparam \POWERLED.G_11_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_11_LC_5_6_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \POWERLED.G_11_LC_5_6_4  (
            .in0(N__17651),
            .in1(N__17621),
            .in2(_gnd_net_),
            .in3(N__29539),
            .lcout(G_11),
            .ltout(G_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_6_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_6_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_6_5  (
            .in0(N__29540),
            .in1(_gnd_net_),
            .in2(N__17615),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.N_27_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_209_i_LC_5_6_6 .C_ON=1'b0;
    defparam \POWERLED.N_209_i_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_209_i_LC_5_6_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.N_209_i_LC_5_6_6  (
            .in0(N__27890),
            .in1(N__28056),
            .in2(_gnd_net_),
            .in3(N__31993),
            .lcout(\POWERLED.N_209_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI0LHN_4_LC_5_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI0LHN_4_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI0LHN_4_LC_5_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI0LHN_4_LC_5_6_7  (
            .in0(N__31992),
            .in1(N__17612),
            .in2(_gnd_net_),
            .in3(N__19222),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIJKSP_10_LC_5_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIJKSP_10_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIJKSP_10_LC_5_7_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \POWERLED.count_RNIJKSP_10_LC_5_7_0  (
            .in0(N__17858),
            .in1(_gnd_net_),
            .in2(N__19438),
            .in3(N__31997),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNISEFN_2_LC_5_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNISEFN_2_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNISEFN_2_LC_5_7_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNISEFN_2_LC_5_7_2  (
            .in0(N__17606),
            .in1(N__31994),
            .in2(_gnd_net_),
            .in3(N__19306),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_5_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_2_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_5_7_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_2_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19310),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33016),
            .ce(N__31768),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNISF4O_11_LC_5_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNISF4O_11_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNISF4O_11_LC_5_7_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \POWERLED.count_RNISF4O_11_LC_5_7_4  (
            .in0(N__17690),
            .in1(_gnd_net_),
            .in2(N__19394),
            .in3(N__31996),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_11_LC_5_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_11_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_5_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_11_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19393),
            .lcout(\POWERLED.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33016),
            .ce(N__31768),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUHGN_3_LC_5_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUHGN_3_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUHGN_3_LC_5_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIUHGN_3_LC_5_7_6  (
            .in0(N__17684),
            .in1(N__31995),
            .in2(_gnd_net_),
            .in3(N__19267),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_3_LC_5_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_3_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_5_7_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_3_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19271),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33016),
            .ce(N__31768),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI4S8O_15_LC_5_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI4S8O_15_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI4S8O_15_LC_5_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI4S8O_15_LC_5_8_0  (
            .in0(N__17678),
            .in1(N__31989),
            .in2(_gnd_net_),
            .in3(N__19621),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_15_LC_5_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_15_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_15_LC_5_8_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_15_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19625),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33070),
            .ce(N__31770),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI6UKN_7_LC_5_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI6UKN_7_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI6UKN_7_LC_5_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI6UKN_7_LC_5_8_2  (
            .in0(N__17672),
            .in1(N__31990),
            .in2(_gnd_net_),
            .in3(N__19525),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_7_LC_5_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_7_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_5_8_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_7_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19529),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33070),
            .ce(N__31770),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI81MN_8_LC_5_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI81MN_8_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI81MN_8_LC_5_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI81MN_8_LC_5_8_4  (
            .in0(N__17864),
            .in1(N__31991),
            .in2(_gnd_net_),
            .in3(N__19483),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_8_LC_5_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_8_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_5_8_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_8_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19487),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33070),
            .ce(N__31770),
            .sr(_gnd_net_));
    defparam \POWERLED.count_9_LC_5_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_9_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_5_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_9_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19607),
            .lcout(\POWERLED.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33070),
            .ce(N__31770),
            .sr(_gnd_net_));
    defparam \POWERLED.count_10_LC_5_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_10_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_5_9_6 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_10_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19439),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33078),
            .ce(N__31769),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_LC_5_10_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_2_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_LC_5_10_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26241),
            .in3(N__26739),
            .lcout(\POWERLED.N_337 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__17727),
            .in2(N__17849),
            .in3(N__17834),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__17831),
            .in2(N__17732),
            .in3(N__17810),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__17807),
            .in2(N__17789),
            .in3(N__17792),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__17788),
            .in2(N__17759),
            .in3(N__17735),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_10_5  (
            .in0(N__18022),
            .in1(N__17731),
            .in2(N__17711),
            .in3(N__17693),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_10_6  (
            .in0(N__18041),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18032),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_LC_5_10_7 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_fast_LC_5_10_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.tmp_0_fast_LC_5_10_7  (
            .in0(N__26000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22072),
            .lcout(SUSWARN_N_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33071),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_3_LC_5_11_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_5_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_3_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__26695),
            .in2(N__26942),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_5_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__26937),
            .in2(N__20951),
            .in3(N__17960),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_5_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__26278),
            .in2(N__27194),
            .in3(N__17939),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_5_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__26804),
            .in2(N__26287),
            .in3(N__17918),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_5_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__20963),
            .in2(N__22543),
            .in3(N__17891),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_5_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__26194),
            .in2(N__23153),
            .in3(N__17867),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_5_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__20915),
            .in2(N__26198),
            .in3(N__18131),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_5_11_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__24263),
            .in2(N__20933),
            .in3(N__18107),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_5_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__23471),
            .in2(N__21035),
            .in3(N__18083),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_5_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__24175),
            .in2(N__20297),
            .in3(N__18080),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_8_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_5_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__23036),
            .in2(N__19859),
            .in3(N__18077),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_9_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_5_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__18074),
            .in2(N__21200),
            .in3(N__18068),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_5_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__23318),
            .in2(N__23378),
            .in3(N__18065),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_5_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_5_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__21257),
            .in2(N__23044),
            .in3(N__18047),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_5_12_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_5_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__21189),
            .in2(N__21146),
            .in3(N__18044),
            .lcout(\POWERLED.mult1_un47_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_5_12_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_5_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__23366),
            .in2(N__19763),
            .in3(N__18218),
            .lcout(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_5_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_5_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__23367),
            .in2(N__19805),
            .in3(N__18215),
            .lcout(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_5_13_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18212),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_13_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_13_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__18232),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_5_13_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_5_13_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_5_13_3  (
            .in0(N__20046),
            .in1(N__20047),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_13_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_13_4 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_13_4  (
            .in0(N__19952),
            .in1(_gnd_net_),
            .in2(N__18173),
            .in3(N__19974),
            .lcout(\POWERLED.mult1_un40_sum_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19879),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18187),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_13_7 .LUT_INIT=16'b1100110011000011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__18169),
            .in2(N__19976),
            .in3(N__19951),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__20074),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__18344),
            .in2(N__18268),
            .in3(N__18338),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2_c ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__18264),
            .in2(N__18335),
            .in3(N__18326),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3_c ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__18323),
            .in2(N__18313),
            .in3(N__18317),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4_c ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__18309),
            .in2(N__18287),
            .in3(N__18278),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5_c ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_14_5  (
            .in0(N__20195),
            .in1(N__18275),
            .in2(N__18269),
            .in3(N__18251),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6_c ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18248),
            .in3(N__18239),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(\POWERLED.mult1_un68_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18236),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__18233),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__18461),
            .in2(N__18361),
            .in3(N__18443),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__18357),
            .in2(N__20252),
            .in3(N__18431),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__20099),
            .in2(N__20231),
            .in3(N__18422),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__20213),
            .in2(N__20107),
            .in3(N__18413),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_15_5  (
            .in0(N__18387),
            .in1(N__20168),
            .in2(N__18362),
            .in3(N__18401),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20135),
            .in3(N__18398),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20098),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_12_LC_6_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_12_LC_6_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_12_LC_6_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_12_LC_6_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18779),
            .lcout(\PCH_PWRGD.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32489),
            .ce(N__18716),
            .sr(N__18936));
    defparam \PCH_PWRGD.count_2_LC_6_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_2_LC_6_2_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_2_LC_6_2_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \PCH_PWRGD.count_2_LC_6_2_0  (
            .in0(N__18841),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18882),
            .lcout(\PCH_PWRGD.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32686),
            .ce(N__18714),
            .sr(N__18935));
    defparam \PCH_PWRGD.count_RNIFV674_2_LC_6_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIFV674_2_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIFV674_2_LC_6_2_2 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \PCH_PWRGD.count_RNIFV674_2_LC_6_2_2  (
            .in0(N__18677),
            .in1(N__18829),
            .in2(N__18845),
            .in3(N__18880),
            .lcout(\PCH_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_6_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_6_2_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_6_2_3  (
            .in0(N__18881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18840),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIFV674_0_2_LC_6_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIFV674_0_2_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIFV674_0_2_LC_6_2_4 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \PCH_PWRGD.count_RNIFV674_0_2_LC_6_2_4  (
            .in0(N__18679),
            .in1(N__18830),
            .in2(N__18821),
            .in3(N__18818),
            .lcout(\PCH_PWRGD.un12_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI37554_12_LC_6_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI37554_12_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI37554_12_LC_6_2_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNI37554_12_LC_6_2_6  (
            .in0(N__18678),
            .in1(N__18785),
            .in2(_gnd_net_),
            .in3(N__18775),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(\PCH_PWRGD.countZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIORHA4_0_10_LC_6_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIORHA4_0_10_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIORHA4_0_10_LC_6_2_7 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \PCH_PWRGD.count_RNIORHA4_0_10_LC_6_2_7  (
            .in0(N__18756),
            .in1(N__18740),
            .in2(N__18722),
            .in3(N__18676),
            .lcout(\PCH_PWRGD.un12_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_6_3_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_6_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_6_3_0  (
            .in0(N__29549),
            .in1(N__18488),
            .in2(N__18509),
            .in3(N__18508),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_1_LC_6_3_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_6_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_6_3_1  (
            .in0(N__29543),
            .in1(N__18476),
            .in2(_gnd_net_),
            .in3(N__18464),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_2_LC_6_3_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_6_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_6_3_2  (
            .in0(N__29550),
            .in1(N__19085),
            .in2(_gnd_net_),
            .in3(N__19073),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_3_LC_6_3_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_6_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_6_3_3  (
            .in0(N__29544),
            .in1(N__19069),
            .in2(_gnd_net_),
            .in3(N__19055),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_4_LC_6_3_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_6_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_6_3_4  (
            .in0(N__29551),
            .in1(N__19052),
            .in2(_gnd_net_),
            .in3(N__19040),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_5_LC_6_3_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_6_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_6_3_5  (
            .in0(N__29545),
            .in1(N__19037),
            .in2(_gnd_net_),
            .in3(N__19025),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_6_LC_6_3_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_6_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_6_3_6  (
            .in0(N__29552),
            .in1(N__19022),
            .in2(_gnd_net_),
            .in3(N__19010),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_7_LC_6_3_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_6_3_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_6_3_7  (
            .in0(N__29546),
            .in1(N__19007),
            .in2(_gnd_net_),
            .in3(N__18995),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__32634),
            .ce(),
            .sr(N__19114));
    defparam \RSMRST_PWRGD.count_8_LC_6_4_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_6_4_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_6_4_0  (
            .in0(N__29567),
            .in1(N__18991),
            .in2(_gnd_net_),
            .in3(N__18977),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__32887),
            .ce(),
            .sr(N__19115));
    defparam \RSMRST_PWRGD.count_9_LC_6_4_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_6_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_6_4_1  (
            .in0(N__29563),
            .in1(N__18974),
            .in2(_gnd_net_),
            .in3(N__18962),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__32887),
            .ce(),
            .sr(N__19115));
    defparam \RSMRST_PWRGD.count_10_LC_6_4_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_6_4_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_6_4_2  (
            .in0(N__29564),
            .in1(N__18959),
            .in2(_gnd_net_),
            .in3(N__18947),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__32887),
            .ce(),
            .sr(N__19115));
    defparam \RSMRST_PWRGD.count_11_LC_6_4_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_6_4_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_6_4_3  (
            .in0(N__29561),
            .in1(N__19208),
            .in2(_gnd_net_),
            .in3(N__19196),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__32887),
            .ce(),
            .sr(N__19115));
    defparam \RSMRST_PWRGD.count_12_LC_6_4_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_6_4_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_6_4_4  (
            .in0(N__29565),
            .in1(N__19192),
            .in2(_gnd_net_),
            .in3(N__19178),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__32887),
            .ce(),
            .sr(N__19115));
    defparam \RSMRST_PWRGD.count_13_LC_6_4_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_6_4_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_6_4_5  (
            .in0(N__29562),
            .in1(N__19174),
            .in2(_gnd_net_),
            .in3(N__19160),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__32887),
            .ce(),
            .sr(N__19115));
    defparam \RSMRST_PWRGD.count_14_LC_6_4_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_6_4_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_6_4_6  (
            .in0(N__29566),
            .in1(N__19157),
            .in2(_gnd_net_),
            .in3(N__19145),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__32887),
            .ce(),
            .sr(N__19115));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(N__27453),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_6_5_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_6_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__19139),
            .in2(_gnd_net_),
            .in3(N__19142),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32899),
            .ce(N__19127),
            .sr(N__19104));
    defparam \POWERLED.count_RNI_2_LC_6_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_2_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_2_LC_6_6_0 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.count_RNI_2_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19252),
            .in3(N__19326),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_3_LC_6_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_3_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_3_LC_6_6_1 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \POWERLED.count_RNI_3_LC_6_6_1  (
            .in0(N__20640),
            .in1(N__20730),
            .in2(N__19088),
            .in3(N__19287),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlt15_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_7_LC_6_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_7_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_7_LC_6_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_7_LC_6_6_2  (
            .in0(N__19513),
            .in1(N__19548),
            .in2(N__19376),
            .in3(N__19591),
            .lcout(\POWERLED.un79_clk_100khzlto15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_6_6_3 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_6_6_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_6_6_3  (
            .in0(N__31998),
            .in1(N__25218),
            .in2(_gnd_net_),
            .in3(N__25183),
            .lcout(\POWERLED.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_10_LC_6_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_10_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_10_LC_6_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_10_LC_6_6_4  (
            .in0(N__19410),
            .in1(N__20475),
            .in2(N__19464),
            .in3(N__21994),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_15_LC_6_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_15_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_15_LC_6_6_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.count_RNI_15_LC_6_6_5  (
            .in0(N__20685),
            .in1(N__19358),
            .in2(N__19352),
            .in3(N__19650),
            .lcout(\POWERLED.count_RNIZ0Z_15 ),
            .ltout(\POWERLED.count_RNIZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_6_6_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_6_6_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.curr_state_RNIFPNR_0_LC_6_6_6  (
            .in0(N__25219),
            .in1(N__31799),
            .in2(N__19349),
            .in3(N__31999),
            .lcout(\POWERLED.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_LC_6_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_LC_6_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__25140),
            .in2(N__25098),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\POWERLED.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_6_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_6_7_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_RNIB209_LC_6_7_1  (
            .in0(N__25030),
            .in1(N__19327),
            .in2(_gnd_net_),
            .in3(N__19298),
            .lcout(\POWERLED.un1_count_cry_1_c_RNIBZ0Z209 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_1 ),
            .carryout(\POWERLED.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_6_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_6_7_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_2_c_RNIC419_LC_6_7_2  (
            .in0(N__25036),
            .in1(N__19288),
            .in2(_gnd_net_),
            .in3(N__19259),
            .lcout(\POWERLED.un1_count_cry_2_c_RNICZ0Z419 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_2 ),
            .carryout(\POWERLED.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_6_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_6_7_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_3_c_RNID629_LC_6_7_3  (
            .in0(N__25031),
            .in1(N__19248),
            .in2(_gnd_net_),
            .in3(N__19211),
            .lcout(\POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_3 ),
            .carryout(\POWERLED.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_6_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_6_7_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNIE839_LC_6_7_4  (
            .in0(N__25034),
            .in1(N__20731),
            .in2(_gnd_net_),
            .in3(N__19559),
            .lcout(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_4 ),
            .carryout(\POWERLED.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_6_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_6_7_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNIFA49_LC_6_7_5  (
            .in0(N__25033),
            .in1(N__20641),
            .in2(_gnd_net_),
            .in3(N__19556),
            .lcout(\POWERLED.un1_count_cry_5_c_RNIFAZ0Z49 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_5 ),
            .carryout(\POWERLED.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_6_7_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_6_7_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_6_c_RNIGC59_LC_6_7_6  (
            .in0(N__25035),
            .in1(N__19549),
            .in2(_gnd_net_),
            .in3(N__19517),
            .lcout(\POWERLED.un1_count_cry_6_c_RNIGCZ0Z59 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_6 ),
            .carryout(\POWERLED.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_6_7_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_6_7_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_7_c_RNIHE69_LC_6_7_7  (
            .in0(N__25032),
            .in1(N__19506),
            .in2(_gnd_net_),
            .in3(N__19475),
            .lcout(\POWERLED.un1_count_cry_7_c_RNIHEZ0Z69 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_7 ),
            .carryout(\POWERLED.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_6_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_6_8_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_8_c_RNIIG79_LC_6_8_0  (
            .in0(N__25041),
            .in1(N__19587),
            .in2(_gnd_net_),
            .in3(N__19472),
            .lcout(\POWERLED.un1_count_cry_8_c_RNIIGZ0Z79 ),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(\POWERLED.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_6_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_6_8_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_9_c_RNIJI89_LC_6_8_1  (
            .in0(N__25038),
            .in1(_gnd_net_),
            .in2(N__19465),
            .in3(N__19421),
            .lcout(\POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_9 ),
            .carryout(\POWERLED.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_6_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_6_8_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_6_8_2  (
            .in0(N__25043),
            .in1(N__19411),
            .in2(_gnd_net_),
            .in3(N__19382),
            .lcout(\POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_10 ),
            .carryout(\POWERLED.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_6_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_6_8_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_11_c_RNISEH7_LC_6_8_3  (
            .in0(N__25037),
            .in1(N__21990),
            .in2(_gnd_net_),
            .in3(N__19379),
            .lcout(\POWERLED.un1_count_cry_11_c_RNISEHZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_11 ),
            .carryout(\POWERLED.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_6_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_6_8_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_12_c_RNITGI7_LC_6_8_4  (
            .in0(N__25042),
            .in1(N__20476),
            .in2(_gnd_net_),
            .in3(N__19661),
            .lcout(\POWERLED.un1_count_cry_12_c_RNITGIZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_12 ),
            .carryout(\POWERLED.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_6_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_6_8_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_6_8_5  (
            .in0(N__25039),
            .in1(N__20686),
            .in2(_gnd_net_),
            .in3(N__19658),
            .lcout(\POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_13 ),
            .carryout(\POWERLED.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_6_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_6_8_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_6_8_6  (
            .in0(N__19651),
            .in1(N__25040),
            .in2(_gnd_net_),
            .in3(N__19628),
            .lcout(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIA4NN_9_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIA4NN_9_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIA4NN_9_LC_6_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIA4NN_9_LC_6_8_7  (
            .in0(N__19613),
            .in1(N__31988),
            .in2(_gnd_net_),
            .in3(N__19606),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI496F5_2_LC_6_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI496F5_2_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI496F5_2_LC_6_9_0 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \POWERLED.dutycycle_RNI496F5_2_LC_6_9_0  (
            .in0(N__23884),
            .in1(N__20870),
            .in2(N__21786),
            .in3(N__20879),
            .lcout(\POWERLED.dutycycle_eena_1 ),
            .ltout(\POWERLED.dutycycle_eena_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN2MP8_2_LC_6_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN2MP8_2_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN2MP8_2_LC_6_9_1 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \POWERLED.dutycycle_RNIN2MP8_2_LC_6_9_1  (
            .in0(N__23778),
            .in1(N__19693),
            .in2(N__19568),
            .in3(N__20413),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNINQPO7_1_LC_6_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNINQPO7_1_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNINQPO7_1_LC_6_9_2 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \POWERLED.dutycycle_RNINQPO7_1_LC_6_9_2  (
            .in0(N__19711),
            .in1(N__23777),
            .in2(N__20510),
            .in3(N__19721),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIP27U5_0_LC_6_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIP27U5_0_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIP27U5_0_LC_6_9_3 .LUT_INIT=16'b0011000111111111;
    LogicCell40 \POWERLED.dutycycle_RNIP27U5_0_LC_6_9_3  (
            .in0(N__30524),
            .in1(N__19565),
            .in2(N__26941),
            .in3(N__23883),
            .lcout(\POWERLED.dutycycle_eena ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIELPT3_1_LC_6_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIELPT3_1_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIELPT3_1_LC_6_9_4 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \POWERLED.func_state_RNIELPT3_1_LC_6_9_4  (
            .in0(N__21776),
            .in1(N__30522),
            .in2(N__28124),
            .in3(N__20878),
            .lcout(\POWERLED.N_108_f0_1 ),
            .ltout(\POWERLED.N_108_f0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIP27U5_1_LC_6_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIP27U5_1_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIP27U5_1_LC_6_9_5 .LUT_INIT=16'b0011111100110111;
    LogicCell40 \POWERLED.dutycycle_RNIP27U5_1_LC_6_9_5  (
            .in0(N__30523),
            .in1(N__23882),
            .in2(N__19724),
            .in3(N__26475),
            .lcout(\POWERLED.dutycycle_eena_0 ),
            .ltout(\POWERLED.dutycycle_eena_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_6_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_6_9_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_1_LC_6_9_6 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \POWERLED.dutycycle_1_LC_6_9_6  (
            .in0(N__19712),
            .in1(N__20503),
            .in2(N__19715),
            .in3(N__23780),
            .lcout(\POWERLED.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33077),
            .ce(),
            .sr(N__22900));
    defparam \POWERLED.dutycycle_2_LC_6_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_6_9_7 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_2_LC_6_9_7 .LUT_INIT=16'b0111000011111000;
    LogicCell40 \POWERLED.dutycycle_2_LC_6_9_7  (
            .in0(N__23779),
            .in1(N__19703),
            .in2(N__19697),
            .in3(N__20414),
            .lcout(\POWERLED.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33077),
            .ce(),
            .sr(N__22900));
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_x1_LC_6_10_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_x1_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_x1_LC_6_10_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.func_state_0_sqmuxa_0_o2_x1_LC_6_10_0  (
            .in0(N__22484),
            .in1(N__24906),
            .in2(N__28073),
            .in3(N__22068),
            .lcout(),
            .ltout(\POWERLED.func_state_0_sqmuxa_0_o2_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_ns_LC_6_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_ns_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_ns_LC_6_10_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.func_state_0_sqmuxa_0_o2_ns_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__27445),
            .in2(N__19682),
            .in3(N__24857),
            .lcout(\POWERLED.N_209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBK1U_0_1_LC_6_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBK1U_0_1_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBK1U_0_1_LC_6_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.func_state_RNIBK1U_0_1_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__20441),
            .in2(_gnd_net_),
            .in3(N__30550),
            .lcout(),
            .ltout(\POWERLED.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN3GO3_6_LC_6_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN3GO3_6_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN3GO3_6_LC_6_10_3 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \POWERLED.dutycycle_RNIN3GO3_6_LC_6_10_3  (
            .in0(N__19814),
            .in1(N__19673),
            .in2(N__19679),
            .in3(N__26576),
            .lcout(\POWERLED.N_217_N_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIBVNS_0_4_LC_6_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIBVNS_0_4_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIBVNS_0_4_LC_6_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_clk_RNIBVNS_0_4_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__25758),
            .in2(_gnd_net_),
            .in3(N__28472),
            .lcout(),
            .ltout(\POWERLED.N_300_N_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI6K332_4_LC_6_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI6K332_4_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI6K332_4_LC_6_10_5 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \POWERLED.count_clk_RNI6K332_4_LC_6_10_5  (
            .in0(N__28068),
            .in1(N__27885),
            .in2(N__19676),
            .in3(N__27097),
            .lcout(\POWERLED.N_4548_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOBU76_6_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOBU76_6_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOBU76_6_LC_6_10_6 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \POWERLED.dutycycle_RNIOBU76_6_LC_6_10_6  (
            .in0(N__23893),
            .in1(N__19667),
            .in2(_gnd_net_),
            .in3(N__20396),
            .lcout(\POWERLED.dutycycle_eena_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6RAN_0_1_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6RAN_0_1_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6RAN_0_1_LC_6_10_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.func_state_RNI6RAN_0_1_LC_6_10_7  (
            .in0(N__24907),
            .in1(N__28072),
            .in2(_gnd_net_),
            .in3(N__27795),
            .lcout(\POWERLED.N_353_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJ27K7_14_LC_6_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJ27K7_14_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJ27K7_14_LC_6_11_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIJ27K7_14_LC_6_11_0  (
            .in0(N__19781),
            .in1(N__25756),
            .in2(N__21089),
            .in3(N__19790),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(\POWERLED.dutycycleZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_LC_6_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_LC_6_11_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_14_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19808),
            .in3(N__22940),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN3GO3_14_LC_6_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN3GO3_14_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN3GO3_14_LC_6_11_2 .LUT_INIT=16'b1100111111101111;
    LogicCell40 \POWERLED.dutycycle_RNIN3GO3_14_LC_6_11_2  (
            .in0(N__23298),
            .in1(N__24019),
            .in2(N__24107),
            .in3(N__21182),
            .lcout(),
            .ltout(\POWERLED.N_86_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEB706_14_LC_6_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEB706_14_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEB706_14_LC_6_11_3 .LUT_INIT=16'b0011111100000000;
    LogicCell40 \POWERLED.dutycycle_RNIEB706_14_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__23891),
            .in2(N__19793),
            .in3(N__23804),
            .lcout(\POWERLED.dutycycle_en_11 ),
            .ltout(\POWERLED.dutycycle_en_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_6_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_14_LC_6_11_4 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_14_LC_6_11_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.dutycycle_14_LC_6_11_4  (
            .in0(N__21088),
            .in1(N__19777),
            .in2(N__19784),
            .in3(N__25757),
            .lcout(\POWERLED.dutycycleZ1Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33090),
            .ce(),
            .sr(N__22878));
    defparam \POWERLED.dutycycle_RNI_1_15_LC_6_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_6_11_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_15_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(N__23380),
            .in2(N__21199),
            .in3(N__22939),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIN3GO3_1_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIN3GO3_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIN3GO3_1_LC_6_11_6 .LUT_INIT=16'b1110110011111111;
    LogicCell40 \POWERLED.func_state_RNIN3GO3_1_LC_6_11_6  (
            .in0(N__23299),
            .in1(N__24020),
            .in2(N__19754),
            .in3(N__24104),
            .lcout(),
            .ltout(\POWERLED.N_84_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIEB706_1_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIEB706_1_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIEB706_1_LC_6_11_7 .LUT_INIT=16'b0011111100000000;
    LogicCell40 \POWERLED.func_state_RNIEB706_1_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(N__23892),
            .in2(N__19727),
            .in3(N__23805),
            .lcout(\POWERLED.dutycycle_en_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_LC_6_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_LC_6_12_0 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \POWERLED.dutycycle_RNI_10_LC_6_12_0  (
            .in0(N__21019),
            .in1(N__24387),
            .in2(_gnd_net_),
            .in3(N__24248),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_6_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_10_LC_6_12_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_10_LC_6_12_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \POWERLED.dutycycle_10_LC_6_12_1  (
            .in0(N__21325),
            .in1(N__19850),
            .in2(N__25821),
            .in3(N__21122),
            .lcout(\POWERLED.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32949),
            .ce(),
            .sr(N__22879));
    defparam \POWERLED.dutycycle_RNI_0_13_LC_6_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_6_12_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_13_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__24249),
            .in2(_gnd_net_),
            .in3(N__23021),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_10_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_9_LC_6_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_6_12_3 .LUT_INIT=16'b1011010011010010;
    LogicCell40 \POWERLED.dutycycle_RNI_2_9_LC_6_12_3  (
            .in0(N__23256),
            .in1(N__24394),
            .in2(N__19865),
            .in3(N__22969),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_LC_6_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_LC_6_12_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_13_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19862),
            .in3(N__23022),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI45I67_10_LC_6_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI45I67_10_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI45I67_10_LC_6_12_5 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.dutycycle_RNI45I67_10_LC_6_12_5  (
            .in0(N__25797),
            .in1(N__19849),
            .in2(N__21326),
            .in3(N__21121),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(\POWERLED.dutycycleZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_9_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_6_12_6 .LUT_INIT=16'b1111110101000100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_9_LC_6_12_6  (
            .in0(N__21020),
            .in1(N__24388),
            .in2(N__19841),
            .in3(N__23255),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_4Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_11_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_6_12_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_11_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(N__19838),
            .in2(N__19832),
            .in3(N__23468),
            .lcout(\POWERLED.un1_dutycycle_53_50_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_6_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_6_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19829),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_6_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_6_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19985),
            .in3(N__20030),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_6_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_6_13_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19937),
            .in3(N__20015),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_6_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_6_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__27468),
            .in2(N__20012),
            .in3(N__19991),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_6_13_4 .C_ON=1'b0;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_6_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19988),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_6_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_6_13_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19975),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_6_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_6_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__19970),
            .in2(_gnd_net_),
            .in3(N__19950),
            .lcout(\POWERLED.mult1_un47_sum_s_4_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIL58K7_15_LC_6_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIL58K7_15_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIL58K7_15_LC_6_13_7 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIL58K7_15_LC_6_13_7  (
            .in0(N__19927),
            .in1(N__25801),
            .in2(N__19904),
            .in3(N__21061),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__19880),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__20057),
            .in2(N__20152),
            .in3(N__20243),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__20148),
            .in2(N__20240),
            .in3(N__20222),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__20219),
            .in2(N__20203),
            .in3(N__20207),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__20199),
            .in2(N__20177),
            .in3(N__20162),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_14_5  (
            .in0(N__20103),
            .in1(N__20159),
            .in2(N__20153),
            .in3(N__20126),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20123),
            .in3(N__20114),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20078),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_7_LC_6_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_7_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_7_LC_6_15_0 .LUT_INIT=16'b0000110100000100;
    LogicCell40 \POWERLED.dutycycle_RNI_11_7_LC_6_15_0  (
            .in0(N__20285),
            .in1(N__24357),
            .in2(N__20276),
            .in3(N__23100),
            .lcout(\POWERLED.dutycycle_RNI_11Z0Z_7 ),
            .ltout(\POWERLED.dutycycle_RNI_11Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_12_LC_6_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_6_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_12_LC_6_15_1  (
            .in0(N__23230),
            .in1(N__24179),
            .in2(N__20300),
            .in3(N__24344),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_9_LC_6_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_6_15_2 .LUT_INIT=16'b0101000001110101;
    LogicCell40 \POWERLED.dutycycle_RNI_5_9_LC_6_15_2  (
            .in0(N__26599),
            .in1(N__26391),
            .in2(N__24386),
            .in3(N__23228),
            .lcout(\POWERLED.un1_dutycycle_53_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFO3M8_8_LC_6_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFO3M8_8_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFO3M8_8_LC_6_15_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIFO3M8_8_LC_6_15_3  (
            .in0(N__21286),
            .in1(N__21304),
            .in2(N__25820),
            .in3(N__22672),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(\POWERLED.dutycycleZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_LC_6_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_LC_6_15_4 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.dutycycle_RNI_4_LC_6_15_4  (
            .in0(N__26600),
            .in1(_gnd_net_),
            .in2(N__20279),
            .in3(N__26392),
            .lcout(\POWERLED.un1_dutycycle_53_45_a0_1 ),
            .ltout(\POWERLED.un1_dutycycle_53_45_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_7_LC_6_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_6_15_5 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \POWERLED.dutycycle_RNI_3_7_LC_6_15_5  (
            .in0(N__24267),
            .in1(N__23108),
            .in2(N__20267),
            .in3(N__24343),
            .lcout(\POWERLED.un1_dutycycle_53_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_7_LC_6_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_7_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_7_LC_6_15_6 .LUT_INIT=16'b0010000011011000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_7_LC_6_15_6  (
            .in0(N__26601),
            .in1(N__23099),
            .in2(N__26405),
            .in3(N__24356),
            .lcout(\POWERLED.un1_dutycycle_53_13_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_LC_6_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_LC_6_15_7 .LUT_INIT=16'b1111011110111111;
    LogicCell40 \POWERLED.dutycycle_RNI_9_LC_6_15_7  (
            .in0(N__23229),
            .in1(N__24342),
            .in2(N__23128),
            .in3(N__26602),
            .lcout(\POWERLED.un1_dutycycle_53_13_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_7_1_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_7_1_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIB5IA5_2_LC_7_1_1  (
            .in0(N__21386),
            .in1(N__21380),
            .in2(N__21275),
            .in3(N__21392),
            .lcout(\HDA_STRAP.un4_count ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_7_2_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_7_2_0 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \HDA_STRAP.count_17_LC_7_2_0  (
            .in0(N__21445),
            .in1(N__24623),
            .in2(N__21578),
            .in3(N__21506),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32685),
            .ce(N__29397),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_1_2_LC_7_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_1_2_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_1_2_LC_7_2_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \HDA_STRAP.curr_state_RNO_1_2_LC_7_2_1  (
            .in0(N__21504),
            .in1(N__21564),
            .in2(_gnd_net_),
            .in3(N__21444),
            .lcout(),
            .ltout(\HDA_STRAP.N_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_7_2_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_7_2_2 .LUT_INIT=16'b0010111000001100;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_7_2_2  (
            .in0(N__21565),
            .in1(N__20374),
            .in2(N__20378),
            .in3(N__20309),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32685),
            .ce(N__29397),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_7_2_3 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_7_2_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_7_2_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_LC_7_2_3  (
            .in0(N__20375),
            .in1(N__21503),
            .in2(_gnd_net_),
            .in3(N__21570),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32685),
            .ce(N__29397),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_1_0_LC_7_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_1_0_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_1_0_LC_7_2_4 .LUT_INIT=16'b0011111110101010;
    LogicCell40 \HDA_STRAP.curr_state_RNO_1_0_LC_7_2_4  (
            .in0(N__20348),
            .in1(N__20333),
            .in2(N__30586),
            .in3(N__21505),
            .lcout(),
            .ltout(\HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_7_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_7_2_5 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_7_2_5  (
            .in0(_gnd_net_),
            .in1(N__21569),
            .in2(N__20336),
            .in3(N__20315),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32685),
            .ce(N__29397),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_7_2_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_7_2_6 .LUT_INIT=16'b1010001110101111;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_0_LC_7_2_6  (
            .in0(N__21443),
            .in1(N__20332),
            .in2(N__21523),
            .in3(N__30576),
            .lcout(\HDA_STRAP.curr_state_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_7  (
            .in0(_gnd_net_),
            .in1(N__21499),
            .in2(_gnd_net_),
            .in3(N__30302),
            .lcout(\HDA_STRAP.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_1_LC_7_3_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_1_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_1_LC_7_3_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.func_state_RNI_3_1_LC_7_3_0  (
            .in0(N__28177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27778),
            .lcout(\POWERLED.N_341 ),
            .ltout(\POWERLED.N_341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_7_3_1 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_7_3_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_7_3_1  (
            .in0(N__29249),
            .in1(_gnd_net_),
            .in2(N__20303),
            .in3(N__25595),
            .lcout(\POWERLED.un1_func_state25_6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_LC_7_3_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_LC_7_3_2 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \POWERLED.func_state_RNI_1_LC_7_3_2  (
            .in0(N__27103),
            .in1(N__27777),
            .in2(N__20816),
            .in3(N__22141),
            .lcout(\POWERLED.func_state_1_m2s2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_1_LC_7_3_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_1_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_1_LC_7_3_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.func_state_RNI_4_1_LC_7_3_3  (
            .in0(N__27779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25594),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_a3_1_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI2AJD2_LC_7_3_4 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI2AJD2_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI2AJD2_LC_7_3_4 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI2AJD2_LC_7_3_4  (
            .in0(N__28054),
            .in1(N__24778),
            .in2(N__20417),
            .in3(N__20384),
            .lcout(\POWERLED.N_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0RLE1_1_LC_7_3_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0RLE1_1_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0RLE1_1_LC_7_3_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.func_state_RNI0RLE1_1_LC_7_3_5  (
            .in0(N__28053),
            .in1(N__27876),
            .in2(N__22049),
            .in3(N__27102),
            .lcout(\POWERLED.N_275_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_LC_7_3_6 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_LC_7_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_LC_7_3_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.tmp_0_LC_7_3_6  (
            .in0(N__31885),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26032),
            .lcout(suswarn_n),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32569),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJ9IE1_0_11_LC_7_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJ9IE1_0_11_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJ9IE1_0_11_LC_7_4_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.count_off_RNIJ9IE1_0_11_LC_7_4_0  (
            .in0(N__28031),
            .in1(N__24779),
            .in2(_gnd_net_),
            .in3(N__21630),
            .lcout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMJCH1_1_LC_7_4_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMJCH1_1_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMJCH1_1_LC_7_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNIMJCH1_1_LC_7_4_2  (
            .in0(_gnd_net_),
            .in1(N__23949),
            .in2(_gnd_net_),
            .in3(N__28242),
            .lcout(\POWERLED.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_6_1_LC_7_4_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_6_1_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_6_1_LC_7_4_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.func_state_RNI_6_1_LC_7_4_3  (
            .in0(N__22190),
            .in1(N__22140),
            .in2(_gnd_net_),
            .in3(N__27775),
            .lcout(),
            .ltout(\POWERLED.g0_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBK1U_1_LC_7_4_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBK1U_1_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBK1U_1_LC_7_4_4 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \POWERLED.func_state_RNIBK1U_1_LC_7_4_4  (
            .in0(N__21827),
            .in1(N__30555),
            .in2(N__20399),
            .in3(N__29242),
            .lcout(\POWERLED.g0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHL0V1_0_LC_7_4_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHL0V1_0_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHL0V1_0_LC_7_4_5 .LUT_INIT=16'b0111001101110111;
    LogicCell40 \POWERLED.func_state_RNIHL0V1_0_LC_7_4_5  (
            .in0(N__21914),
            .in1(N__20761),
            .in2(N__27889),
            .in3(N__22230),
            .lcout(\POWERLED.func_state_1_m0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_4_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_4_6 .LUT_INIT=16'b0000001100010011;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_4_6  (
            .in0(N__27776),
            .in1(N__30554),
            .in2(N__29250),
            .in3(N__20999),
            .lcout(\POWERLED.dutycycle_1_0_iv_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_7_5_0 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_7_5_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_7_5_0  (
            .in0(N__22474),
            .in1(N__24946),
            .in2(_gnd_net_),
            .in3(N__22384),
            .lcout(\POWERLED.N_326_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_7_5_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_7_5_1 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \POWERLED.func_state_RNIMQ0F_1_LC_7_5_1  (
            .in0(N__28471),
            .in1(N__27740),
            .in2(N__24955),
            .in3(N__24849),
            .lcout(\POWERLED.func_state_RNIMQ0FZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_0_LC_7_5_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_0_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_0_LC_7_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_3_0_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22221),
            .lcout(\POWERLED.N_2171_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9TUV2_0_LC_7_5_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9TUV2_0_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9TUV2_0_LC_7_5_3 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \POWERLED.func_state_RNI9TUV2_0_LC_7_5_3  (
            .in0(N__21653),
            .in1(N__20429),
            .in2(N__21644),
            .in3(N__21811),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIG5G37_1_LC_7_5_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIG5G37_1_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIG5G37_1_LC_7_5_4 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \POWERLED.func_state_RNIG5G37_1_LC_7_5_4  (
            .in0(N__29231),
            .in1(N__21602),
            .in2(N__20423),
            .in3(N__21608),
            .lcout(\POWERLED.func_state_RNIG5G37Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_1_LC_7_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_1_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_1_LC_7_5_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.count_RNI_1_LC_7_5_5  (
            .in0(N__25136),
            .in1(N__25046),
            .in2(_gnd_net_),
            .in3(N__25078),
            .lcout(),
            .ltout(\POWERLED.count_RNI_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGBFE_1_LC_7_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGBFE_1_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGBFE_1_LC_7_5_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIGBFE_1_LC_7_5_6  (
            .in0(N__31890),
            .in1(_gnd_net_),
            .in2(N__20420),
            .in3(N__25109),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_7_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_7_5_7 .LUT_INIT=16'b0101011111010111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_7_5_7  (
            .in0(N__22385),
            .in1(N__22475),
            .in2(N__24956),
            .in3(N__31889),
            .lcout(\POWERLED.N_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_7_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_7_6_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_0_LC_7_6_0 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \POWERLED.dutycycle_0_LC_7_6_0  (
            .in0(N__20585),
            .in1(N__20591),
            .in2(N__23789),
            .in3(N__20570),
            .lcout(\POWERLED.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32776),
            .ce(),
            .sr(N__22903));
    defparam \POWERLED.func_state_RNIBVNS_0_LC_7_6_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_7_6_1 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_LC_7_6_1  (
            .in0(N__26884),
            .in1(N__25869),
            .in2(N__22247),
            .in3(N__27737),
            .lcout(\POWERLED.dutycycle_1_0_0 ),
            .ltout(\POWERLED.dutycycle_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJFRN7_0_LC_7_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJFRN7_0_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJFRN7_0_LC_7_6_2 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \POWERLED.dutycycle_RNIJFRN7_0_LC_7_6_2  (
            .in0(N__23758),
            .in1(N__20584),
            .in2(N__20573),
            .in3(N__20569),
            .lcout(\POWERLED.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_0_LC_7_6_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_0_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_0_LC_7_6_3 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \POWERLED.func_state_RNI_4_0_LC_7_6_3  (
            .in0(N__22243),
            .in1(N__21640),
            .in2(_gnd_net_),
            .in3(N__27739),
            .lcout(\POWERLED.un1_func_state25_4_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI12UT8_1_LC_7_6_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI12UT8_1_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI12UT8_1_LC_7_6_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \POWERLED.func_state_RNI12UT8_1_LC_7_6_4  (
            .in0(N__23757),
            .in1(N__21763),
            .in2(N__20555),
            .in3(N__20524),
            .lcout(\POWERLED.func_state ),
            .ltout(\POWERLED.func_state_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_1_LC_7_6_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_1_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_1_LC_7_6_5 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \POWERLED.func_state_RNIBVNS_1_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20513),
            .in3(N__25865),
            .lcout(\POWERLED.func_state_RNIBVNSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_7_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_7_6_6 .LUT_INIT=16'b1011111100011111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_7_6_6  (
            .in0(N__27738),
            .in1(N__21011),
            .in2(N__25871),
            .in3(N__22242),
            .lcout(\POWERLED.dutycycle_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_1_LC_7_6_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_1_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_1_LC_7_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNI_2_1_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__21639),
            .in2(_gnd_net_),
            .in3(N__27736),
            .lcout(\POWERLED.func_state_RNI_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI0M6O_13_LC_7_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI0M6O_13_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI0M6O_13_LC_7_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI0M6O_13_LC_7_7_0  (
            .in0(N__31987),
            .in1(N__20447),
            .in2(_gnd_net_),
            .in3(N__20455),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_13_LC_7_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_13_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_7_7_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_13_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20459),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32798),
            .ce(N__31763),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI2OIN_5_LC_7_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI2OIN_5_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI2OIN_5_LC_7_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI2OIN_5_LC_7_7_2  (
            .in0(N__31985),
            .in1(N__20702),
            .in2(_gnd_net_),
            .in3(N__20710),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_5_LC_7_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_5_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_7_7_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_5_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20714),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32798),
            .ce(N__31763),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI2P7O_14_LC_7_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI2P7O_14_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI2P7O_14_LC_7_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI2P7O_14_LC_7_7_4  (
            .in0(N__20657),
            .in1(N__32003),
            .in2(_gnd_net_),
            .in3(N__20665),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_14_LC_7_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_14_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_7_7_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_14_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20669),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32798),
            .ce(N__31763),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI4RJN_6_LC_7_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI4RJN_6_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI4RJN_6_LC_7_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI4RJN_6_LC_7_7_6  (
            .in0(N__31986),
            .in1(N__20612),
            .in2(_gnd_net_),
            .in3(N__20620),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_6_LC_7_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_6_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_7_7_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_6_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20624),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32798),
            .ce(N__31763),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHV5K7_13_LC_7_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHV5K7_13_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHV5K7_13_LC_7_8_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIHV5K7_13_LC_7_8_0  (
            .in0(N__20788),
            .in1(N__25717),
            .in2(N__20600),
            .in3(N__21103),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(\POWERLED.dutycycleZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN3GO3_13_LC_7_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN3GO3_13_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN3GO3_13_LC_7_8_1 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \POWERLED.dutycycle_RNIN3GO3_13_LC_7_8_1  (
            .in0(N__25718),
            .in1(N__24099),
            .in2(N__20606),
            .in3(N__28449),
            .lcout(),
            .ltout(\POWERLED.N_148_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEB706_13_LC_7_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEB706_13_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEB706_13_LC_7_8_2 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIEB706_13_LC_7_8_2  (
            .in0(N__23975),
            .in1(N__23948),
            .in2(N__20603),
            .in3(N__23742),
            .lcout(\POWERLED.dutycycle_en_10 ),
            .ltout(\POWERLED.dutycycle_en_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_7_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_13_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_13_LC_7_8_3 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \POWERLED.dutycycle_13_LC_7_8_3  (
            .in0(N__21104),
            .in1(N__25722),
            .in2(N__20792),
            .in3(N__20789),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32794),
            .ce(),
            .sr(N__22880));
    defparam \POWERLED.func_state_RNIOTGO_0_LC_7_8_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOTGO_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOTGO_0_LC_7_8_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.func_state_RNIOTGO_0_LC_7_8_4  (
            .in0(N__28055),
            .in1(N__20780),
            .in2(N__28250),
            .in3(N__30509),
            .lcout(),
            .ltout(\POWERLED.N_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIES0I2_0_LC_7_8_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIES0I2_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIES0I2_0_LC_7_8_5 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \POWERLED.func_state_RNIES0I2_0_LC_7_8_5  (
            .in0(N__21775),
            .in1(N__25723),
            .in2(N__20771),
            .in3(N__23974),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQF354_1_LC_7_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQF354_1_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQF354_1_LC_7_8_6 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \POWERLED.func_state_RNIQF354_1_LC_7_8_6  (
            .in0(N__28207),
            .in1(N__20768),
            .in2(N__20750),
            .in3(N__23741),
            .lcout(\POWERLED.count_clk_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_0_1_LC_7_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_1_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_1_LC_7_8_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_1_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23297),
            .in3(_gnd_net_),
            .lcout(\POWERLED.func_state_RNIBVNS_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIBVNS_1_4_LC_7_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIBVNS_1_4_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIBVNS_1_4_LC_7_9_0 .LUT_INIT=16'b0011011101110111;
    LogicCell40 \POWERLED.count_clk_RNIBVNS_1_4_LC_7_9_0  (
            .in0(N__28456),
            .in1(N__25854),
            .in2(N__22172),
            .in3(N__22131),
            .lcout(\POWERLED.un1_count_off_1_sqmuxa_8_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_0_LC_7_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_7_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_0_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__25581),
            .in2(_gnd_net_),
            .in3(N__20803),
            .lcout(\POWERLED.dutycycle_RNI_8Z0Z_0 ),
            .ltout(\POWERLED.dutycycle_RNI_8Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_2_LC_7_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_7_9_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_2_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20747),
            .in3(N__22132),
            .lcout(),
            .ltout(\POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_1_0_LC_7_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_1_0_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_1_0_LC_7_9_3 .LUT_INIT=16'b0011011110111111;
    LogicCell40 \POWERLED.func_state_RNIBVNS_1_0_LC_7_9_3  (
            .in0(N__25900),
            .in1(N__25728),
            .in2(N__20744),
            .in3(N__25582),
            .lcout(),
            .ltout(\POWERLED.func_state_RNIBVNS_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMUFP1_1_LC_7_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMUFP1_1_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMUFP1_1_LC_7_9_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \POWERLED.func_state_RNIMUFP1_1_LC_7_9_4  (
            .in0(N__26769),
            .in1(N__25901),
            .in2(N__20891),
            .in3(N__20888),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIES0I2_1_LC_7_9_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIES0I2_1_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIES0I2_1_LC_7_9_5 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \POWERLED.func_state_RNIES0I2_1_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__28066),
            .in2(N__20882),
            .in3(N__30484),
            .lcout(\POWERLED.N_171 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILP0F_2_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILP0F_2_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILP0F_2_LC_7_9_6 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \POWERLED.dutycycle_RNILP0F_2_LC_7_9_6  (
            .in0(N__26240),
            .in1(N__27768),
            .in2(N__30521),
            .in3(N__27092),
            .lcout(\POWERLED.N_283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_7_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_0_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(N__25727),
            .in2(_gnd_net_),
            .in3(N__25583),
            .lcout(\POWERLED.func_state_RNIBVNS_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_7_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_7_10_0 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_6_LC_7_10_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \POWERLED.dutycycle_6_LC_7_10_0  (
            .in0(N__23740),
            .in1(N__20839),
            .in2(N__20849),
            .in3(N__20828),
            .lcout(\POWERLED.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32948),
            .ce(),
            .sr(N__22905));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI92UT3_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI92UT3_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI92UT3_LC_7_10_1 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI92UT3_LC_7_10_1  (
            .in0(N__23904),
            .in1(N__25759),
            .in2(N__20864),
            .in3(N__20978),
            .lcout(\POWERLED.dutycycle_set_0_0 ),
            .ltout(\POWERLED.dutycycle_set_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM1P2B_6_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM1P2B_6_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM1P2B_6_LC_7_10_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \POWERLED.dutycycle_RNIM1P2B_6_LC_7_10_2  (
            .in0(N__23739),
            .in1(N__20840),
            .in2(N__20831),
            .in3(N__20827),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(\POWERLED.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_LC_7_10_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_LC_7_10_3  (
            .in0(N__26921),
            .in1(_gnd_net_),
            .in2(N__20819),
            .in3(N__26456),
            .lcout(\POWERLED.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_0_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_7_10_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_0_LC_7_10_4  (
            .in0(N__26457),
            .in1(N__26922),
            .in2(N__26184),
            .in3(N__26554),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_10_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_0_LC_7_10_5  (
            .in0(N__26923),
            .in1(N__26577),
            .in2(N__26750),
            .in3(N__26458),
            .lcout(\POWERLED.N_392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_3_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_7_10_6 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_3_LC_7_10_6  (
            .in0(N__26455),
            .in1(N__26682),
            .in2(_gnd_net_),
            .in3(N__26555),
            .lcout(),
            .ltout(\POWERLED.d_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_5_LC_7_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_7_10_7 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_5_LC_7_10_7  (
            .in0(N__26165),
            .in1(N__22547),
            .in2(N__20966),
            .in3(N__26504),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_0_LC_7_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_7_11_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_0_LC_7_11_0  (
            .in0(N__26389),
            .in1(N__26932),
            .in2(_gnd_net_),
            .in3(N__26462),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_3_LC_7_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_7_11_1 .LUT_INIT=16'b1110110011001000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_3_LC_7_11_1  (
            .in0(N__23131),
            .in1(N__26388),
            .in2(N__24424),
            .in3(N__26677),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_3 ),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_9_LC_7_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_7_11_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_9_LC_7_11_2  (
            .in0(N__26565),
            .in1(_gnd_net_),
            .in2(N__20939),
            .in3(N__23258),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_7_LC_7_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_7_11_3 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_7_LC_7_11_3  (
            .in0(N__23132),
            .in1(N__26568),
            .in2(N__20936),
            .in3(N__24264),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_LC_7_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_LC_7_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_5_LC_7_11_4  (
            .in0(N__26567),
            .in1(N__20921),
            .in2(N__26190),
            .in3(N__23259),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_9_LC_7_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_7_11_5 .LUT_INIT=16'b0001111100001010;
    LogicCell40 \POWERLED.dutycycle_RNI_6_9_LC_7_11_5  (
            .in0(N__23257),
            .in1(N__26566),
            .in2(N__20906),
            .in3(N__22505),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_13_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_11_LC_7_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_7_11_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_11_LC_7_11_6  (
            .in0(N__23467),
            .in1(N__22511),
            .in2(N__21050),
            .in3(N__21047),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_7_LC_7_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_7_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_7_LC_7_11_7 .LUT_INIT=16'b0001010100010111;
    LogicCell40 \POWERLED.dutycycle_RNI_10_7_LC_7_11_7  (
            .in0(N__23130),
            .in1(N__26387),
            .in2(N__24423),
            .in3(N__26564),
            .lcout(\POWERLED.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_7_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_7_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__26938),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__27019),
            .in2(N__26482),
            .in3(N__21002),
            .lcout(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__26265),
            .in2(N__27053),
            .in3(N__20990),
            .lcout(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_1 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_7_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__27017),
            .in2(N__26696),
            .in3(N__20987),
            .lcout(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_7_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__27042),
            .in2(N__26358),
            .in3(N__20984),
            .lcout(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__27018),
            .in2(N__26191),
            .in3(N__20981),
            .lcout(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_12_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__26578),
            .in2(N__27052),
            .in3(N__20969),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_7_12_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_7_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__27013),
            .in2(N__23129),
            .in3(N__21131),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_7_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_7_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__27020),
            .in2(N__24406),
            .in3(N__21128),
            .lcout(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIMPUT_LC_7_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIMPUT_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIMPUT_LC_7_13_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_8_c_RNIMPUT_LC_7_13_1  (
            .in0(N__25738),
            .in1(N__27024),
            .in2(N__23254),
            .in3(N__21125),
            .lcout(\POWERLED.dutycycle_rst_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_7_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__27021),
            .in2(N__24265),
            .in3(N__21113),
            .lcout(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__27025),
            .in2(N__23453),
            .in3(N__21110),
            .lcout(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__24152),
            .in2(N__27054),
            .in3(N__21107),
            .lcout(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__27029),
            .in2(N__23020),
            .in3(N__21092),
            .lcout(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_13_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__27022),
            .in2(N__21204),
            .in3(N__21074),
            .lcout(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_13_7  (
            .in0(N__27023),
            .in1(N__23371),
            .in2(_gnd_net_),
            .in3(N__21071),
            .lcout(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_LC_7_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_LC_7_14_0 .LUT_INIT=16'b1111100000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_12_LC_7_14_0  (
            .in0(N__23249),
            .in1(N__24268),
            .in2(N__23466),
            .in3(N__24158),
            .lcout(\POWERLED.g0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_9_LC_7_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_9_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_9_LC_7_14_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_9_LC_7_14_1  (
            .in0(N__23811),
            .in1(N__21245),
            .in2(N__23525),
            .in3(N__21232),
            .lcout(\POWERLED.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33050),
            .ce(),
            .sr(N__22902));
    defparam \POWERLED.dutycycle_RNI_6_12_LC_7_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_12_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_12_LC_7_14_2 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \POWERLED.dutycycle_RNI_6_12_LC_7_14_2  (
            .in0(N__23250),
            .in1(N__24269),
            .in2(N__23162),
            .in3(N__24159),
            .lcout(),
            .ltout(\POWERLED.g0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_13_LC_7_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_7_14_3 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_13_LC_7_14_3  (
            .in0(N__23040),
            .in1(N__24185),
            .in2(N__21266),
            .in3(N__21263),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI67G18_9_LC_7_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI67G18_9_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI67G18_9_LC_7_14_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.dutycycle_RNI67G18_9_LC_7_14_4  (
            .in0(N__21244),
            .in1(N__23521),
            .in2(N__21233),
            .in3(N__23810),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(\POWERLED.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_9_LC_7_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_7_14_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_9_LC_7_14_5  (
            .in0(N__23168),
            .in1(_gnd_net_),
            .in2(N__21221),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.g0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_12_LC_7_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_7_14_6 .LUT_INIT=16'b1010111000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_12_LC_7_14_6  (
            .in0(N__23449),
            .in1(N__24270),
            .in2(N__21218),
            .in3(N__24160),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_14_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_14_LC_7_14_7  (
            .in0(N__21205),
            .in1(_gnd_net_),
            .in2(N__21149),
            .in3(N__23035),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_7_LC_7_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_7_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_7_LC_7_15_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.dutycycle_7_LC_7_15_0  (
            .in0(N__21350),
            .in1(N__21362),
            .in2(N__21371),
            .in3(N__25805),
            .lcout(\POWERLED.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33139),
            .ce(),
            .sr(N__22907));
    defparam \POWERLED.count_clk_RNI1J4E2_0_4_LC_7_15_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI1J4E2_0_4_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI1J4E2_0_4_LC_7_15_1 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \POWERLED.count_clk_RNI1J4E2_0_4_LC_7_15_1  (
            .in0(N__24009),
            .in1(N__23946),
            .in2(N__28475),
            .in3(N__25734),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_36_and_i_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEB706_7_LC_7_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEB706_7_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEB706_7_LC_7_15_2 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \POWERLED.dutycycle_RNIEB706_7_LC_7_15_2  (
            .in0(N__24105),
            .in1(N__23809),
            .in2(N__21374),
            .in3(N__21335),
            .lcout(\POWERLED.dutycycle_RNIEB706Z0Z_7 ),
            .ltout(\POWERLED.dutycycle_RNIEB706Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN1M47_7_LC_7_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN1M47_7_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN1M47_7_LC_7_15_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIN1M47_7_LC_7_15_3  (
            .in0(N__21361),
            .in1(N__25733),
            .in2(N__21353),
            .in3(N__21349),
            .lcout(\POWERLED.dutycycleZ1Z_6 ),
            .ltout(\POWERLED.dutycycleZ1Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_7_LC_7_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_7_15_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_7_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21338),
            .in3(N__24008),
            .lcout(\POWERLED.un1_clk_100khz_36_and_i_0_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI1J4E2_4_LC_7_15_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI1J4E2_4_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI1J4E2_4_LC_7_15_5 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \POWERLED.count_clk_RNI1J4E2_4_LC_7_15_5  (
            .in0(N__28466),
            .in1(N__23945),
            .in2(_gnd_net_),
            .in3(N__25732),
            .lcout(\POWERLED.dutycycle_eena_3_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN3GO3_10_LC_7_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN3GO3_10_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN3GO3_10_LC_7_15_6 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \POWERLED.dutycycle_RNIN3GO3_10_LC_7_15_6  (
            .in0(N__24106),
            .in1(N__28470),
            .in2(N__25793),
            .in3(N__24266),
            .lcout(),
            .ltout(\POWERLED.N_143_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEB706_10_LC_7_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEB706_10_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEB706_10_LC_7_15_7 .LUT_INIT=16'b0100000011001100;
    LogicCell40 \POWERLED.dutycycle_RNIEB706_10_LC_7_15_7  (
            .in0(N__24010),
            .in1(N__23812),
            .in2(N__21329),
            .in3(N__23947),
            .lcout(\POWERLED.dutycycle_en_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_7_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_8_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_8_LC_7_16_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \POWERLED.dutycycle_8_LC_7_16_5  (
            .in0(N__21308),
            .in1(N__22673),
            .in2(N__21290),
            .in3(N__25822),
            .lcout(\POWERLED.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33052),
            .ce(),
            .sr(N__22868));
    defparam \HDA_STRAP.count_RNI5DB61_6_LC_8_1_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI5DB61_6_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI5DB61_6_LC_8_1_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNI5DB61_6_LC_8_1_0  (
            .in0(N__24484),
            .in1(N__24568),
            .in2(N__24524),
            .in3(N__24460),
            .lcout(\HDA_STRAP.un4_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_8_1_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_8_1_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNIBJB61_7_LC_8_1_1  (
            .in0(N__24439),
            .in1(N__24499),
            .in2(N__24545),
            .in3(N__24709),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI0NIR1_14_LC_8_1_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI0NIR1_14_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI0NIR1_14_LC_8_1_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \HDA_STRAP.count_RNI0NIR1_14_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__24679),
            .in2(N__21395),
            .in3(N__24694),
            .lcout(\HDA_STRAP.un4_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_8_1_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_8_1_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \HDA_STRAP.count_RNI4CB61_17_LC_8_1_3  (
            .in0(N__23587),
            .in1(N__24664),
            .in2(N__23624),
            .in3(N__24637),
            .lcout(\HDA_STRAP.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI2L821_2_LC_8_1_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_8_1_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNI2L821_2_LC_8_1_4  (
            .in0(N__23539),
            .in1(N__23554),
            .in2(N__23573),
            .in3(N__24583),
            .lcout(\HDA_STRAP.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIH91A_1_LC_8_1_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIH91A_1_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIH91A_1_LC_8_1_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \HDA_STRAP.curr_state_RNIH91A_1_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(N__21522),
            .in2(_gnd_net_),
            .in3(N__21563),
            .lcout(\HDA_STRAP.curr_state_RNIH91AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_8_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_8_2_1 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \HDA_STRAP.count_6_LC_8_2_1  (
            .in0(N__21574),
            .in1(N__21508),
            .in2(N__24557),
            .in3(N__21452),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32748),
            .ce(N__29396),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_8_2_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_8_2_2 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \HDA_STRAP.count_8_LC_8_2_2  (
            .in0(N__21448),
            .in1(N__21577),
            .in2(N__21526),
            .in3(N__24509),
            .lcout(\HDA_STRAP.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32748),
            .ce(N__29396),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_8_2_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_8_2_3 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \HDA_STRAP.count_10_LC_8_2_3  (
            .in0(N__21572),
            .in1(N__21507),
            .in2(N__24473),
            .in3(N__21450),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32748),
            .ce(N__29396),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_8_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_8_2_4 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \HDA_STRAP.count_11_LC_8_2_4  (
            .in0(N__21447),
            .in1(N__21576),
            .in2(N__21525),
            .in3(N__24449),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32748),
            .ce(N__29396),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_8_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_8_2_5 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_8_2_5  (
            .in0(N__21571),
            .in1(N__21449),
            .in2(N__30310),
            .in3(N__21518),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32748),
            .ce(N__29396),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_0_LC_8_2_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_8_2_6 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \HDA_STRAP.count_0_LC_8_2_6  (
            .in0(N__21446),
            .in1(N__21575),
            .in2(N__21524),
            .in3(N__23594),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32748),
            .ce(N__29396),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_8_2_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_8_2_7 .LUT_INIT=16'b1000110011001100;
    LogicCell40 \HDA_STRAP.count_16_LC_8_2_7  (
            .in0(N__21573),
            .in1(N__24653),
            .in2(N__21527),
            .in3(N__21451),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32748),
            .ce(N__29396),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_3_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_3_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_3_0  (
            .in0(N__24952),
            .in1(N__22485),
            .in2(N__22040),
            .in3(N__22391),
            .lcout(\POWERLED.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_2_0_LC_8_3_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_2_0_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_2_0_LC_8_3_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_2_0_LC_8_3_1  (
            .in0(N__22392),
            .in1(N__24954),
            .in2(N__22490),
            .in3(N__25584),
            .lcout(\POWERLED.func_state_RNIBVNS_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6RAN_1_LC_8_3_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6RAN_1_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6RAN_1_LC_8_3_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.func_state_RNI6RAN_1_LC_8_3_2  (
            .in0(N__24953),
            .in1(N__28027),
            .in2(_gnd_net_),
            .in3(N__27797),
            .lcout(\POWERLED.func_state_RNI6RANZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBK1U_1_1_LC_8_3_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBK1U_1_1_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBK1U_1_1_LC_8_3_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \POWERLED.func_state_RNIBK1U_1_1_LC_8_3_4  (
            .in0(N__21416),
            .in1(N__28249),
            .in2(N__25596),
            .in3(N__24809),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m2s2_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHDGK3_1_LC_8_3_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHDGK3_1_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHDGK3_1_LC_8_3_5 .LUT_INIT=16'b1111000111111111;
    LogicCell40 \POWERLED.func_state_RNIHDGK3_1_LC_8_3_5  (
            .in0(N__27798),
            .in1(N__24780),
            .in2(N__21410),
            .in3(N__23954),
            .lcout(\POWERLED.N_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_rep1_LC_8_3_6 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_rep1_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_rep1_LC_8_3_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.tmp_0_rep1_LC_8_3_6  (
            .in0(N__22029),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26033),
            .lcout(SUSWARN_N_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32981),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI4VID3_0_LC_8_3_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI4VID3_0_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI4VID3_0_LC_8_3_7 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \POWERLED.func_state_RNI4VID3_0_LC_8_3_7  (
            .in0(N__21407),
            .in1(N__24746),
            .in2(N__21818),
            .in3(N__28160),
            .lcout(\POWERLED.func_state_1_m0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_en_LC_8_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_en_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_en_LC_8_4_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \POWERLED.count_off_en_LC_8_4_0  (
            .in0(N__21833),
            .in1(N__23695),
            .in2(N__24596),
            .in3(N__27902),
            .lcout(\POWERLED.count_off_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_154_LC_8_4_1 .C_ON=1'b0;
    defparam \POWERLED.G_154_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_154_LC_8_4_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.G_154_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(N__22030),
            .in2(_gnd_net_),
            .in3(N__26001),
            .lcout(G_154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_11_LC_8_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_11_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_11_LC_8_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.count_off_RNI_11_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28156),
            .lcout(\POWERLED.count_off_RNIZ0Z_11 ),
            .ltout(\POWERLED.count_off_RNIZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIJ9IE1_0_0_LC_8_4_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIJ9IE1_0_0_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIJ9IE1_0_0_LC_8_4_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.func_state_RNIJ9IE1_0_0_LC_8_4_3  (
            .in0(N__25579),
            .in1(N__27979),
            .in2(N__21656),
            .in3(N__24788),
            .lcout(\POWERLED.N_310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIBK1U_11_LC_8_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIBK1U_11_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIBK1U_11_LC_8_4_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.count_off_RNIBK1U_11_LC_8_4_4  (
            .in0(N__24808),
            .in1(N__25578),
            .in2(_gnd_net_),
            .in3(N__28157),
            .lcout(),
            .ltout(\POWERLED.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI18EF2_11_LC_8_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI18EF2_11_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI18EF2_11_LC_8_4_5 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \POWERLED.count_off_RNI18EF2_11_LC_8_4_5  (
            .in0(N__27106),
            .in1(N__23952),
            .in2(N__21647),
            .in3(N__21629),
            .lcout(),
            .ltout(\POWERLED.func_state_1_ss0_i_0_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHDGK3_0_1_LC_8_4_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHDGK3_0_1_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHDGK3_0_1_LC_8_4_6 .LUT_INIT=16'b1111111100001011;
    LogicCell40 \POWERLED.func_state_RNIHDGK3_0_1_LC_8_4_6  (
            .in0(N__27796),
            .in1(N__24777),
            .in2(N__21611),
            .in3(N__21810),
            .lcout(\POWERLED.func_state_RNIHDGK3_0Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNIHDGK3_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIB74H7_1_LC_8_4_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIB74H7_1_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIB74H7_1_LC_8_4_7 .LUT_INIT=16'b0100111000000000;
    LogicCell40 \POWERLED.func_state_RNIB74H7_1_LC_8_4_7  (
            .in0(N__21598),
            .in1(N__21587),
            .in2(N__21581),
            .in3(N__29200),
            .lcout(\POWERLED.func_state_RNIB74H7Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_8_5_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_8_5_0 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_8_5_0  (
            .in0(N__32402),
            .in1(N__28799),
            .in2(N__31517),
            .in3(N__32150),
            .lcout(\VPP_VDDQ.un9_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_LC_8_5_1 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_LC_8_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_LC_8_5_1  (
            .in0(N__22171),
            .in1(N__25870),
            .in2(N__22142),
            .in3(N__27105),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_287_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_0_LC_8_5_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_0_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_0_LC_8_5_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI_1_0_LC_8_5_2  (
            .in0(N__22222),
            .in1(N__22136),
            .in2(_gnd_net_),
            .in3(N__22170),
            .lcout(\POWERLED.func_state_RNI_1Z0Z_0 ),
            .ltout(\POWERLED.func_state_RNI_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBK1U_0_LC_8_5_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBK1U_0_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBK1U_0_LC_8_5_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.func_state_RNIBK1U_0_LC_8_5_3  (
            .in0(N__24807),
            .in1(_gnd_net_),
            .in2(N__21821),
            .in3(_gnd_net_),
            .lcout(\POWERLED.func_state_RNIBK1UZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIR2IB9_0_LC_8_5_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIR2IB9_0_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIR2IB9_0_LC_8_5_4 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \POWERLED.func_state_RNIR2IB9_0_LC_8_5_4  (
            .in0(N__21751),
            .in1(N__21728),
            .in2(N__23699),
            .in3(N__21694),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(\POWERLED.func_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1GMT1_0_LC_8_5_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1GMT1_0_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1GMT1_0_LC_8_5_5 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \POWERLED.func_state_RNI1GMT1_0_LC_8_5_5  (
            .in0(N__28048),
            .in1(N__21683),
            .in2(N__21674),
            .in3(N__27835),
            .lcout(\POWERLED.un1_clk_100khz_48_and_i_o2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_m1_0_a2_0_LC_8_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_m1_0_a2_0_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_m1_0_a2_0_LC_8_5_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.un1_m1_0_a2_0_LC_8_5_6  (
            .in0(N__22473),
            .in1(N__24951),
            .in2(_gnd_net_),
            .in3(N__24845),
            .lcout(\POWERLED.un1_N_3_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_52_and_i_0_0_LC_8_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_52_and_i_0_0_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_52_and_i_0_0_LC_8_5_7 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \POWERLED.un1_clk_100khz_52_and_i_0_0_LC_8_5_7  (
            .in0(N__24950),
            .in1(N__22472),
            .in2(N__28067),
            .in3(N__22386),
            .lcout(\POWERLED.un1_clk_100khz_52_and_i_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0RLE1_0_1_LC_8_6_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0RLE1_0_1_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0RLE1_0_1_LC_8_6_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.func_state_RNI0RLE1_0_1_LC_8_6_0  (
            .in0(N__28052),
            .in1(N__22048),
            .in2(N__27880),
            .in3(N__27104),
            .lcout(),
            .ltout(\POWERLED.N_275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI80TT3_LC_8_6_1 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI80TT3_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI80TT3_LC_8_6_1 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI80TT3_LC_8_6_1  (
            .in0(N__23953),
            .in1(N__21671),
            .in2(N__21659),
            .in3(N__25782),
            .lcout(\POWERLED.dutycycle_set_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_0_LC_8_6_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_0_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_0_LC_8_6_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.func_state_RNI_2_0_LC_8_6_2  (
            .in0(N__27733),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22245),
            .lcout(\POWERLED.func_state_RNI_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_5_1_LC_8_6_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_5_1_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_5_1_LC_8_6_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI_5_1_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__25580),
            .in2(_gnd_net_),
            .in3(N__27732),
            .lcout(\POWERLED.func_state_RNI_5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_1_LC_8_6_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_1_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_1_LC_8_6_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \POWERLED.func_state_RNI_1_1_LC_8_6_4  (
            .in0(N__27735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28460),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_48_and_i_o2_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIC4OR2_0_LC_8_6_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIC4OR2_0_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIC4OR2_0_LC_8_6_5 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \POWERLED.func_state_RNIC4OR2_0_LC_8_6_5  (
            .in0(N__30515),
            .in1(N__29201),
            .in2(N__21923),
            .in3(N__21920),
            .lcout(\POWERLED.func_state_RNIC4OR2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_0_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_0_LC_8_6_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \POWERLED.func_state_RNI_0_0_LC_8_6_6  (
            .in0(N__27734),
            .in1(N__22246),
            .in2(_gnd_net_),
            .in3(N__28170),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNICAC53_0_LC_8_6_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNICAC53_0_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNICAC53_0_LC_8_6_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.func_state_RNICAC53_0_LC_8_6_7  (
            .in0(N__21913),
            .in1(N__28097),
            .in2(N__21902),
            .in3(N__27659),
            .lcout(\POWERLED.func_state_RNICAC53_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_8_7_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_8_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21899),
            .lcout(\POWERLED.un85_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_13_LC_8_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_13_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_8_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_13_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25523),
            .lcout(\POWERLED.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32935),
            .ce(N__31218),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_14_LC_8_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_14_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_8_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_14_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25508),
            .lcout(\POWERLED.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32935),
            .ce(N__31218),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_2_LC_8_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_2_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_8_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_2_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25276),
            .lcout(\POWERLED.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32935),
            .ce(N__31218),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_3_LC_8_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_3_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_8_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_3_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25391),
            .lcout(\POWERLED.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32935),
            .ce(N__31218),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_4_LC_8_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_4_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_8_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_4_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25376),
            .lcout(\POWERLED.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32935),
            .ce(N__31218),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_8_7_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_7_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUI5O_12_LC_8_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUI5O_12_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUI5O_12_LC_8_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIUI5O_12_LC_8_8_0  (
            .in0(N__21950),
            .in1(N__32002),
            .in2(_gnd_net_),
            .in3(N__21961),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_12_LC_8_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_12_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_8_8_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_12_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21965),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32944),
            .ce(N__31767),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIHTPD_2_LC_8_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIHTPD_2_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIHTPD_2_LC_8_8_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNIHTPD_2_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__21944),
            .in2(N__25277),
            .in3(N__31143),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIL756_13_LC_8_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIL756_13_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIL756_13_LC_8_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIL756_13_LC_8_8_3  (
            .in0(N__31146),
            .in1(N__21938),
            .in2(_gnd_net_),
            .in3(N__25522),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINA66_14_LC_8_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINA66_14_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINA66_14_LC_8_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNINA66_14_LC_8_8_4  (
            .in0(N__21932),
            .in1(N__31147),
            .in2(_gnd_net_),
            .in3(N__25507),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPD76_15_LC_8_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPD76_15_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPD76_15_LC_8_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIPD76_15_LC_8_8_5  (
            .in0(N__31148),
            .in1(N__25478),
            .in2(_gnd_net_),
            .in3(N__25489),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIJ0RD_3_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIJ0RD_3_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIJ0RD_3_LC_8_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNIJ0RD_3_LC_8_8_6  (
            .in0(N__22262),
            .in1(N__31144),
            .in2(_gnd_net_),
            .in3(N__25390),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIL3SD_4_LC_8_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIL3SD_4_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIL3SD_4_LC_8_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIL3SD_4_LC_8_8_7  (
            .in0(N__31145),
            .in1(N__22256),
            .in2(_gnd_net_),
            .in3(N__25375),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_5_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26153),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_5 ),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_0_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_0_LC_8_9_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_0_LC_8_9_1  (
            .in0(N__26788),
            .in1(_gnd_net_),
            .in2(N__22250),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_10Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_1_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_1_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_1_LC_8_9_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \POWERLED.func_state_RNI_0_1_LC_8_9_2  (
            .in0(N__25597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27767),
            .lcout(\POWERLED.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_LC_8_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_LC_8_9_3 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_LC_8_9_3  (
            .in0(N__22244),
            .in1(N__22183),
            .in2(N__22169),
            .in3(N__22122),
            .lcout(\POWERLED.N_390 ),
            .ltout(\POWERLED.N_390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI39RS_0_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI39RS_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI39RS_0_LC_8_9_4 .LUT_INIT=16'b0111000011111111;
    LogicCell40 \POWERLED.func_state_RNI39RS_0_LC_8_9_4  (
            .in0(N__28065),
            .in1(N__22076),
            .in2(N__22052),
            .in3(N__22041),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_3_0_0_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIN7N72_0_LC_8_9_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIN7N72_0_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIN7N72_0_LC_8_9_5 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \POWERLED.func_state_RNIN7N72_0_LC_8_9_5  (
            .in0(N__24004),
            .in1(N__27859),
            .in2(N__22001),
            .in3(N__26016),
            .lcout(\POWERLED.dutycycle_eena_3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.slp_s3n_signal_2_LC_8_9_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.slp_s3n_signal_2_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.slp_s3n_signal_2_LC_8_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.slp_s3n_signal_2_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__22464),
            .in2(_gnd_net_),
            .in3(N__24853),
            .lcout(slp_s3n_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_m1_e_LC_8_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_m1_e_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_m1_e_LC_8_9_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \POWERLED.dutycycle_m1_e_LC_8_9_7  (
            .in0(N__22465),
            .in1(N__24922),
            .in2(_gnd_net_),
            .in3(N__22399),
            .lcout(\POWERLED.dutycycle_N_3_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILP0F_5_LC_8_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILP0F_5_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILP0F_5_LC_8_10_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \POWERLED.dutycycle_RNILP0F_5_LC_8_10_0  (
            .in0(N__22334),
            .in1(N__22328),
            .in2(_gnd_net_),
            .in3(N__30483),
            .lcout(\POWERLED.un1_clk_100khz_52_and_i_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_5_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_8_10_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_5_LC_8_10_1  (
            .in0(N__27794),
            .in1(_gnd_net_),
            .in2(N__26193),
            .in3(N__27093),
            .lcout(\POWERLED.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_0_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_8_10_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \POWERLED.dutycycle_RNI_6_0_LC_8_10_2  (
            .in0(N__22556),
            .in1(N__25447),
            .in2(_gnd_net_),
            .in3(N__28473),
            .lcout(\POWERLED.un1_dutycycle_172_sm3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI1U7M2_5_LC_8_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI1U7M2_5_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI1U7M2_5_LC_8_10_3 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \POWERLED.dutycycle_RNI1U7M2_5_LC_8_10_3  (
            .in0(N__26053),
            .in1(N__22555),
            .in2(N__26192),
            .in3(N__26039),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNICFHA6_5_LC_8_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNICFHA6_5_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNICFHA6_5_LC_8_10_4 .LUT_INIT=16'b0011001110111000;
    LogicCell40 \POWERLED.dutycycle_RNICFHA6_5_LC_8_10_4  (
            .in0(N__27113),
            .in1(N__22322),
            .in2(N__22316),
            .in3(N__30482),
            .lcout(),
            .ltout(\POWERLED.N_225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIG6629_5_LC_8_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIG6629_5_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIG6629_5_LC_8_10_5 .LUT_INIT=16'b0011000011111111;
    LogicCell40 \POWERLED.dutycycle_RNIG6629_5_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__22313),
            .in2(N__22304),
            .in3(N__23903),
            .lcout(\POWERLED.dutycycle_eena_14 ),
            .ltout(\POWERLED.dutycycle_eena_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNICPVSD_5_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNICPVSD_5_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNICPVSD_5_LC_8_10_6 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \POWERLED.dutycycle_RNICPVSD_5_LC_8_10_6  (
            .in0(N__22286),
            .in1(N__22270),
            .in2(N__22301),
            .in3(N__23703),
            .lcout(\POWERLED.dutycycleZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_8_10_7 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_5_LC_8_10_7 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_5_LC_8_10_7  (
            .in0(N__22271),
            .in1(N__22298),
            .in2(N__23738),
            .in3(N__22285),
            .lcout(\POWERLED.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33110),
            .ce(),
            .sr(N__22906));
    defparam \POWERLED.dutycycle_3_LC_8_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_3_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_3_LC_8_11_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \POWERLED.dutycycle_3_LC_8_11_0  (
            .in0(N__25767),
            .in1(N__22499),
            .in2(N__22582),
            .in3(N__22595),
            .lcout(\POWERLED.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33123),
            .ce(),
            .sr(N__22904));
    defparam \POWERLED.dutycycle_RNI59UL8_3_LC_8_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI59UL8_3_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI59UL8_3_LC_8_11_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.dutycycle_RNI59UL8_3_LC_8_11_1  (
            .in0(N__22498),
            .in1(N__22594),
            .in2(N__22583),
            .in3(N__25766),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(\POWERLED.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_11_2 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \POWERLED.dutycycle_RNI_7_3_LC_8_11_2  (
            .in0(N__26394),
            .in1(_gnd_net_),
            .in2(N__22562),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_3 ),
            .ltout(\POWERLED.dutycycle_RNI_7Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_0_LC_8_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_8_11_3 .LUT_INIT=16'b1110101011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_0_LC_8_11_3  (
            .in0(N__25891),
            .in1(N__26948),
            .in2(N__22559),
            .in3(N__26711),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_3_LC_8_11_4  (
            .in0(N__26395),
            .in1(N__26681),
            .in2(_gnd_net_),
            .in3(N__23134),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_7_LC_8_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_8_11_5 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \POWERLED.dutycycle_RNI_6_7_LC_8_11_5  (
            .in0(N__22520),
            .in1(_gnd_net_),
            .in2(N__23138),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_11_6 .LUT_INIT=16'b1011111111111010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_7_LC_8_11_6  (
            .in0(N__26575),
            .in1(N__22519),
            .in2(N__24425),
            .in3(N__23133),
            .lcout(\POWERLED.un1_dutycycle_53_13_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_LC_8_11_7 .LUT_INIT=16'b1110110011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_LC_8_11_7  (
            .in0(N__26390),
            .in1(N__24416),
            .in2(N__26693),
            .in3(N__26574),
            .lcout(\POWERLED.un1_dutycycle_53_31_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4VJH7_3_LC_8_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4VJH7_3_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4VJH7_3_LC_8_12_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI4VJH7_3_LC_8_12_0  (
            .in0(N__24083),
            .in1(N__22687),
            .in2(N__26692),
            .in3(N__22708),
            .lcout(\POWERLED.dutycycle_en_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4VJH7_4_LC_8_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4VJH7_4_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4VJH7_4_LC_8_12_1 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI4VJH7_4_LC_8_12_1  (
            .in0(N__22688),
            .in1(N__24081),
            .in2(N__26401),
            .in3(N__22704),
            .lcout(\POWERLED.dutycycle_RNI4VJH7Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4VJH7_8_LC_8_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4VJH7_8_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4VJH7_8_LC_8_12_2 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \POWERLED.dutycycle_RNI4VJH7_8_LC_8_12_2  (
            .in0(N__24082),
            .in1(N__24414),
            .in2(N__22709),
            .in3(N__22686),
            .lcout(\POWERLED.dutycycle_en_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_7_LC_8_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_8_12_3 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_7_LC_8_12_3  (
            .in0(N__24413),
            .in1(N__26357),
            .in2(_gnd_net_),
            .in3(N__23120),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_10_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_9_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_8_12_4 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_3_9_LC_8_12_4  (
            .in0(N__22741),
            .in1(N__23260),
            .in2(N__22652),
            .in3(N__24281),
            .lcout(\POWERLED.un1_dutycycle_53_10_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_7_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_8_12_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.dutycycle_RNI_7_7_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__26613),
            .in2(_gnd_net_),
            .in3(N__23119),
            .lcout(\POWERLED.un1_dutycycle_53_31_a7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_9_1_LC_8_12_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_9_1_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_9_1_LC_8_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_9_1_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26770),
            .lcout(\POWERLED.N_2200_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_12_LC_8_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_8_12_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \POWERLED.dutycycle_RNI_5_12_LC_8_12_7  (
            .in0(N__26852),
            .in1(N__24415),
            .in2(_gnd_net_),
            .in3(N__24167),
            .lcout(\POWERLED.un2_count_clk_17_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI7CVL8_4_LC_8_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI7CVL8_4_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI7CVL8_4_LC_8_13_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \POWERLED.dutycycle_RNI7CVL8_4_LC_8_13_0  (
            .in0(N__22631),
            .in1(N__25815),
            .in2(N__22619),
            .in3(N__22603),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_8_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_4_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_4_LC_8_13_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.dutycycle_4_LC_8_13_1  (
            .in0(N__25813),
            .in1(N__22630),
            .in2(N__22607),
            .in3(N__22618),
            .lcout(\POWERLED.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33128),
            .ce(),
            .sr(N__22901));
    defparam \POWERLED.dutycycle_RNIDP3K7_11_LC_8_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIDP3K7_11_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIDP3K7_11_LC_8_13_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.dutycycle_RNIDP3K7_11_LC_8_13_2  (
            .in0(N__22915),
            .in1(N__22720),
            .in2(N__25823),
            .in3(N__22924),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(\POWERLED.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_11_LC_8_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_8_13_3 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_11_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23048),
            .in3(N__23244),
            .lcout(\POWERLED.un1_dutycycle_53_50_a0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_12_LC_8_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_8_13_4 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_12_LC_8_13_4  (
            .in0(N__24168),
            .in1(N__24283),
            .in2(N__23465),
            .in3(N__23034),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_LC_8_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_LC_8_13_5 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_LC_8_13_5  (
            .in0(N__22970),
            .in1(N__22949),
            .in2(N__22943),
            .in3(N__24422),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_8_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_11_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_11_LC_8_13_6 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_11_LC_8_13_6  (
            .in0(N__22916),
            .in1(N__25814),
            .in2(N__22727),
            .in3(N__22925),
            .lcout(\POWERLED.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33128),
            .ce(),
            .sr(N__22901));
    defparam \POWERLED.dutycycle_RNI_11_LC_8_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_LC_8_13_7 .LUT_INIT=16'b1110111010001010;
    LogicCell40 \POWERLED.dutycycle_RNI_11_LC_8_13_7  (
            .in0(N__24282),
            .in1(N__23442),
            .in2(N__22745),
            .in3(N__23245),
            .lcout(\POWERLED.un1_dutycycle_53_50_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN3GO3_11_LC_8_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN3GO3_11_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN3GO3_11_LC_8_14_0 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \POWERLED.dutycycle_RNIN3GO3_11_LC_8_14_0  (
            .in0(N__28446),
            .in1(N__25810),
            .in2(N__24100),
            .in3(N__23433),
            .lcout(),
            .ltout(\POWERLED.N_144_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEB706_11_LC_8_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEB706_11_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEB706_11_LC_8_14_1 .LUT_INIT=16'b0100010011000100;
    LogicCell40 \POWERLED.dutycycle_RNIEB706_11_LC_8_14_1  (
            .in0(N__23944),
            .in1(N__23813),
            .in2(N__22730),
            .in3(N__24011),
            .lcout(\POWERLED.dutycycle_en_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIBVNS_4_LC_8_14_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIBVNS_4_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIBVNS_4_LC_8_14_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_clk_RNIBVNS_4_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__28448),
            .in2(_gnd_net_),
            .in3(N__25811),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNIBVNSZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOMK66_9_LC_8_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOMK66_9_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOMK66_9_LC_8_14_3 .LUT_INIT=16'b0011001011111111;
    LogicCell40 \POWERLED.dutycycle_RNIOMK66_9_LC_8_14_3  (
            .in0(N__24087),
            .in1(N__23174),
            .in2(N__23528),
            .in3(N__23951),
            .lcout(\POWERLED.dutycycle_eena_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFS4K7_12_LC_8_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFS4K7_12_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFS4K7_12_LC_8_14_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIFS4K7_12_LC_8_14_4  (
            .in0(N__23513),
            .in1(N__25812),
            .in2(N__23488),
            .in3(N__23635),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(\POWERLED.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_12_LC_8_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_8_14_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI_4_12_LC_8_14_5  (
            .in0(N__23434),
            .in1(_gnd_net_),
            .in2(N__23393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_51_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_14_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_15_LC_8_14_6  (
            .in0(N__23390),
            .in1(N__23384),
            .in2(N__23333),
            .in3(N__23330),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBVNS_9_LC_8_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBVNS_9_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBVNS_9_LC_8_14_7 .LUT_INIT=16'b1100110011111110;
    LogicCell40 \POWERLED.dutycycle_RNIBVNS_9_LC_8_14_7  (
            .in0(N__28447),
            .in1(N__24012),
            .in2(N__23306),
            .in3(N__23231),
            .lcout(\POWERLED.un1_clk_100khz_30_and_i_o2_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_7_LC_8_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_7_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_7_LC_8_15_0 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_8_7_LC_8_15_0  (
            .in0(N__23104),
            .in1(N__26622),
            .in2(N__24420),
            .in3(N__26380),
            .lcout(\POWERLED.dutycycle_RNI_8Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_LC_8_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_LC_8_15_1 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_LC_8_15_1  (
            .in0(N__26381),
            .in1(N__23106),
            .in2(N__26627),
            .in3(N__24398),
            .lcout(\POWERLED.N_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_3_LC_8_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_8_15_2 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_3_LC_8_15_2  (
            .in0(N__23107),
            .in1(N__26694),
            .in2(N__24421),
            .in3(N__26383),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_7_LC_8_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_8_15_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_7_LC_8_15_3  (
            .in0(N__26382),
            .in1(N__23105),
            .in2(_gnd_net_),
            .in3(N__26626),
            .lcout(),
            .ltout(\POWERLED.g0_i_a6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_12_LC_8_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_8_15_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_12_LC_8_15_4  (
            .in0(N__24402),
            .in1(N__24284),
            .in2(N__24188),
            .in3(N__24156),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIN3GO3_12_LC_8_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN3GO3_12_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN3GO3_12_LC_8_15_6 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \POWERLED.dutycycle_RNIN3GO3_12_LC_8_15_6  (
            .in0(N__25809),
            .in1(N__24157),
            .in2(N__28474),
            .in3(N__24080),
            .lcout(),
            .ltout(\POWERLED.N_145_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEB706_12_LC_8_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEB706_12_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEB706_12_LC_8_15_7 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIEB706_12_LC_8_15_7  (
            .in0(N__24013),
            .in1(N__23950),
            .in2(N__23816),
            .in3(N__23737),
            .lcout(\POWERLED.dutycycle_en_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_0_LC_9_1_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_0_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_0_LC_9_1_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_0_LC_9_1_0  (
            .in0(_gnd_net_),
            .in1(N__23620),
            .in2(N__23609),
            .in3(N__23608),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_9_1_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_1_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_9_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_1_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__23588),
            .in2(_gnd_net_),
            .in3(N__23576),
            .lcout(\HDA_STRAP.countZ0Z_1 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_0 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_1 ),
            .clk(N__32747),
            .ce(N__29395),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_9_1_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_2_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_9_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_2_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(N__23569),
            .in2(_gnd_net_),
            .in3(N__23558),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_2 ),
            .clk(N__32747),
            .ce(N__29395),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_9_1_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_3_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_9_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_3_LC_9_1_3  (
            .in0(_gnd_net_),
            .in1(N__23555),
            .in2(_gnd_net_),
            .in3(N__23543),
            .lcout(\HDA_STRAP.countZ0Z_3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_3 ),
            .clk(N__32747),
            .ce(N__29395),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_9_1_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_4_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_9_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_4_LC_9_1_4  (
            .in0(_gnd_net_),
            .in1(N__23540),
            .in2(_gnd_net_),
            .in3(N__24587),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_4 ),
            .clk(N__32747),
            .ce(N__29395),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_9_1_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_5_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_9_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_5_LC_9_1_5  (
            .in0(_gnd_net_),
            .in1(N__24584),
            .in2(_gnd_net_),
            .in3(N__24572),
            .lcout(\HDA_STRAP.countZ0Z_5 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_5 ),
            .clk(N__32747),
            .ce(N__29395),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_6_LC_9_1_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_6_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_6_LC_9_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_6_LC_9_1_6  (
            .in0(_gnd_net_),
            .in1(N__24569),
            .in2(_gnd_net_),
            .in3(N__24548),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_5 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_9_1_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_7_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_9_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_7_LC_9_1_7  (
            .in0(_gnd_net_),
            .in1(N__24538),
            .in2(_gnd_net_),
            .in3(N__24527),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_7 ),
            .clk(N__32747),
            .ce(N__29395),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_8_LC_9_2_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_8_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_8_LC_9_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_8_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(N__24520),
            .in2(_gnd_net_),
            .in3(N__24503),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_9_2_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_9_LC_9_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_9_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_9_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__24500),
            .in2(_gnd_net_),
            .in3(N__24488),
            .lcout(\HDA_STRAP.countZ0Z_9 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_8 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_9 ),
            .clk(N__32911),
            .ce(N__29401),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_10_LC_9_2_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_10_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_10_LC_9_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_10_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__24485),
            .in2(_gnd_net_),
            .in3(N__24464),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_11_LC_9_2_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_11_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_11_LC_9_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_11_LC_9_2_3  (
            .in0(_gnd_net_),
            .in1(N__24461),
            .in2(_gnd_net_),
            .in3(N__24443),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_9_2_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_12_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_9_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_12_LC_9_2_4  (
            .in0(_gnd_net_),
            .in1(N__24440),
            .in2(_gnd_net_),
            .in3(N__24428),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_12 ),
            .clk(N__32911),
            .ce(N__29401),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_9_2_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_13_LC_9_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_9_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_13_LC_9_2_5  (
            .in0(_gnd_net_),
            .in1(N__24710),
            .in2(_gnd_net_),
            .in3(N__24698),
            .lcout(\HDA_STRAP.countZ0Z_13 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_13 ),
            .clk(N__32911),
            .ce(N__29401),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_9_2_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_14_LC_9_2_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_9_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_14_LC_9_2_6  (
            .in0(_gnd_net_),
            .in1(N__24695),
            .in2(_gnd_net_),
            .in3(N__24683),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_14 ),
            .clk(N__32911),
            .ce(N__29401),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_9_2_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_15_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_9_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_15_LC_9_2_7  (
            .in0(_gnd_net_),
            .in1(N__24680),
            .in2(_gnd_net_),
            .in3(N__24668),
            .lcout(\HDA_STRAP.countZ0Z_15 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_15 ),
            .clk(N__32911),
            .ce(N__29401),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_16_LC_9_3_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_16_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_16_LC_9_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_16_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__24665),
            .in2(_gnd_net_),
            .in3(N__24647),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_17_LC_9_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNO_0_17_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_17_LC_9_3_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \HDA_STRAP.count_RNO_0_17_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(N__24644),
            .in2(_gnd_net_),
            .in3(N__24626),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_9_3_3 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_9_3_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_9_3_3  (
            .in0(N__27107),
            .in1(N__28030),
            .in2(N__27884),
            .in3(N__28159),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_o_N_305_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_9_3_4 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_9_3_4 .LUT_INIT=16'b1111010011111100;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_9_3_4  (
            .in0(N__28029),
            .in1(N__24611),
            .in2(N__24602),
            .in3(N__30547),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_3_5 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_3_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_3_5  (
            .in0(N__28200),
            .in1(N__28640),
            .in2(N__24599),
            .in3(N__27800),
            .lcout(\POWERLED.un1_func_state25_6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_ss0_i_0_x2_LC_9_3_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_ss0_i_0_x2_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_1_ss0_i_0_x2_LC_9_3_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.func_state_1_ss0_i_0_x2_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29238),
            .in3(N__30546),
            .lcout(\POWERLED.N_150_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJ9IE1_11_LC_9_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJ9IE1_11_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJ9IE1_11_LC_9_3_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.count_off_RNIJ9IE1_11_LC_9_3_7  (
            .in0(N__24781),
            .in1(N__28028),
            .in2(_gnd_net_),
            .in3(N__28158),
            .lcout(\POWERLED.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIR1479_9_LC_9_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIR1479_9_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIR1479_9_LC_9_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIR1479_9_LC_9_4_0  (
            .in0(N__24724),
            .in1(N__24733),
            .in2(_gnd_net_),
            .in3(N__30715),
            .lcout(\POWERLED.un3_count_off_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_9_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_10_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_9_4_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_10_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__30925),
            .in2(_gnd_net_),
            .in3(N__29944),
            .lcout(\POWERLED.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32942),
            .ce(N__30751),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_9_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_9_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_9_4_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.count_off_9_LC_9_4_2  (
            .in0(N__29980),
            .in1(_gnd_net_),
            .in2(N__30932),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32942),
            .ce(N__30751),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNISUHQ2_LC_9_4_3 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNISUHQ2_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNISUHQ2_LC_9_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNISUHQ2_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(N__30923),
            .in2(_gnd_net_),
            .in3(N__29981),
            .lcout(\POWERLED.count_off_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI4C959_10_LC_9_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI4C959_10_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI4C959_10_LC_9_4_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \POWERLED.count_off_RNI4C959_10_LC_9_4_4  (
            .in0(N__30924),
            .in1(N__24740),
            .in2(N__29948),
            .in3(N__30714),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(\POWERLED.count_offZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIR1479_0_9_LC_9_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIR1479_0_9_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIR1479_0_9_LC_9_4_5 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \POWERLED.count_off_RNIR1479_0_9_LC_9_4_5  (
            .in0(N__24734),
            .in1(N__24725),
            .in2(N__24716),
            .in3(N__30753),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIG5N6N1_11_LC_9_4_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIG5N6N1_11_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIG5N6N1_11_LC_9_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNIG5N6N1_11_LC_9_4_6  (
            .in0(N__25259),
            .in1(N__27548),
            .in2(N__24713),
            .in3(N__29831),
            .lcout(\POWERLED.count_off_RNIG5N6N1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDJM39_0_11_LC_9_4_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDJM39_0_11_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDJM39_0_11_LC_9_4_7 .LUT_INIT=16'b0001000100000101;
    LogicCell40 \POWERLED.count_off_RNIDJM39_0_11_LC_9_4_7  (
            .in0(N__29909),
            .in1(N__27599),
            .in2(N__27584),
            .in3(N__30752),
            .lcout(\POWERLED.un34_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_9_5_0 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_9_5_0 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \POWERLED.curr_state_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__25253),
            .in2(N__25223),
            .in3(N__25190),
            .lcout(\POWERLED.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32971),
            .ce(N__31766),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIHTOU_8_LC_9_5_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIHTOU_8_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIHTOU_8_LC_9_5_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNIHTOU_8_LC_9_5_1  (
            .in0(N__32401),
            .in1(N__32234),
            .in2(_gnd_net_),
            .in3(N__32207),
            .lcout(\VPP_VDDQ.count_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIM9AN_1_LC_9_5_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIM9AN_1_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIM9AN_1_LC_9_5_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIM9AN_1_LC_9_5_2  (
            .in0(N__28795),
            .in1(N__32400),
            .in2(_gnd_net_),
            .in3(N__31510),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_1 ),
            .ltout(\VPP_VDDQ.un1_count_2_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_1_LC_9_5_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_9_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \VPP_VDDQ.count_2_RNI_1_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25151),
            .in3(N__32149),
            .lcout(\VPP_VDDQ.count_2_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_9_5_4 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_9_5_4 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \POWERLED.count_1_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__25141),
            .in2(N__25099),
            .in3(N__25044),
            .lcout(\POWERLED.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32971),
            .ce(N__31766),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_9_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_9_5_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_0_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__25091),
            .in2(_gnd_net_),
            .in3(N__25045),
            .lcout(\POWERLED.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32971),
            .ce(N__31766),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.VCCST_EN_0_LC_9_5_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.VCCST_EN_0_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.VCCST_EN_0_LC_9_5_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.VCCST_EN_0_LC_9_5_7  (
            .in0(N__24942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24844),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIN6TD_5_LC_9_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIN6TD_5_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIN6TD_5_LC_9_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIN6TD_5_LC_9_6_0  (
            .in0(N__31202),
            .in1(N__25301),
            .in2(_gnd_net_),
            .in3(N__25360),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_5_LC_9_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_5_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_9_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_5_LC_9_6_1  (
            .in0(N__25361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33099),
            .ce(N__31223),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIP9UD_6_LC_9_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIP9UD_6_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIP9UD_6_LC_9_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIP9UD_6_LC_9_6_2  (
            .in0(N__31203),
            .in1(N__25295),
            .in2(_gnd_net_),
            .in3(N__25348),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_6_LC_9_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_6_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_9_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_6_LC_9_6_3  (
            .in0(N__25349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33099),
            .ce(N__31223),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNITF0E_8_LC_9_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNITF0E_8_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNITF0E_8_LC_9_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNITF0E_8_LC_9_6_4  (
            .in0(N__31204),
            .in1(N__25289),
            .in2(_gnd_net_),
            .in3(N__25333),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_8_LC_9_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_8_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_9_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_8_LC_9_6_5  (
            .in0(N__25334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33099),
            .ce(N__31223),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIVI1E_9_LC_9_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIVI1E_9_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIVI1E_9_LC_9_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIVI1E_9_LC_9_6_6  (
            .in0(N__31205),
            .in1(N__25283),
            .in2(_gnd_net_),
            .in3(N__25321),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_9_LC_9_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_9_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_9_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_9_LC_9_6_7  (
            .in0(N__25322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33099),
            .ce(N__31223),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_9_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_9_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__31352),
            .in2(N__31085),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_9_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_9_7_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_9_7_1  (
            .in0(N__31315),
            .in1(_gnd_net_),
            .in2(N__28609),
            .in3(N__25262),
            .lcout(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_9_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_9_7_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_9_7_2  (
            .in0(N__31251),
            .in1(_gnd_net_),
            .in2(N__28585),
            .in3(N__25379),
            .lcout(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_9_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_9_7_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_9_7_3  (
            .in0(N__31316),
            .in1(_gnd_net_),
            .in2(N__28503),
            .in3(N__25364),
            .lcout(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_9_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_9_7_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_9_7_4  (
            .in0(N__31252),
            .in1(_gnd_net_),
            .in2(N__31032),
            .in3(N__25352),
            .lcout(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_9_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_9_7_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_9_7_5  (
            .in0(N__31317),
            .in1(_gnd_net_),
            .in2(N__28560),
            .in3(N__25340),
            .lcout(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_9_7_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_9_7_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_9_7_6  (
            .in0(N__31253),
            .in1(_gnd_net_),
            .in2(N__28313),
            .in3(N__25337),
            .lcout(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_9_7_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_9_7_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_9_7_7  (
            .in0(N__31318),
            .in1(_gnd_net_),
            .in2(N__28528),
            .in3(N__25325),
            .lcout(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_7_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_9_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_9_8_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_9_8_0  (
            .in0(N__31319),
            .in1(_gnd_net_),
            .in2(N__31002),
            .in3(N__25310),
            .lcout(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_9_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_9_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28724),
            .in3(N__25307),
            .lcout(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_9_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_9_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_9_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__31424),
            .in2(_gnd_net_),
            .in3(N__25304),
            .lcout(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_10_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_9_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_9_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__31366),
            .in2(_gnd_net_),
            .in3(N__25526),
            .lcout(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_9_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_9_8_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_9_8_4  (
            .in0(N__31320),
            .in1(_gnd_net_),
            .in2(N__28693),
            .in3(N__25511),
            .lcout(\POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_9_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_9_8_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_9_8_5  (
            .in0(N__31321),
            .in1(_gnd_net_),
            .in2(N__28672),
            .in3(N__25496),
            .lcout(\POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_9_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_9_8_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_9_8_6  (
            .in0(N__28708),
            .in1(N__31322),
            .in2(_gnd_net_),
            .in3(N__25493),
            .lcout(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_15_LC_9_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_15_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_15_LC_9_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_15_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25490),
            .lcout(\POWERLED.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32943),
            .ce(N__31217),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0  (
            .in0(N__31206),
            .in1(N__25460),
            .in2(_gnd_net_),
            .in3(N__25471),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_7_LC_9_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_7_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_9_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_7_LC_9_9_1  (
            .in0(N__25472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32972),
            .ce(N__31207),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_0_LC_9_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_9_9_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_0_LC_9_9_2  (
            .in0(N__25454),
            .in1(N__26831),
            .in2(_gnd_net_),
            .in3(N__28424),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_9_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_9_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25436),
            .in3(N__25412),
            .lcout(\POWERLED.mult1_un47_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_9_6 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_9_6  (
            .in0(N__26097),
            .in1(N__26098),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBVNS_5_LC_9_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBVNS_5_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBVNS_5_LC_9_10_0 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \POWERLED.dutycycle_RNIBVNS_5_LC_9_10_0  (
            .in0(N__26170),
            .in1(N__25889),
            .in2(N__26063),
            .in3(N__26832),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m4_bm_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMUFP1_2_LC_9_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMUFP1_2_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMUFP1_2_LC_9_10_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \POWERLED.dutycycle_RNIMUFP1_2_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__25846),
            .in2(N__26042),
            .in3(N__25907),
            .lcout(\POWERLED.dutycycle_RNIMUFP1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_9_LC_9_10_2 .C_ON=1'b0;
    defparam \POWERLED.G_9_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_9_LC_9_10_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.G_9_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__32008),
            .in2(_gnd_net_),
            .in3(N__26031),
            .lcout(G_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_2_LC_9_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_9_10_3 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \POWERLED.dutycycle_RNI_1_2_LC_9_10_3  (
            .in0(N__25890),
            .in1(N__26171),
            .in2(N__26288),
            .in3(N__26707),
            .lcout(\POWERLED.un1_dutycycle_172_m4_bm_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_4_LC_9_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_4_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_4_LC_9_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_clk_RNI_1_4_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__28428),
            .in2(_gnd_net_),
            .in3(N__27077),
            .lcout(\POWERLED.N_20_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBVNS_2_LC_9_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBVNS_2_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBVNS_2_LC_9_10_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNIBVNS_2_LC_9_10_5  (
            .in0(N__25818),
            .in1(N__25603),
            .in2(_gnd_net_),
            .in3(N__26282),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMUFP1_0_LC_9_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMUFP1_0_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMUFP1_0_LC_9_10_6 .LUT_INIT=16'b0000110000011101;
    LogicCell40 \POWERLED.dutycycle_RNIMUFP1_0_LC_9_10_6  (
            .in0(N__25847),
            .in1(N__26840),
            .in2(N__25826),
            .in3(N__26833),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m3_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1U7M2_0_LC_9_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1U7M2_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1U7M2_0_LC_9_10_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.func_state_RNI1U7M2_0_LC_9_10_7  (
            .in0(N__25819),
            .in1(N__25604),
            .in2(N__25529),
            .in3(N__27119),
            .lcout(\POWERLED.un1_dutycycle_172_m3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_0_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_9_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_0_LC_9_11_0  (
            .in0(N__26487),
            .in1(N__26939),
            .in2(N__27098),
            .in3(N__28429),
            .lcout(\POWERLED.un1_dutycycle_96_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_0_LC_9_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_9_11_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_0_LC_9_11_1  (
            .in0(N__26940),
            .in1(N__26851),
            .in2(N__28461),
            .in3(N__26488),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_3_LC_9_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_9_11_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \POWERLED.dutycycle_RNI_3_3_LC_9_11_2  (
            .in0(N__26675),
            .in1(N__26273),
            .in2(_gnd_net_),
            .in3(N__26607),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_1_LC_9_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_9_11_3 .LUT_INIT=16'b1100001101001011;
    LogicCell40 \POWERLED.dutycycle_RNI_0_1_LC_9_11_3  (
            .in0(N__26834),
            .in1(N__26483),
            .in2(N__26810),
            .in3(N__26396),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_2_LC_9_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_9_11_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_2_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26807),
            .in3(N__26274),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_0_LC_9_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_0_LC_9_11_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.dutycycle_RNI_9_0_LC_9_11_5  (
            .in0(N__26795),
            .in1(N__26777),
            .in2(N__28462),
            .in3(N__26749),
            .lcout(\POWERLED.dutycycle_RNI_9Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_3_LC_9_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_9_11_6 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_3_LC_9_11_6  (
            .in0(N__26676),
            .in1(N__26393),
            .in2(N__26492),
            .in3(N__26606),
            .lcout(\POWERLED.un1_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_LC_9_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_LC_9_11_7 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_LC_9_11_7  (
            .in0(N__26489),
            .in1(N__26397),
            .in2(N__26286),
            .in3(N__26166),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_12_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_12_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_9_12_0  (
            .in0(N__27272),
            .in1(N__27254),
            .in2(N__27215),
            .in3(N__27160),
            .lcout(\VPP_VDDQ.un6_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_12_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_12_1  (
            .in0(N__27488),
            .in1(N__27506),
            .in2(N__27377),
            .in3(N__27524),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_12_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_12_2  (
            .in0(N__27173),
            .in1(N__27182),
            .in2(N__27176),
            .in3(N__27167),
            .lcout(\VPP_VDDQ.un6_count ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_12_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_9_12_3  (
            .in0(N__27319),
            .in1(N__27334),
            .in2(N__27290),
            .in3(N__27349),
            .lcout(\VPP_VDDQ.un6_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_12_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_9_12_4  (
            .in0(N__27304),
            .in1(N__27148),
            .in2(N__27236),
            .in3(N__27133),
            .lcout(\VPP_VDDQ.un6_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_9_13_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_9_13_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_9_13_0  (
            .in0(N__29588),
            .in1(N__27161),
            .in2(N__29162),
            .in3(N__29161),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_1_LC_9_13_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_9_13_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_9_13_1  (
            .in0(N__29584),
            .in1(N__27149),
            .in2(_gnd_net_),
            .in3(N__27137),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_2_LC_9_13_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_9_13_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_9_13_2  (
            .in0(N__29589),
            .in1(N__27134),
            .in2(_gnd_net_),
            .in3(N__27122),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_3_LC_9_13_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_9_13_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_9_13_3  (
            .in0(N__29585),
            .in1(N__27350),
            .in2(_gnd_net_),
            .in3(N__27338),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_4_LC_9_13_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_9_13_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_9_13_4  (
            .in0(N__29590),
            .in1(N__27335),
            .in2(_gnd_net_),
            .in3(N__27323),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_5_LC_9_13_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_9_13_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_9_13_5  (
            .in0(N__29586),
            .in1(N__27320),
            .in2(_gnd_net_),
            .in3(N__27308),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_6_LC_9_13_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_9_13_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_9_13_6  (
            .in0(N__29591),
            .in1(N__27305),
            .in2(_gnd_net_),
            .in3(N__27293),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_7_LC_9_13_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_9_13_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_9_13_7  (
            .in0(N__29587),
            .in1(N__27289),
            .in2(_gnd_net_),
            .in3(N__27275),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__33142),
            .ce(),
            .sr(N__29129));
    defparam \VPP_VDDQ.count_8_LC_9_14_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_9_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_9_14_0  (
            .in0(N__29583),
            .in1(N__27271),
            .in2(_gnd_net_),
            .in3(N__27257),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__33138),
            .ce(),
            .sr(N__29128));
    defparam \VPP_VDDQ.count_9_LC_9_14_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_9_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_9_14_1  (
            .in0(N__29579),
            .in1(N__27253),
            .in2(_gnd_net_),
            .in3(N__27239),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__33138),
            .ce(),
            .sr(N__29128));
    defparam \VPP_VDDQ.count_10_LC_9_14_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_9_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_9_14_2  (
            .in0(N__29580),
            .in1(N__27232),
            .in2(_gnd_net_),
            .in3(N__27218),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__33138),
            .ce(),
            .sr(N__29128));
    defparam \VPP_VDDQ.count_11_LC_9_14_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_9_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_9_14_3  (
            .in0(N__29577),
            .in1(N__27211),
            .in2(_gnd_net_),
            .in3(N__27197),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__33138),
            .ce(),
            .sr(N__29128));
    defparam \VPP_VDDQ.count_12_LC_9_14_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_9_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_9_14_4  (
            .in0(N__29581),
            .in1(N__27523),
            .in2(_gnd_net_),
            .in3(N__27509),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__33138),
            .ce(),
            .sr(N__29128));
    defparam \VPP_VDDQ.count_13_LC_9_14_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_9_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_9_14_5  (
            .in0(N__29578),
            .in1(N__27505),
            .in2(_gnd_net_),
            .in3(N__27491),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__33138),
            .ce(),
            .sr(N__29128));
    defparam \VPP_VDDQ.count_14_LC_9_14_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_9_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_9_14_6  (
            .in0(N__29582),
            .in1(N__27487),
            .in2(_gnd_net_),
            .in3(N__27473),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__33138),
            .ce(),
            .sr(N__29128));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_9_14_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_9_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__27449),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_9_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_9_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__27373),
            .in2(_gnd_net_),
            .in3(N__27380),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33140),
            .ce(N__29093),
            .sr(N__29121));
    defparam \POWERLED.count_off_RNIJLV69_5_LC_11_3_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJLV69_5_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJLV69_5_LC_11_3_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.count_off_RNIJLV69_5_LC_11_3_0  (
            .in0(N__30921),
            .in1(N__29761),
            .in2(N__27359),
            .in3(N__30761),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_11_3_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_11_3_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.count_off_5_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29762),
            .in3(N__30922),
            .lcout(\POWERLED.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32906),
            .ce(N__30782),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_11_3_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_14_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_11_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_14_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__30160),
            .in2(_gnd_net_),
            .in3(N__30917),
            .lcout(\POWERLED.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32906),
            .ce(N__30782),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_11_3_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_11_3_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_15_LC_11_3_4  (
            .in0(N__30185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30918),
            .lcout(\POWERLED.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32906),
            .ce(N__30782),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNILVQ39_15_LC_11_3_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNILVQ39_15_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNILVQ39_15_LC_11_3_5 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.count_off_RNILVQ39_15_LC_11_3_5  (
            .in0(N__30920),
            .in1(N__27563),
            .in2(N__30784),
            .in3(N__30184),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_11_3_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_8_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_11_3_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_8_LC_11_3_6  (
            .in0(N__30004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30919),
            .lcout(\POWERLED.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32906),
            .ce(N__30782),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIPU279_8_LC_11_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIPU279_8_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIPU279_8_LC_11_3_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.count_off_RNIPU279_8_LC_11_3_7  (
            .in0(N__30916),
            .in1(N__27557),
            .in2(N__30785),
            .in3(N__30005),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_11_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_11_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_2_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__29794),
            .in2(_gnd_net_),
            .in3(N__30931),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33029),
            .ce(N__30765),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDCS69_0_2_LC_11_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDCS69_0_2_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDCS69_0_2_LC_11_4_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \POWERLED.count_off_RNIDCS69_0_2_LC_11_4_1  (
            .in0(N__29776),
            .in1(N__27641),
            .in2(N__30777),
            .in3(N__27632),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI8GSR41_2_LC_11_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI8GSR41_2_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI8GSR41_2_LC_11_4_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNI8GSR41_2_LC_11_4_2  (
            .in0(N__27614),
            .in1(N__30116),
            .in2(N__27551),
            .in3(N__27539),
            .lcout(\POWERLED.un34_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNILO079_0_6_LC_11_4_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNILO079_0_6_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNILO079_0_6_LC_11_4_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \POWERLED.count_off_RNILO079_0_6_LC_11_4_3  (
            .in0(N__29819),
            .in1(N__27533),
            .in2(N__30778),
            .in3(N__28271),
            .lcout(\POWERLED.un34_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNIPOEQ2_LC_11_4_4 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNIPOEQ2_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNIPOEQ2_LC_11_4_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNIPOEQ2_LC_11_4_4  (
            .in0(N__29741),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30929),
            .lcout(\POWERLED.count_off_1_6 ),
            .ltout(\POWERLED.count_off_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNILO079_6_LC_11_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNILO079_6_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNILO079_6_LC_11_4_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \POWERLED.count_off_RNILO079_6_LC_11_4_5  (
            .in0(N__30734),
            .in1(N__28270),
            .in2(N__27527),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un3_count_off_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNILGAQ2_LC_11_4_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNILGAQ2_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNILGAQ2_LC_11_4_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNILGAQ2_LC_11_4_6  (
            .in0(_gnd_net_),
            .in1(N__29795),
            .in2(_gnd_net_),
            .in3(N__30930),
            .lcout(\POWERLED.count_off_1_2 ),
            .ltout(\POWERLED.count_off_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDCS69_2_LC_11_4_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDCS69_2_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDCS69_2_LC_11_4_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_off_RNIDCS69_2_LC_11_4_7  (
            .in0(N__30735),
            .in1(_gnd_net_),
            .in2(N__27635),
            .in3(N__27631),
            .lcout(\POWERLED.un3_count_off_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNINR179_7_LC_11_5_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNINR179_7_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNINR179_7_LC_11_5_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNINR179_7_LC_11_5_0  (
            .in0(N__30766),
            .in1(N__27607),
            .in2(_gnd_net_),
            .in3(N__27623),
            .lcout(\POWERLED.un3_count_off_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIQQFQ2_LC_11_5_1 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIQQFQ2_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIQQFQ2_LC_11_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNIQQFQ2_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__30032),
            .in2(_gnd_net_),
            .in3(N__30853),
            .lcout(\POWERLED.count_off_1_7 ),
            .ltout(\POWERLED.count_off_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNINR179_0_7_LC_11_5_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNINR179_0_7_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNINR179_0_7_LC_11_5_2 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \POWERLED.count_off_RNINR179_0_7_LC_11_5_2  (
            .in0(N__30787),
            .in1(N__27608),
            .in2(N__27617),
            .in3(N__30020),
            .lcout(\POWERLED.un34_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_11_5_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_7_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_11_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_7_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__30031),
            .in2(_gnd_net_),
            .in3(N__30857),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32907),
            .ce(N__30786),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNI570P2_LC_11_5_4 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNI570P2_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNI570P2_LC_11_5_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNI570P2_LC_11_5_4  (
            .in0(N__30854),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29921),
            .lcout(\POWERLED.count_off_1_11 ),
            .ltout(\POWERLED.count_off_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDJM39_11_LC_11_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDJM39_11_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDJM39_11_LC_11_5_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_off_RNIDJM39_11_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__27574),
            .in2(N__27587),
            .in3(N__30767),
            .lcout(\POWERLED.un3_count_off_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_11_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_11_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_11_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_11_LC_11_5_6  (
            .in0(N__30855),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29920),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32907),
            .ce(N__30786),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_11_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_11_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_6_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__29740),
            .in2(_gnd_net_),
            .in3(N__30856),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32907),
            .ce(N__30786),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIJ9IE1_0_LC_11_6_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIJ9IE1_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIJ9IE1_0_LC_11_6_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNIJ9IE1_0_LC_11_6_0  (
            .in0(N__28282),
            .in1(N__28262),
            .in2(_gnd_net_),
            .in3(N__28087),
            .lcout(),
            .ltout(\POWERLED.N_289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIU8AB2_7_LC_11_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIU8AB2_7_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIU8AB2_7_LC_11_6_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \POWERLED.count_clk_RNIU8AB2_7_LC_11_6_1  (
            .in0(N__28632),
            .in1(N__28241),
            .in2(N__28211),
            .in3(N__28208),
            .lcout(\POWERLED.N_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_8_1_LC_11_6_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_8_1_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_8_1_LC_11_6_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \POWERLED.func_state_RNI_8_1_LC_11_6_3  (
            .in0(N__28178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28120),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_2_tz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIRKB61_1_LC_11_6_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIRKB61_1_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIRKB61_1_LC_11_6_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \POWERLED.func_state_RNIRKB61_1_LC_11_6_4  (
            .in0(N__28283),
            .in1(N__28001),
            .in2(N__28100),
            .in3(N__27883),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_11_6_5 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_11_6_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_11_6_5  (
            .in0(N__27882),
            .in1(N__28088),
            .in2(N__28041),
            .in3(N__28281),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_304_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_1_LC_11_6_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_11_6_6 .LUT_INIT=16'b0010000000100011;
    LogicCell40 \POWERLED.func_state_RNIOGRS_1_LC_11_6_6  (
            .in0(N__28633),
            .in1(N__27881),
            .in2(N__27799),
            .in3(N__28340),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_4_LC_11_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_4_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_4_LC_11_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_4_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__28561),
            .in2(_gnd_net_),
            .in3(N__28510),
            .lcout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_2_LC_11_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_2_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_2_LC_11_7_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_2_LC_11_7_0  (
            .in0(N__28615),
            .in1(N__28534),
            .in2(N__27650),
            .in3(N__28591),
            .lcout(\POWERLED.N_352 ),
            .ltout(\POWERLED.N_352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_7_LC_11_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_7_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_7_LC_11_7_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \POWERLED.count_clk_RNI_7_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__28315),
            .in2(N__28643),
            .in3(N__30968),
            .lcout(\POWERLED.N_394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_11_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_11_7_2 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_11_7_2  (
            .in0(N__31607),
            .in1(N__33660),
            .in2(_gnd_net_),
            .in3(N__32001),
            .lcout(\VPP_VDDQ.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_11_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_11_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_1_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33431),
            .lcout(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_2_LC_11_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_2_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_2_LC_11_7_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \POWERLED.count_clk_RNI_2_LC_11_7_4  (
            .in0(N__28616),
            .in1(N__28592),
            .in2(N__28568),
            .in3(N__28535),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_4_LC_11_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_4_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_4_LC_11_7_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \POWERLED.count_clk_RNI_4_LC_11_7_5  (
            .in0(N__28511),
            .in1(N__28316),
            .in2(N__28478),
            .in3(N__30967),
            .lcout(\POWERLED.N_2182_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_7_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.count_clk_RNI_0_1_LC_11_7_6  (
            .in0(N__31039),
            .in1(N__31076),
            .in2(_gnd_net_),
            .in3(N__31051),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_9_LC_11_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_9_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_9_LC_11_7_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNI_9_LC_11_7_7  (
            .in0(N__28322),
            .in1(N__28314),
            .in2(N__28286),
            .in3(N__31003),
            .lcout(\POWERLED.count_clk_RNIZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_10_LC_11_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_10_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_11_8_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.count_clk_10_LC_11_8_0  (
            .in0(N__28736),
            .in1(_gnd_net_),
            .in2(N__31314),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33048),
            .ce(N__31201),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8SH6_10_LC_11_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8SH6_10_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8SH6_10_LC_11_8_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.count_clk_RNI8SH6_10_LC_11_8_1  (
            .in0(N__31162),
            .in1(N__31285),
            .in2(N__28745),
            .in3(N__28735),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(\POWERLED.count_clkZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_15_LC_11_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_15_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_15_LC_11_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_15_LC_11_8_2  (
            .in0(N__31367),
            .in1(N__31423),
            .in2(N__28712),
            .in3(N__28709),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_13_LC_11_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_13_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_13_LC_11_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_13_LC_11_8_3  (
            .in0(N__31345),
            .in1(N__28694),
            .in2(N__28676),
            .in3(N__28673),
            .lcout(\POWERLED.N_163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_11_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_0_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_11_8_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_clk_0_LC_11_8_4  (
            .in0(N__31286),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31346),
            .lcout(\POWERLED.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33048),
            .ce(N__31201),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_8_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_0_LC_11_8_5  (
            .in0(N__31347),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31283),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIQF8B_0_LC_11_8_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIQF8B_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIQF8B_0_LC_11_8_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNIQF8B_0_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__28655),
            .in2(N__28649),
            .in3(N__31161),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(\POWERLED.count_clkZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_LC_11_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_LC_11_8_7 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_LC_11_8_7  (
            .in0(N__31078),
            .in1(_gnd_net_),
            .in2(N__28646),
            .in3(N__31284),
            .lcout(\POWERLED.count_clk_RNIZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_11_9_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_11_9_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_11_9_0  (
            .in0(N__33397),
            .in1(N__33557),
            .in2(N__33297),
            .in3(N__28822),
            .lcout(\VPP_VDDQ.count_2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_4_LC_11_9_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_4_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_4_LC_11_9_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_4_LC_11_9_1  (
            .in0(N__33558),
            .in1(N__33277),
            .in2(N__28826),
            .in3(N__33402),
            .lcout(\VPP_VDDQ.count_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33100),
            .ce(N__32429),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_11_9_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_11_9_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_11_9_2  (
            .in0(N__28948),
            .in1(N__33567),
            .in2(N__33451),
            .in3(N__33282),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJ0QU_9_LC_11_9_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJ0QU_9_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJ0QU_9_LC_11_9_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIJ0QU_9_LC_11_9_3  (
            .in0(N__28805),
            .in1(_gnd_net_),
            .in2(N__28808),
            .in3(N__32363),
            .lcout(\VPP_VDDQ.count_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_9_LC_11_9_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_9_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_9_LC_11_9_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_9_LC_11_9_4  (
            .in0(N__33399),
            .in1(N__33560),
            .in2(N__28949),
            .in3(N__33281),
            .lcout(\VPP_VDDQ.count_2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33100),
            .ce(N__32429),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_1_LC_11_9_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_1_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_1_LC_11_9_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_1_LC_11_9_5  (
            .in0(N__33278),
            .in1(N__31541),
            .in2(N__33620),
            .in3(N__33401),
            .lcout(\VPP_VDDQ.count_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33100),
            .ce(N__32429),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_2_LC_11_9_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_2_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_2_LC_11_9_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_2_LC_11_9_6  (
            .in0(N__33398),
            .in1(N__33559),
            .in2(N__31484),
            .in3(N__33280),
            .lcout(\VPP_VDDQ.count_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33100),
            .ce(N__32429),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_5_LC_11_9_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_5_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_5_LC_11_9_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_5_LC_11_9_7  (
            .in0(N__33279),
            .in1(N__33400),
            .in2(N__33621),
            .in3(N__29006),
            .lcout(\VPP_VDDQ.count_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33100),
            .ce(N__32429),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI5BIU_0_2_LC_11_10_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI5BIU_0_2_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI5BIU_0_2_LC_11_10_0 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI5BIU_0_2_LC_11_10_0  (
            .in0(N__32359),
            .in1(N__31460),
            .in2(N__28874),
            .in3(N__31447),
            .lcout(\VPP_VDDQ.un9_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIBKLU_0_5_LC_11_10_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIBKLU_0_5_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIBKLU_0_5_LC_11_10_1 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIBKLU_0_5_LC_11_10_1  (
            .in0(N__28981),
            .in1(N__32361),
            .in2(N__28889),
            .in3(N__28898),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFQ6J3_1_LC_11_10_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFQ6J3_1_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFQ6J3_1_LC_11_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIFQ6J3_1_LC_11_10_2  (
            .in0(N__28775),
            .in1(N__28760),
            .in2(N__28754),
            .in3(N__28751),
            .lcout(\VPP_VDDQ.un9_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI9HKU_0_4_LC_11_10_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI9HKU_0_4_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI9HKU_0_4_LC_11_10_3 .LUT_INIT=16'b0000010000000111;
    LogicCell40 \VPP_VDDQ.count_2_RNI9HKU_0_4_LC_11_10_3  (
            .in0(N__28907),
            .in1(N__32360),
            .in2(N__31703),
            .in3(N__28918),
            .lcout(\VPP_VDDQ.un9_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI9HKU_4_LC_11_10_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI9HKU_4_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI9HKU_4_LC_11_10_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \VPP_VDDQ.count_2_RNI9HKU_4_LC_11_10_4  (
            .in0(N__32357),
            .in1(_gnd_net_),
            .in2(N__28919),
            .in3(N__28906),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_11_10_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_11_10_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_11_10_5  (
            .in0(N__33428),
            .in1(N__33268),
            .in2(N__33657),
            .in3(N__29002),
            .lcout(\VPP_VDDQ.count_2_1_5 ),
            .ltout(\VPP_VDDQ.count_2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIBKLU_5_LC_11_10_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIBKLU_5_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIBKLU_5_LC_11_10_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIBKLU_5_LC_11_10_6  (
            .in0(N__32358),
            .in1(_gnd_net_),
            .in2(N__28892),
            .in3(N__28885),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI5BIU_2_LC_11_10_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI5BIU_2_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI5BIU_2_LC_11_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI5BIU_2_LC_11_10_7  (
            .in0(N__31459),
            .in1(N__28870),
            .in2(_gnd_net_),
            .in3(N__32356),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_11_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__32135),
            .in2(N__28862),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_11_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__28844),
            .in2(_gnd_net_),
            .in3(N__28838),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_11_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__31448),
            .in2(_gnd_net_),
            .in3(N__28835),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_11_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__28832),
            .in2(_gnd_net_),
            .in3(N__28811),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_11_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__29012),
            .in2(_gnd_net_),
            .in3(N__28991),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_LC_11_11_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_LC_11_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__31696),
            .in2(_gnd_net_),
            .in3(N__28988),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8CZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_11_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__32075),
            .in2(_gnd_net_),
            .in3(N__28985),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_11_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__28982),
            .in2(_gnd_net_),
            .in3(N__28952),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_12_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__31574),
            .in2(_gnd_net_),
            .in3(N__28934),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_12_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__33671),
            .in2(_gnd_net_),
            .in3(N__28931),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_12_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__32192),
            .in2(_gnd_net_),
            .in3(N__28928),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_12_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__32065),
            .in2(_gnd_net_),
            .in3(N__28925),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_12_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_12_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29054),
            .in3(N__28922),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_12_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__32029),
            .in2(_gnd_net_),
            .in3(N__29078),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_12_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__29038),
            .in2(_gnd_net_),
            .in3(N__29075),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_15_LC_11_12_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_11_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_2_RNI_15_LC_11_12_7  (
            .in0(N__32030),
            .in1(N__32066),
            .in2(N__29039),
            .in3(N__29053),
            .lcout(\VPP_VDDQ.un9_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_13_LC_11_13_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_13_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_13_LC_11_13_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_13_LC_11_13_0  (
            .in0(N__33290),
            .in1(N__33465),
            .in2(N__33664),
            .in3(N__29071),
            .lcout(\VPP_VDDQ.count_2_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33136),
            .ce(N__32418),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_13_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_13_1  (
            .in0(N__29072),
            .in1(N__33654),
            .in2(N__33473),
            .in3(N__33293),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI98N41_13_LC_11_13_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI98N41_13_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI98N41_13_LC_11_13_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNI98N41_13_LC_11_13_2  (
            .in0(N__32381),
            .in1(_gnd_net_),
            .in2(N__29063),
            .in3(N__29060),
            .lcout(\VPP_VDDQ.count_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_13_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_13_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_13_4  (
            .in0(N__33655),
            .in1(N__33470),
            .in2(N__33299),
            .in3(N__29026),
            .lcout(),
            .ltout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIDEP41_15_LC_11_13_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIDEP41_15_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIDEP41_15_LC_11_13_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIDEP41_15_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__29018),
            .in2(N__29042),
            .in3(N__32382),
            .lcout(\VPP_VDDQ.count_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_15_LC_11_13_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_15_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_15_LC_11_13_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_15_LC_11_13_6  (
            .in0(N__33291),
            .in1(N__33466),
            .in2(N__33665),
            .in3(N__29027),
            .lcout(\VPP_VDDQ.count_2_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33136),
            .ce(N__32418),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_14_LC_11_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_14_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_14_LC_11_13_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_14_LC_11_13_7  (
            .in0(N__33464),
            .in1(N__33647),
            .in2(N__32056),
            .in3(N__33292),
            .lcout(\VPP_VDDQ.count_2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33136),
            .ce(N__32418),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_14_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_14_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_14_0  (
            .in0(N__29268),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29138),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_11_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_11_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_11_14_3  (
            .in0(N__31629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29267),
            .lcout(\VPP_VDDQ.N_360 ),
            .ltout(\VPP_VDDQ.N_360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_4 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__29620),
            .in2(N__29165),
            .in3(N__29681),
            .lcout(\VPP_VDDQ.N_264_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_14_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_14_5 .LUT_INIT=16'b0010110010101010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_14_5  (
            .in0(N__29137),
            .in1(N__29726),
            .in2(N__29624),
            .in3(N__29575),
            .lcout(),
            .ltout(\VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_14_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_14_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_14_6  (
            .in0(N__29576),
            .in1(N__29084),
            .in2(N__29141),
            .in3(N__29646),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33137),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNITROD7_0_LC_11_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNITROD7_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNITROD7_0_LC_11_15_0 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNITROD7_0_LC_11_15_0  (
            .in0(N__29725),
            .in1(N__29617),
            .in2(N__29714),
            .in3(N__29547),
            .lcout(\VPP_VDDQ.curr_state_RNITROD7Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_RNITROD7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_11_15_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_11_15_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_11_15_1  (
            .in0(N__29548),
            .in1(_gnd_net_),
            .in2(N__29096),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.N_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_15_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_15_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_15_2  (
            .in0(N__29675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29618),
            .lcout(\VPP_VDDQ.N_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_15_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__29673),
            .in2(_gnd_net_),
            .in3(N__29640),
            .lcout(\VPP_VDDQ.N_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_11_15_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_11_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.curr_state_RNI8I855_0_LC_11_15_4  (
            .in0(N__29674),
            .in1(N__29616),
            .in2(_gnd_net_),
            .in3(N__29704),
            .lcout(\VPP_VDDQ.N_214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_11_16_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_11_16_0 .LUT_INIT=16'b0000010010101110;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_11_16_0  (
            .in0(N__29680),
            .in1(N__29619),
            .in2(N__29651),
            .in3(N__29705),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33112),
            .ce(N__29416),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_11_16_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_11_16_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__29679),
            .in2(_gnd_net_),
            .in3(N__29650),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33112),
            .ce(N__29416),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIFMN39_12_LC_12_3_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIFMN39_12_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIFMN39_12_LC_12_3_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.count_off_RNIFMN39_12_LC_12_3_0  (
            .in0(N__29306),
            .in1(N__30911),
            .in2(N__29888),
            .in3(N__30775),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_1_LC_12_3_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_1_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_1_LC_12_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.count_off_RNI_1_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__29817),
            .in2(_gnd_net_),
            .in3(N__30066),
            .lcout(\POWERLED.count_off_RNIZ0Z_1 ),
            .ltout(\POWERLED.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIL3SN8_1_LC_12_3_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIL3SN8_1_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIL3SN8_1_LC_12_3_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.count_off_RNIL3SN8_1_LC_12_3_2  (
            .in0(N__29294),
            .in1(N__30912),
            .in2(N__29309),
            .in3(N__30776),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_12_3_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_12_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_12_3_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_12_LC_12_3_3  (
            .in0(N__30913),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29884),
            .lcout(\POWERLED.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33068),
            .ce(N__30783),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_12_3_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_1_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_12_3_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_1_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__29300),
            .in2(_gnd_net_),
            .in3(N__30915),
            .lcout(\POWERLED.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33068),
            .ce(N__30783),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_12_3_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_13_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_12_3_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_13_LC_12_3_5  (
            .in0(N__30914),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29857),
            .lcout(\POWERLED.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33068),
            .ce(N__30783),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHPO39_13_LC_12_3_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHPO39_13_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHPO39_13_LC_12_3_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.count_off_RNIHPO39_13_LC_12_3_6  (
            .in0(N__29840),
            .in1(N__30910),
            .in2(N__29861),
            .in3(N__30774),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(\POWERLED.count_offZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_15_LC_12_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_15_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_15_LC_12_3_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_15_LC_12_3_7  (
            .in0(N__30143),
            .in1(N__30065),
            .in2(N__29834),
            .in3(N__30199),
            .lcout(\POWERLED.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_12_4_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_12_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(N__29818),
            .in2(N__30068),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNIN70F_LC_12_4_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNIN70F_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNIN70F_LC_12_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNIN70F_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(N__29801),
            .in2(_gnd_net_),
            .in3(N__29786),
            .lcout(\POWERLED.un3_count_off_1_cry_1_c_RNIN70FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_1 ),
            .carryout(\POWERLED.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_12_4_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_12_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(N__30077),
            .in2(_gnd_net_),
            .in3(N__29783),
            .lcout(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_2 ),
            .carryout(\POWERLED.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_12_4_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_12_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_12_4_3  (
            .in0(_gnd_net_),
            .in1(N__30128),
            .in2(_gnd_net_),
            .in3(N__29780),
            .lcout(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_3 ),
            .carryout(\POWERLED.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNIQD3F_LC_12_4_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNIQD3F_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNIQD3F_LC_12_4_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un3_count_off_1_cry_4_c_RNIQD3F_LC_12_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29777),
            .in3(N__29750),
            .lcout(\POWERLED.un3_count_off_1_cry_4_c_RNIQD3FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_4 ),
            .carryout(\POWERLED.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNIRF4F_LC_12_4_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNIRF4F_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNIRF4F_LC_12_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNIRF4F_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(N__29747),
            .in2(_gnd_net_),
            .in3(N__29729),
            .lcout(\POWERLED.un3_count_off_1_cry_5_c_RNIRF4FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_5 ),
            .carryout(\POWERLED.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNISH5F_LC_12_4_6 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNISH5F_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNISH5F_LC_12_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNISH5F_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(N__30038),
            .in2(_gnd_net_),
            .in3(N__30023),
            .lcout(\POWERLED.un3_count_off_1_cry_6_c_RNISH5FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_6 ),
            .carryout(\POWERLED.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNITJ6F_LC_12_4_7 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNITJ6F_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNITJ6F_LC_12_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_7_c_RNITJ6F_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(N__30016),
            .in2(_gnd_net_),
            .in3(N__29996),
            .lcout(\POWERLED.un3_count_off_1_cry_7_c_RNITJ6FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_7 ),
            .carryout(\POWERLED.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIUL7F_LC_12_5_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIUL7F_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIUL7F_LC_12_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNIUL7F_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__29993),
            .in2(_gnd_net_),
            .in3(N__29966),
            .lcout(\POWERLED.un3_count_off_1_cry_8_c_RNIUL7FZ0 ),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIVN8F_LC_12_5_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIVN8F_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIVN8F_LC_12_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_9_c_RNIVN8F_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__29963),
            .in2(_gnd_net_),
            .in3(N__29930),
            .lcout(\POWERLED.un3_count_off_1_cry_9_c_RNIVN8FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_9 ),
            .carryout(\POWERLED.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNI7ULD_LC_12_5_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNI7ULD_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNI7ULD_LC_12_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNI7ULD_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__29927),
            .in2(_gnd_net_),
            .in3(N__29912),
            .lcout(\POWERLED.un3_count_off_1_cry_10_c_RNI7ULDZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_10 ),
            .carryout(\POWERLED.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNI80ND_LC_12_5_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNI80ND_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNI80ND_LC_12_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_11_c_RNI80ND_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__29905),
            .in2(_gnd_net_),
            .in3(N__29873),
            .lcout(\POWERLED.un3_count_off_1_cry_11_c_RNI80NDZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_11 ),
            .carryout(\POWERLED.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNI92OD_LC_12_5_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNI92OD_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNI92OD_LC_12_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_12_c_RNI92OD_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__29870),
            .in2(_gnd_net_),
            .in3(N__29846),
            .lcout(\POWERLED.un3_count_off_1_cry_12_c_RNI92ODZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_12 ),
            .carryout(\POWERLED.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIA4PD_LC_12_5_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIA4PD_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIA4PD_LC_12_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_13_c_RNIA4PD_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(N__30139),
            .in2(_gnd_net_),
            .in3(N__29843),
            .lcout(\POWERLED.un3_count_off_1_cry_13_c_RNIA4PDZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_13 ),
            .carryout(\POWERLED.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIB6QD_LC_12_5_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIB6QD_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIB6QD_LC_12_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un3_count_off_1_cry_14_c_RNIB6QD_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(N__30203),
            .in2(_gnd_net_),
            .in3(N__30188),
            .lcout(\POWERLED.un3_count_off_1_cry_14_c_RNIB6QDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJSP39_14_LC_12_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJSP39_14_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJSP39_14_LC_12_5_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.count_off_RNIJSP39_14_LC_12_5_7  (
            .in0(N__30173),
            .in1(N__30888),
            .in2(N__30161),
            .in3(N__30773),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_12_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_3_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_12_6_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_3_LC_12_6_0  (
            .in0(N__30862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30106),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33028),
            .ce(N__30788),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHIU69_4_LC_12_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHIU69_4_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHIU69_4_LC_12_6_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.count_off_RNIHIU69_4_LC_12_6_1  (
            .in0(N__30794),
            .in1(N__30859),
            .in2(N__30950),
            .in3(N__30756),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(\POWERLED.count_offZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIFFT69_0_3_LC_12_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIFFT69_0_3_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIFFT69_0_3_LC_12_6_2 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \POWERLED.count_off_RNIFFT69_0_3_LC_12_6_2  (
            .in0(N__30757),
            .in1(N__30095),
            .in2(N__30119),
            .in3(N__30086),
            .lcout(\POWERLED.un34_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIMIBQ2_LC_12_6_3 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIMIBQ2_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIMIBQ2_LC_12_6_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNIMIBQ2_LC_12_6_3  (
            .in0(N__30107),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30858),
            .lcout(\POWERLED.count_off_1_3 ),
            .ltout(\POWERLED.count_off_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIFFT69_3_LC_12_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIFFT69_3_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIFFT69_3_LC_12_6_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_off_RNIFFT69_3_LC_12_6_4  (
            .in0(N__30755),
            .in1(_gnd_net_),
            .in2(N__30089),
            .in3(N__30085),
            .lcout(\POWERLED.un3_count_off_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIK2SN8_0_LC_12_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIK2SN8_0_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIK2SN8_0_LC_12_6_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \POWERLED.count_off_RNIK2SN8_0_LC_12_6_5  (
            .in0(N__30956),
            .in1(N__30860),
            .in2(N__30067),
            .in3(N__30754),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(\POWERLED.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_12_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_12_6_6 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \POWERLED.count_off_0_LC_12_6_6  (
            .in0(N__30861),
            .in1(_gnd_net_),
            .in2(N__30959),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33028),
            .ce(N__30788),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_12_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_4_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_12_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_4_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__30946),
            .in2(_gnd_net_),
            .in3(N__30863),
            .lcout(\POWERLED.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33028),
            .ce(N__30788),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_3_LC_12_7_0 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_LC_12_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_LC_12_7_0  (
            .in0(N__30611),
            .in1(N__30599),
            .in2(N__30587),
            .in3(N__30428),
            .lcout(),
            .ltout(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_LC_12_7_1 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_LC_12_7_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__30398),
            .in2(N__30392),
            .in3(N__30389),
            .lcout(vccin_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_12_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_12_7_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_12_7_2  (
            .in0(N__30254),
            .in1(N__31659),
            .in2(N__30245),
            .in3(N__30230),
            .lcout(),
            .ltout(\VPP_VDDQ.delayed_vddq_okZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI9SRO4_LC_12_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI9SRO4_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI9SRO4_LC_12_7_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNI9SRO4_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30338),
            .in3(N__30328),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_12_7_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_12_7_5 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNINI731_0_LC_12_7_5  (
            .in0(N__30227),
            .in1(N__33661),
            .in2(N__31661),
            .in3(N__31801),
            .lcout(\VPP_VDDQ.delayed_vddq_ok_en ),
            .ltout(\VPP_VDDQ.delayed_vddq_ok_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_7_6 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_7_6 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_LC_12_7_6  (
            .in0(N__30241),
            .in1(N__31658),
            .in2(N__30248),
            .in3(N__30229),
            .lcout(\VPP_VDDQ.delayed_vddq_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33049),
            .ce(),
            .sr(N__30215));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_7_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_7_7  (
            .in0(N__30228),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.N_53_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIH136_11_LC_12_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIH136_11_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIH136_11_LC_12_8_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.count_clk_RNIH136_11_LC_12_8_0  (
            .in0(N__31394),
            .in1(N__31160),
            .in2(N__31409),
            .in3(N__31309),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_11_LC_12_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_11_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_12_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_clk_11_LC_12_8_1  (
            .in0(N__31311),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31405),
            .lcout(\POWERLED.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33051),
            .ce(N__31219),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_12_LC_12_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_12_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_12_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_12_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__31378),
            .in2(_gnd_net_),
            .in3(N__31313),
            .lcout(\POWERLED.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33051),
            .ce(N__31219),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIJ446_12_LC_12_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIJ446_12_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIJ446_12_LC_12_8_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \POWERLED.count_clk_RNIJ446_12_LC_12_8_3  (
            .in0(N__31310),
            .in1(N__31388),
            .in2(N__31382),
            .in3(N__31192),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_LC_12_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_12_8_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.count_clk_1_LC_12_8_4  (
            .in0(N__31348),
            .in1(N__31312),
            .in2(_gnd_net_),
            .in3(N__31077),
            .lcout(\POWERLED.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33051),
            .ce(N__31219),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIRG8B_1_LC_12_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIRG8B_1_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIRG8B_1_LC_12_8_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \POWERLED.count_clk_RNIRG8B_1_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__31229),
            .in2(N__31191),
            .in3(N__31091),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(\POWERLED.count_clkZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_LC_12_8_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_LC_12_8_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \POWERLED.count_clk_RNI_1_LC_12_8_6  (
            .in0(N__31052),
            .in1(N__31040),
            .in2(N__31007),
            .in3(N__31004),
            .lcout(\POWERLED.N_176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_9_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_9_0 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_9_0  (
            .in0(N__31599),
            .in1(N__33545),
            .in2(N__33450),
            .in3(N__33269),
            .lcout(),
            .ltout(\VPP_VDDQ.N_47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_12_9_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_12_9_1 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__31490),
            .in2(N__31544),
            .in3(N__32000),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_9_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_9_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_9_2  (
            .in0(N__33555),
            .in1(N__31540),
            .in2(N__31520),
            .in3(N__33270),
            .lcout(\VPP_VDDQ.count_2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_1_LC_12_9_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_1_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_1_LC_12_9_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \VPP_VDDQ.curr_state_2_1_LC_12_9_4  (
            .in0(N__33393),
            .in1(N__33547),
            .in2(N__31603),
            .in3(N__33273),
            .lcout(\VPP_VDDQ.curr_state_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33127),
            .ce(N__31772),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_12_9_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_12_9_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_12_9_5  (
            .in0(N__33271),
            .in1(N__33556),
            .in2(N__31483),
            .in3(N__33391),
            .lcout(\VPP_VDDQ.count_2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_12_9_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_12_9_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_12_9_6  (
            .in0(N__33392),
            .in1(N__33546),
            .in2(N__32285),
            .in3(N__33272),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI7EJU_3_LC_12_9_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI7EJU_3_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI7EJU_3_LC_12_9_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNI7EJU_3_LC_12_9_7  (
            .in0(N__32362),
            .in1(_gnd_net_),
            .in2(N__31451),
            .in3(N__32267),
            .lcout(\VPP_VDDQ.count_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_0_LC_12_10_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_0_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_0_LC_12_10_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \VPP_VDDQ.curr_state_2_0_LC_12_10_0  (
            .in0(N__31433),
            .in1(N__33615),
            .in2(N__31660),
            .in3(N__31677),
            .lcout(\VPP_VDDQ.curr_state_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33135),
            .ce(N__31771),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_12_10_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_12_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_12_10_1  (
            .in0(N__33429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33207),
            .lcout(\VPP_VDDQ.N_385 ),
            .ltout(\VPP_VDDQ.N_385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_12_10_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_12_10_2 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_12_10_2  (
            .in0(N__31653),
            .in1(N__33616),
            .in2(N__31427),
            .in3(N__31678),
            .lcout(),
            .ltout(\VPP_VDDQ.m4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_12_10_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_12_10_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__32018),
            .in2(N__32012),
            .in3(N__32009),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_12_10_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_12_10_4 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_12_10_4  (
            .in0(N__31595),
            .in1(N__31676),
            .in2(N__31805),
            .in3(N__31794),
            .lcout(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIDNMU_6_LC_12_10_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIDNMU_6_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIDNMU_6_LC_12_10_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIDNMU_6_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__31685),
            .in2(N__31706),
            .in3(N__32243),
            .lcout(\VPP_VDDQ.count_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_0_LC_12_10_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_0_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_0_LC_12_10_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNII8C7_0_LC_12_10_6  (
            .in0(N__33208),
            .in1(N__33430),
            .in2(N__32258),
            .in3(N__33617),
            .lcout(\VPP_VDDQ.count_2_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_a2_0_LC_12_10_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_a2_0_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_a2_0_LC_12_10_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_a2_0_LC_12_10_7  (
            .in0(N__31679),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31654),
            .lcout(N_362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_0_LC_12_11_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_12_11_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \VPP_VDDQ.count_2_RNI_0_LC_12_11_0  (
            .in0(N__33432),
            .in1(N__32137),
            .in2(N__33618),
            .in3(N__33236),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIL8AN_0_LC_12_11_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIL8AN_0_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIL8AN_0_LC_12_11_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIL8AN_0_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__32114),
            .in2(N__31577),
            .in3(N__32331),
            .lcout(\VPP_VDDQ.count_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_12_11_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_12_11_2 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_12_11_2  (
            .in0(N__32333),
            .in1(N__31573),
            .in2(N__32090),
            .in3(N__32096),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIQODG5_10_LC_12_11_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIQODG5_10_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIQODG5_10_LC_12_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIQODG5_10_LC_12_11_3  (
            .in0(N__32183),
            .in1(N__31559),
            .in2(N__31553),
            .in3(N__31550),
            .lcout(\VPP_VDDQ.N_1_i ),
            .ltout(\VPP_VDDQ.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_0_LC_12_11_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_0_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_0_LC_12_11_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \VPP_VDDQ.count_2_0_LC_12_11_4  (
            .in0(N__33434),
            .in1(N__33656),
            .in2(N__32153),
            .in3(N__32136),
            .lcout(\VPP_VDDQ.count_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33141),
            .ce(N__32403),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_7_LC_12_11_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_7_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_7_LC_12_11_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_7_LC_12_11_5  (
            .in0(N__33238),
            .in1(N__33554),
            .in2(N__32108),
            .in3(N__33435),
            .lcout(\VPP_VDDQ.count_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33141),
            .ce(N__32403),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_11_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_11_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_11_6  (
            .in0(N__33433),
            .in1(N__32104),
            .in2(N__33619),
            .in3(N__33237),
            .lcout(\VPP_VDDQ.count_2_1_7 ),
            .ltout(\VPP_VDDQ.count_2_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFQNU_7_LC_12_11_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFQNU_7_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFQNU_7_LC_12_11_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIFQNU_7_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__32086),
            .in2(N__32078),
            .in3(N__32332),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_12_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_12_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_12_0  (
            .in0(N__33241),
            .in1(N__33313),
            .in2(N__33662),
            .in3(N__33454),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI75M41_12_LC_12_12_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI75M41_12_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI75M41_12_LC_12_12_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI75M41_12_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__32380),
            .in2(N__32069),
            .in3(N__33152),
            .lcout(\VPP_VDDQ.count_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_12_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_12_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_12_2  (
            .in0(N__33240),
            .in1(N__33625),
            .in2(N__32057),
            .in3(N__33453),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIBBO41_14_LC_12_12_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIBBO41_14_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIBBO41_14_LC_12_12_3 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIBBO41_14_LC_12_12_3  (
            .in0(N__32039),
            .in1(N__32379),
            .in2(N__32033),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_3_LC_12_12_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_3_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_3_LC_12_12_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_3_LC_12_12_4  (
            .in0(N__33242),
            .in1(N__32281),
            .in2(N__33663),
            .in3(N__33456),
            .lcout(\VPP_VDDQ.count_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33111),
            .ce(N__32425),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_6_LC_12_12_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_6_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_6_LC_12_12_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.count_2_6_LC_12_12_5  (
            .in0(N__33455),
            .in1(N__33244),
            .in2(N__33659),
            .in3(N__32254),
            .lcout(\VPP_VDDQ.count_2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33111),
            .ce(N__32425),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_8_LC_12_12_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_8_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_8_LC_12_12_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_8_LC_12_12_6  (
            .in0(N__33243),
            .in1(N__33626),
            .in2(N__32219),
            .in3(N__33457),
            .lcout(\VPP_VDDQ.count_2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33111),
            .ce(N__32425),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_12_12_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_12_12_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_12_12_7  (
            .in0(N__33452),
            .in1(N__33239),
            .in2(N__33658),
            .in3(N__32218),
            .lcout(\VPP_VDDQ.count_2_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_10_LC_12_13_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_10_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_10_LC_12_13_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_10_LC_12_13_0  (
            .in0(N__33284),
            .in1(N__33703),
            .in2(N__33472),
            .in3(N__33634),
            .lcout(\VPP_VDDQ.count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33146),
            .ce(N__32409),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_13_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_13_1  (
            .in0(N__33631),
            .in1(N__33459),
            .in2(N__33298),
            .in3(N__32173),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI52L41_11_LC_12_13_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI52L41_11_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI52L41_11_LC_12_13_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI52L41_11_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__32159),
            .in2(N__32195),
            .in3(N__32377),
            .lcout(\VPP_VDDQ.count_2Z0Z_11 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIS3FU_0_10_LC_12_13_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIS3FU_0_10_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIS3FU_0_10_LC_12_13_3 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \VPP_VDDQ.count_2_RNIS3FU_0_10_LC_12_13_3  (
            .in0(N__32378),
            .in1(N__33686),
            .in2(N__32186),
            .in3(N__33692),
            .lcout(\VPP_VDDQ.un9_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_11_LC_12_13_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_11_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_11_LC_12_13_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_11_LC_12_13_4  (
            .in0(N__33285),
            .in1(N__33633),
            .in2(N__32174),
            .in3(N__33471),
            .lcout(\VPP_VDDQ.count_2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33146),
            .ce(N__32409),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_12_13_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_12_13_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_12_13_5  (
            .in0(N__33630),
            .in1(N__33458),
            .in2(N__33704),
            .in3(N__33283),
            .lcout(\VPP_VDDQ.count_2_1_10 ),
            .ltout(\VPP_VDDQ.count_2_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIS3FU_10_LC_12_13_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIS3FU_10_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIS3FU_10_LC_12_13_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIS3FU_10_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__33685),
            .in2(N__33674),
            .in3(N__32376),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_12_LC_12_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_12_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_12_LC_12_13_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_12_LC_12_13_7  (
            .in0(N__33632),
            .in1(N__33460),
            .in2(N__33314),
            .in3(N__33286),
            .lcout(\VPP_VDDQ.count_2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33146),
            .ce(N__32409),
            .sr(_gnd_net_));
endmodule // TOP
