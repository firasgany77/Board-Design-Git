-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 9 2022 14:41:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "pwrbtn_block" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of pwrbtn_block
entity pwrbtn_block is
port (
    rsmrst_n : in std_logic;
    pwrbtn : out std_logic;
    clk_100k : in std_logic);
end pwrbtn_block;

-- Architecture of pwrbtn_block
-- View name is \INTERFACE\
architecture \INTERFACE\ of pwrbtn_block is

signal \N__1865\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1856\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1827\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1810\ : std_logic;
signal \N__1807\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1801\ : std_logic;
signal \N__1798\ : std_logic;
signal \N__1795\ : std_logic;
signal \N__1792\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1785\ : std_logic;
signal \N__1784\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1775\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1753\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1719\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1716\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1711\ : std_logic;
signal \N__1708\ : std_logic;
signal \N__1701\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1694\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1685\ : std_logic;
signal \N__1682\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1655\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1632\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1630\ : std_logic;
signal \N__1629\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1618\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1604\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1601\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1546\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1534\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1525\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1512\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1509\ : std_logic;
signal \N__1506\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1501\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1465\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1443\ : std_logic;
signal \N__1440\ : std_logic;
signal \N__1437\ : std_logic;
signal \N__1432\ : std_logic;
signal \N__1431\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1429\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1426\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1408\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1402\ : std_logic;
signal \N__1401\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1398\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1393\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1385\ : std_logic;
signal \N__1380\ : std_logic;
signal \N__1373\ : std_logic;
signal \N__1370\ : std_logic;
signal \N__1357\ : std_logic;
signal \N__1354\ : std_logic;
signal \N__1353\ : std_logic;
signal \N__1352\ : std_logic;
signal \N__1351\ : std_logic;
signal \N__1348\ : std_logic;
signal \N__1347\ : std_logic;
signal \N__1346\ : std_logic;
signal \N__1345\ : std_logic;
signal \N__1344\ : std_logic;
signal \N__1343\ : std_logic;
signal \N__1340\ : std_logic;
signal \N__1339\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1333\ : std_logic;
signal \N__1330\ : std_logic;
signal \N__1321\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1319\ : std_logic;
signal \N__1318\ : std_logic;
signal \N__1317\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1307\ : std_logic;
signal \N__1300\ : std_logic;
signal \N__1293\ : std_logic;
signal \N__1288\ : std_logic;
signal \N__1285\ : std_logic;
signal \N__1278\ : std_logic;
signal \N__1277\ : std_logic;
signal \N__1276\ : std_logic;
signal \N__1275\ : std_logic;
signal \N__1272\ : std_logic;
signal \N__1269\ : std_logic;
signal \N__1262\ : std_logic;
signal \N__1255\ : std_logic;
signal \N__1254\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1250\ : std_logic;
signal \N__1247\ : std_logic;
signal \N__1244\ : std_logic;
signal \N__1241\ : std_logic;
signal \N__1234\ : std_logic;
signal \N__1233\ : std_logic;
signal \N__1232\ : std_logic;
signal \N__1229\ : std_logic;
signal \N__1226\ : std_logic;
signal \N__1223\ : std_logic;
signal \N__1216\ : std_logic;
signal \N__1213\ : std_logic;
signal \N__1210\ : std_logic;
signal \N__1207\ : std_logic;
signal \N__1204\ : std_logic;
signal \N__1201\ : std_logic;
signal \N__1200\ : std_logic;
signal \N__1197\ : std_logic;
signal \N__1196\ : std_logic;
signal \N__1193\ : std_logic;
signal \N__1190\ : std_logic;
signal \N__1187\ : std_logic;
signal \N__1180\ : std_logic;
signal \N__1177\ : std_logic;
signal \N__1174\ : std_logic;
signal \N__1171\ : std_logic;
signal \N__1168\ : std_logic;
signal \N__1165\ : std_logic;
signal \N__1162\ : std_logic;
signal \N__1159\ : std_logic;
signal \N__1156\ : std_logic;
signal \N__1153\ : std_logic;
signal \N__1150\ : std_logic;
signal \N__1147\ : std_logic;
signal \N__1144\ : std_logic;
signal \N__1141\ : std_logic;
signal \N__1138\ : std_logic;
signal \N__1135\ : std_logic;
signal \N__1132\ : std_logic;
signal \N__1131\ : std_logic;
signal \N__1130\ : std_logic;
signal \N__1125\ : std_logic;
signal \N__1122\ : std_logic;
signal \N__1117\ : std_logic;
signal \N__1116\ : std_logic;
signal \N__1113\ : std_logic;
signal \N__1110\ : std_logic;
signal \N__1107\ : std_logic;
signal \N__1106\ : std_logic;
signal \N__1101\ : std_logic;
signal \N__1098\ : std_logic;
signal \N__1093\ : std_logic;
signal \N__1092\ : std_logic;
signal \N__1091\ : std_logic;
signal \N__1086\ : std_logic;
signal \N__1083\ : std_logic;
signal \N__1078\ : std_logic;
signal \N__1075\ : std_logic;
signal \N__1072\ : std_logic;
signal \N__1071\ : std_logic;
signal \N__1068\ : std_logic;
signal \N__1067\ : std_logic;
signal \N__1066\ : std_logic;
signal \N__1063\ : std_logic;
signal \N__1060\ : std_logic;
signal \N__1057\ : std_logic;
signal \N__1054\ : std_logic;
signal \N__1045\ : std_logic;
signal \N__1044\ : std_logic;
signal \N__1041\ : std_logic;
signal \N__1040\ : std_logic;
signal \N__1037\ : std_logic;
signal \N__1036\ : std_logic;
signal \N__1033\ : std_logic;
signal \N__1026\ : std_logic;
signal \N__1021\ : std_logic;
signal \N__1020\ : std_logic;
signal \N__1017\ : std_logic;
signal \N__1014\ : std_logic;
signal \N__1009\ : std_logic;
signal \N__1006\ : std_logic;
signal \N__1003\ : std_logic;
signal \N__1000\ : std_logic;
signal \N__999\ : std_logic;
signal \N__998\ : std_logic;
signal \N__995\ : std_logic;
signal \N__992\ : std_logic;
signal \N__989\ : std_logic;
signal \N__982\ : std_logic;
signal \N__979\ : std_logic;
signal \N__976\ : std_logic;
signal \N__973\ : std_logic;
signal \N__970\ : std_logic;
signal \N__969\ : std_logic;
signal \N__966\ : std_logic;
signal \N__963\ : std_logic;
signal \N__962\ : std_logic;
signal \N__959\ : std_logic;
signal \N__956\ : std_logic;
signal \N__953\ : std_logic;
signal \N__946\ : std_logic;
signal \N__943\ : std_logic;
signal \N__940\ : std_logic;
signal \N__937\ : std_logic;
signal \N__934\ : std_logic;
signal \N__931\ : std_logic;
signal \N__928\ : std_logic;
signal \N__927\ : std_logic;
signal \N__926\ : std_logic;
signal \N__923\ : std_logic;
signal \N__920\ : std_logic;
signal \N__917\ : std_logic;
signal \N__910\ : std_logic;
signal \N__907\ : std_logic;
signal \N__904\ : std_logic;
signal \N__901\ : std_logic;
signal \N__898\ : std_logic;
signal \N__897\ : std_logic;
signal \N__896\ : std_logic;
signal \N__893\ : std_logic;
signal \N__890\ : std_logic;
signal \N__887\ : std_logic;
signal \N__880\ : std_logic;
signal \N__877\ : std_logic;
signal \N__874\ : std_logic;
signal \N__871\ : std_logic;
signal \N__868\ : std_logic;
signal \N__865\ : std_logic;
signal \N__862\ : std_logic;
signal \N__859\ : std_logic;
signal \N__856\ : std_logic;
signal \N__853\ : std_logic;
signal \N__850\ : std_logic;
signal \N__847\ : std_logic;
signal \N__844\ : std_logic;
signal \N__841\ : std_logic;
signal \N__838\ : std_logic;
signal \N__835\ : std_logic;
signal \N__832\ : std_logic;
signal \N__829\ : std_logic;
signal \N__826\ : std_logic;
signal \N__823\ : std_logic;
signal \N__822\ : std_logic;
signal \N__821\ : std_logic;
signal \N__814\ : std_logic;
signal \N__811\ : std_logic;
signal \N__808\ : std_logic;
signal \N__805\ : std_logic;
signal \N__802\ : std_logic;
signal \N__799\ : std_logic;
signal \N__796\ : std_logic;
signal \N__793\ : std_logic;
signal \N__790\ : std_logic;
signal \N__787\ : std_logic;
signal \N__784\ : std_logic;
signal \N__781\ : std_logic;
signal \N__778\ : std_logic;
signal \N__775\ : std_logic;
signal \N__774\ : std_logic;
signal \N__771\ : std_logic;
signal \N__768\ : std_logic;
signal \N__763\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \curr_state_1_cascade_\ : std_logic;
signal \curr_state_0_cascade_\ : std_logic;
signal pwrbtn_c : std_logic;
signal \count_1_1_cascade_\ : std_logic;
signal curr_state_1 : std_logic;
signal \G_23\ : std_logic;
signal \count_1_0_cascade_\ : std_logic;
signal \count_0_cascade_\ : std_logic;
signal \clk_100k_ibuf_RNIZ0Z_1\ : std_logic;
signal \count_1_15_cascade_\ : std_logic;
signal \count_1_8_cascade_\ : std_logic;
signal un8_clk_100k_11 : std_logic;
signal \un8_clk_100k_10_cascade_\ : std_logic;
signal \un8_clk_100k_cascade_\ : std_logic;
signal \count_1_2_cascade_\ : std_logic;
signal \count_2_cascade_\ : std_logic;
signal un8_clk_100k_9 : std_logic;
signal \count_1_12_cascade_\ : std_logic;
signal \count_1_5_cascade_\ : std_logic;
signal \count_1_9_cascade_\ : std_logic;
signal \count_1_11_cascade_\ : std_logic;
signal \count_1_14_cascade_\ : std_logic;
signal count_1_3 : std_logic;
signal \count_1_7_cascade_\ : std_logic;
signal count_1 : std_logic;
signal count_0 : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal count_2 : std_logic;
signal \un2_count_1_cry_1_c_RNIC3FCZ0\ : std_logic;
signal un2_count_1_cry_1 : std_logic;
signal count_3 : std_logic;
signal \un2_count_1_cry_2_c_RNID5GCZ0\ : std_logic;
signal un2_count_1_cry_2 : std_logic;
signal un2_count_1_cry_3 : std_logic;
signal count_5 : std_logic;
signal \un2_count_1_cry_4_c_RNIF9ICZ0\ : std_logic;
signal un2_count_1_cry_4 : std_logic;
signal un2_count_1_cry_5 : std_logic;
signal count_7 : std_logic;
signal \un2_count_1_cry_6_c_RNIHDKCZ0\ : std_logic;
signal un2_count_1_cry_6 : std_logic;
signal count_8 : std_logic;
signal \un2_count_1_cry_7_c_RNIIFLCZ0\ : std_logic;
signal un2_count_1_cry_7 : std_logic;
signal un2_count_1_cry_8 : std_logic;
signal count_9 : std_logic;
signal \un2_count_1_cry_8_c_RNIJHMCZ0\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal un2_count_1_cry_9 : std_logic;
signal count_11 : std_logic;
signal \un2_count_1_cry_10_c_RNISE0AZ0\ : std_logic;
signal un2_count_1_cry_10 : std_logic;
signal \un2_count_1_cry_11_c_RNITG1AZ0\ : std_logic;
signal un2_count_1_cry_11 : std_logic;
signal un2_count_1_cry_12 : std_logic;
signal \un2_count_1_cry_13_c_RNIVK3AZ0\ : std_logic;
signal un2_count_1_cry_13 : std_logic;
signal un2_count_1_cry_14 : std_logic;
signal \un2_count_1_cry_14_c_RNI0N4AZ0\ : std_logic;
signal count_15 : std_logic;
signal count_14 : std_logic;
signal count_12 : std_logic;
signal un8_clk_100k_8 : std_logic;
signal count_10 : std_logic;
signal \un2_count_1_cry_9_c_RNIKJNCZ0\ : std_logic;
signal count_1_10 : std_logic;
signal \un2_count_1_cry_12_c_RNIUI2AZ0\ : std_logic;
signal \count_1_13_cascade_\ : std_logic;
signal count_13 : std_logic;
signal \un2_count_1_cry_3_c_RNIE7HCZ0\ : std_logic;
signal \count_1_4_cascade_\ : std_logic;
signal count_4 : std_logic;
signal curr_state_0 : std_logic;
signal un8_clk_100k : std_logic;
signal \un2_count_1_cry_5_c_RNIGBJCZ0\ : std_logic;
signal rsmrst_n_c : std_logic;
signal un17_clk_100k_i : std_logic;
signal \count_1_6_cascade_\ : std_logic;
signal clk_100k_c : std_logic;
signal count_6 : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_100k_wire : std_logic;
signal rsmrst_n_wire : std_logic;
signal pwrbtn_wire : std_logic;

begin
    clk_100k_wire <= clk_100k;
    rsmrst_n_wire <= rsmrst_n;
    pwrbtn <= pwrbtn_wire;

    \clk_100k_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1865\,
            DIN => \N__1864\,
            DOUT => \N__1863\,
            PACKAGEPIN => clk_100k_wire
        );

    \clk_100k_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1865\,
            PADOUT => \N__1864\,
            PADIN => \N__1863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_100k_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \rsmrst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1856\,
            DIN => \N__1855\,
            DOUT => \N__1854\,
            PACKAGEPIN => rsmrst_n_wire
        );

    \rsmrst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1856\,
            PADOUT => \N__1855\,
            PADIN => \N__1854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => rsmrst_n_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwrbtn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1847\,
            DIN => \N__1846\,
            DOUT => \N__1845\,
            PACKAGEPIN => pwrbtn_wire
        );

    \pwrbtn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1847\,
            PADOUT => \N__1846\,
            PADIN => \N__1845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__781\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__421\ : InMux
    port map (
            O => \N__1828\,
            I => \N__1823\
        );

    \I__420\ : InMux
    port map (
            O => \N__1827\,
            I => \N__1820\
        );

    \I__419\ : InMux
    port map (
            O => \N__1826\,
            I => \N__1817\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__1823\,
            I => count_10
        );

    \I__417\ : LocalMux
    port map (
            O => \N__1820\,
            I => count_10
        );

    \I__416\ : LocalMux
    port map (
            O => \N__1817\,
            I => count_10
        );

    \I__415\ : InMux
    port map (
            O => \N__1810\,
            I => \N__1807\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__1807\,
            I => \un2_count_1_cry_9_c_RNIKJNCZ0\
        );

    \I__413\ : InMux
    port map (
            O => \N__1804\,
            I => \N__1801\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__1801\,
            I => count_1_10
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__1798\,
            I => \N__1795\
        );

    \I__410\ : InMux
    port map (
            O => \N__1795\,
            I => \N__1792\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__1792\,
            I => \un2_count_1_cry_12_c_RNIUI2AZ0\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__1789\,
            I => \count_1_13_cascade_\
        );

    \I__407\ : InMux
    port map (
            O => \N__1786\,
            I => \N__1781\
        );

    \I__406\ : InMux
    port map (
            O => \N__1785\,
            I => \N__1778\
        );

    \I__405\ : InMux
    port map (
            O => \N__1784\,
            I => \N__1775\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__1781\,
            I => count_13
        );

    \I__403\ : LocalMux
    port map (
            O => \N__1778\,
            I => count_13
        );

    \I__402\ : LocalMux
    port map (
            O => \N__1775\,
            I => count_13
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__1768\,
            I => \N__1765\
        );

    \I__400\ : InMux
    port map (
            O => \N__1765\,
            I => \N__1762\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__1762\,
            I => \N__1759\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__1759\,
            I => \un2_count_1_cry_3_c_RNIE7HCZ0\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__1756\,
            I => \count_1_4_cascade_\
        );

    \I__396\ : InMux
    port map (
            O => \N__1753\,
            I => \N__1749\
        );

    \I__395\ : InMux
    port map (
            O => \N__1752\,
            I => \N__1746\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__1749\,
            I => \N__1740\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__1746\,
            I => \N__1740\
        );

    \I__392\ : InMux
    port map (
            O => \N__1745\,
            I => \N__1737\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__1740\,
            I => count_4
        );

    \I__390\ : LocalMux
    port map (
            O => \N__1737\,
            I => count_4
        );

    \I__389\ : InMux
    port map (
            O => \N__1732\,
            I => \N__1720\
        );

    \I__388\ : InMux
    port map (
            O => \N__1731\,
            I => \N__1720\
        );

    \I__387\ : InMux
    port map (
            O => \N__1730\,
            I => \N__1720\
        );

    \I__386\ : InMux
    port map (
            O => \N__1729\,
            I => \N__1720\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__1720\,
            I => \N__1708\
        );

    \I__384\ : InMux
    port map (
            O => \N__1719\,
            I => \N__1701\
        );

    \I__383\ : InMux
    port map (
            O => \N__1718\,
            I => \N__1701\
        );

    \I__382\ : InMux
    port map (
            O => \N__1717\,
            I => \N__1701\
        );

    \I__381\ : InMux
    port map (
            O => \N__1716\,
            I => \N__1696\
        );

    \I__380\ : InMux
    port map (
            O => \N__1715\,
            I => \N__1696\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__1714\,
            I => \N__1690\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__1713\,
            I => \N__1686\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__1712\,
            I => \N__1682\
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__1711\,
            I => \N__1679\
        );

    \I__375\ : Span4Mux_v
    port map (
            O => \N__1708\,
            I => \N__1675\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__1701\,
            I => \N__1672\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__1696\,
            I => \N__1669\
        );

    \I__372\ : InMux
    port map (
            O => \N__1695\,
            I => \N__1662\
        );

    \I__371\ : InMux
    port map (
            O => \N__1694\,
            I => \N__1662\
        );

    \I__370\ : InMux
    port map (
            O => \N__1693\,
            I => \N__1662\
        );

    \I__369\ : InMux
    port map (
            O => \N__1690\,
            I => \N__1655\
        );

    \I__368\ : InMux
    port map (
            O => \N__1689\,
            I => \N__1655\
        );

    \I__367\ : InMux
    port map (
            O => \N__1686\,
            I => \N__1655\
        );

    \I__366\ : InMux
    port map (
            O => \N__1685\,
            I => \N__1646\
        );

    \I__365\ : InMux
    port map (
            O => \N__1682\,
            I => \N__1646\
        );

    \I__364\ : InMux
    port map (
            O => \N__1679\,
            I => \N__1646\
        );

    \I__363\ : InMux
    port map (
            O => \N__1678\,
            I => \N__1646\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__1675\,
            I => curr_state_0
        );

    \I__361\ : Odrv12
    port map (
            O => \N__1672\,
            I => curr_state_0
        );

    \I__360\ : Odrv4
    port map (
            O => \N__1669\,
            I => curr_state_0
        );

    \I__359\ : LocalMux
    port map (
            O => \N__1662\,
            I => curr_state_0
        );

    \I__358\ : LocalMux
    port map (
            O => \N__1655\,
            I => curr_state_0
        );

    \I__357\ : LocalMux
    port map (
            O => \N__1646\,
            I => curr_state_0
        );

    \I__356\ : InMux
    port map (
            O => \N__1633\,
            I => \N__1620\
        );

    \I__355\ : InMux
    port map (
            O => \N__1632\,
            I => \N__1620\
        );

    \I__354\ : InMux
    port map (
            O => \N__1631\,
            I => \N__1620\
        );

    \I__353\ : InMux
    port map (
            O => \N__1630\,
            I => \N__1609\
        );

    \I__352\ : InMux
    port map (
            O => \N__1629\,
            I => \N__1609\
        );

    \I__351\ : InMux
    port map (
            O => \N__1628\,
            I => \N__1609\
        );

    \I__350\ : CascadeMux
    port map (
            O => \N__1627\,
            I => \N__1606\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__1620\,
            I => \N__1597\
        );

    \I__348\ : InMux
    port map (
            O => \N__1619\,
            I => \N__1588\
        );

    \I__347\ : InMux
    port map (
            O => \N__1618\,
            I => \N__1588\
        );

    \I__346\ : InMux
    port map (
            O => \N__1617\,
            I => \N__1588\
        );

    \I__345\ : InMux
    port map (
            O => \N__1616\,
            I => \N__1588\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__1609\,
            I => \N__1585\
        );

    \I__343\ : InMux
    port map (
            O => \N__1606\,
            I => \N__1578\
        );

    \I__342\ : InMux
    port map (
            O => \N__1605\,
            I => \N__1578\
        );

    \I__341\ : InMux
    port map (
            O => \N__1604\,
            I => \N__1578\
        );

    \I__340\ : InMux
    port map (
            O => \N__1603\,
            I => \N__1571\
        );

    \I__339\ : InMux
    port map (
            O => \N__1602\,
            I => \N__1571\
        );

    \I__338\ : InMux
    port map (
            O => \N__1601\,
            I => \N__1571\
        );

    \I__337\ : InMux
    port map (
            O => \N__1600\,
            I => \N__1568\
        );

    \I__336\ : Odrv4
    port map (
            O => \N__1597\,
            I => un8_clk_100k
        );

    \I__335\ : LocalMux
    port map (
            O => \N__1588\,
            I => un8_clk_100k
        );

    \I__334\ : Odrv4
    port map (
            O => \N__1585\,
            I => un8_clk_100k
        );

    \I__333\ : LocalMux
    port map (
            O => \N__1578\,
            I => un8_clk_100k
        );

    \I__332\ : LocalMux
    port map (
            O => \N__1571\,
            I => un8_clk_100k
        );

    \I__331\ : LocalMux
    port map (
            O => \N__1568\,
            I => un8_clk_100k
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__1555\,
            I => \N__1552\
        );

    \I__329\ : InMux
    port map (
            O => \N__1552\,
            I => \N__1549\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__1549\,
            I => \N__1546\
        );

    \I__327\ : Odrv4
    port map (
            O => \N__1546\,
            I => \un2_count_1_cry_5_c_RNIGBJCZ0\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__1543\,
            I => \N__1537\
        );

    \I__325\ : InMux
    port map (
            O => \N__1542\,
            I => \N__1525\
        );

    \I__324\ : InMux
    port map (
            O => \N__1541\,
            I => \N__1525\
        );

    \I__323\ : InMux
    port map (
            O => \N__1540\,
            I => \N__1525\
        );

    \I__322\ : InMux
    port map (
            O => \N__1537\,
            I => \N__1520\
        );

    \I__321\ : InMux
    port map (
            O => \N__1536\,
            I => \N__1520\
        );

    \I__320\ : CascadeMux
    port map (
            O => \N__1535\,
            I => \N__1517\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__1534\,
            I => \N__1513\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__1533\,
            I => \N__1506\
        );

    \I__317\ : CascadeMux
    port map (
            O => \N__1532\,
            I => \N__1502\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1525\,
            I => \N__1495\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__1520\,
            I => \N__1495\
        );

    \I__314\ : InMux
    port map (
            O => \N__1517\,
            I => \N__1492\
        );

    \I__313\ : InMux
    port map (
            O => \N__1516\,
            I => \N__1487\
        );

    \I__312\ : InMux
    port map (
            O => \N__1513\,
            I => \N__1487\
        );

    \I__311\ : InMux
    port map (
            O => \N__1512\,
            I => \N__1482\
        );

    \I__310\ : InMux
    port map (
            O => \N__1511\,
            I => \N__1482\
        );

    \I__309\ : InMux
    port map (
            O => \N__1510\,
            I => \N__1477\
        );

    \I__308\ : InMux
    port map (
            O => \N__1509\,
            I => \N__1477\
        );

    \I__307\ : InMux
    port map (
            O => \N__1506\,
            I => \N__1474\
        );

    \I__306\ : InMux
    port map (
            O => \N__1505\,
            I => \N__1465\
        );

    \I__305\ : InMux
    port map (
            O => \N__1502\,
            I => \N__1465\
        );

    \I__304\ : InMux
    port map (
            O => \N__1501\,
            I => \N__1465\
        );

    \I__303\ : InMux
    port map (
            O => \N__1500\,
            I => \N__1465\
        );

    \I__302\ : Span4Mux_h
    port map (
            O => \N__1495\,
            I => \N__1458\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__1492\,
            I => \N__1458\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1487\,
            I => \N__1458\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1482\,
            I => \N__1451\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1477\,
            I => \N__1451\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1474\,
            I => \N__1451\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1465\,
            I => \N__1448\
        );

    \I__295\ : Span4Mux_v
    port map (
            O => \N__1458\,
            I => \N__1443\
        );

    \I__294\ : Span4Mux_v
    port map (
            O => \N__1451\,
            I => \N__1443\
        );

    \I__293\ : Span12Mux_v
    port map (
            O => \N__1448\,
            I => \N__1440\
        );

    \I__292\ : Span4Mux_v
    port map (
            O => \N__1443\,
            I => \N__1437\
        );

    \I__291\ : Odrv12
    port map (
            O => \N__1440\,
            I => rsmrst_n_c
        );

    \I__290\ : Odrv4
    port map (
            O => \N__1437\,
            I => rsmrst_n_c
        );

    \I__289\ : InMux
    port map (
            O => \N__1432\,
            I => \N__1415\
        );

    \I__288\ : InMux
    port map (
            O => \N__1431\,
            I => \N__1415\
        );

    \I__287\ : InMux
    port map (
            O => \N__1430\,
            I => \N__1415\
        );

    \I__286\ : InMux
    port map (
            O => \N__1429\,
            I => \N__1415\
        );

    \I__285\ : InMux
    port map (
            O => \N__1428\,
            I => \N__1408\
        );

    \I__284\ : InMux
    port map (
            O => \N__1427\,
            I => \N__1408\
        );

    \I__283\ : InMux
    port map (
            O => \N__1426\,
            I => \N__1408\
        );

    \I__282\ : InMux
    port map (
            O => \N__1425\,
            I => \N__1403\
        );

    \I__281\ : InMux
    port map (
            O => \N__1424\,
            I => \N__1403\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1415\,
            I => \N__1393\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1408\,
            I => \N__1388\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1403\,
            I => \N__1388\
        );

    \I__277\ : InMux
    port map (
            O => \N__1402\,
            I => \N__1385\
        );

    \I__276\ : InMux
    port map (
            O => \N__1401\,
            I => \N__1380\
        );

    \I__275\ : InMux
    port map (
            O => \N__1400\,
            I => \N__1380\
        );

    \I__274\ : InMux
    port map (
            O => \N__1399\,
            I => \N__1373\
        );

    \I__273\ : InMux
    port map (
            O => \N__1398\,
            I => \N__1373\
        );

    \I__272\ : InMux
    port map (
            O => \N__1397\,
            I => \N__1373\
        );

    \I__271\ : InMux
    port map (
            O => \N__1396\,
            I => \N__1370\
        );

    \I__270\ : Odrv4
    port map (
            O => \N__1393\,
            I => un17_clk_100k_i
        );

    \I__269\ : Odrv4
    port map (
            O => \N__1388\,
            I => un17_clk_100k_i
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1385\,
            I => un17_clk_100k_i
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1380\,
            I => un17_clk_100k_i
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1373\,
            I => un17_clk_100k_i
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1370\,
            I => un17_clk_100k_i
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__1357\,
            I => \count_1_6_cascade_\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__1354\,
            I => \N__1348\
        );

    \I__262\ : CascadeMux
    port map (
            O => \N__1353\,
            I => \N__1340\
        );

    \I__261\ : InMux
    port map (
            O => \N__1352\,
            I => \N__1333\
        );

    \I__260\ : InMux
    port map (
            O => \N__1351\,
            I => \N__1333\
        );

    \I__259\ : InMux
    port map (
            O => \N__1348\,
            I => \N__1330\
        );

    \I__258\ : InMux
    port map (
            O => \N__1347\,
            I => \N__1321\
        );

    \I__257\ : InMux
    port map (
            O => \N__1346\,
            I => \N__1321\
        );

    \I__256\ : InMux
    port map (
            O => \N__1345\,
            I => \N__1321\
        );

    \I__255\ : InMux
    port map (
            O => \N__1344\,
            I => \N__1321\
        );

    \I__254\ : InMux
    port map (
            O => \N__1343\,
            I => \N__1307\
        );

    \I__253\ : InMux
    port map (
            O => \N__1340\,
            I => \N__1307\
        );

    \I__252\ : InMux
    port map (
            O => \N__1339\,
            I => \N__1307\
        );

    \I__251\ : InMux
    port map (
            O => \N__1338\,
            I => \N__1307\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1333\,
            I => \N__1300\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1330\,
            I => \N__1300\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1321\,
            I => \N__1300\
        );

    \I__247\ : InMux
    port map (
            O => \N__1320\,
            I => \N__1293\
        );

    \I__246\ : InMux
    port map (
            O => \N__1319\,
            I => \N__1293\
        );

    \I__245\ : InMux
    port map (
            O => \N__1318\,
            I => \N__1293\
        );

    \I__244\ : InMux
    port map (
            O => \N__1317\,
            I => \N__1288\
        );

    \I__243\ : InMux
    port map (
            O => \N__1316\,
            I => \N__1288\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1307\,
            I => \N__1285\
        );

    \I__241\ : Span4Mux_h
    port map (
            O => \N__1300\,
            I => \N__1278\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__1293\,
            I => \N__1278\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1288\,
            I => \N__1278\
        );

    \I__238\ : Span4Mux_v
    port map (
            O => \N__1285\,
            I => \N__1272\
        );

    \I__237\ : Span4Mux_v
    port map (
            O => \N__1278\,
            I => \N__1269\
        );

    \I__236\ : InMux
    port map (
            O => \N__1277\,
            I => \N__1262\
        );

    \I__235\ : InMux
    port map (
            O => \N__1276\,
            I => \N__1262\
        );

    \I__234\ : InMux
    port map (
            O => \N__1275\,
            I => \N__1262\
        );

    \I__233\ : Odrv4
    port map (
            O => \N__1272\,
            I => clk_100k_c
        );

    \I__232\ : Odrv4
    port map (
            O => \N__1269\,
            I => clk_100k_c
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1262\,
            I => clk_100k_c
        );

    \I__230\ : InMux
    port map (
            O => \N__1255\,
            I => \N__1251\
        );

    \I__229\ : InMux
    port map (
            O => \N__1254\,
            I => \N__1247\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1251\,
            I => \N__1244\
        );

    \I__227\ : InMux
    port map (
            O => \N__1250\,
            I => \N__1241\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1247\,
            I => count_6
        );

    \I__225\ : Odrv4
    port map (
            O => \N__1244\,
            I => count_6
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1241\,
            I => count_6
        );

    \I__223\ : InMux
    port map (
            O => \N__1234\,
            I => \N__1229\
        );

    \I__222\ : InMux
    port map (
            O => \N__1233\,
            I => \N__1226\
        );

    \I__221\ : InMux
    port map (
            O => \N__1232\,
            I => \N__1223\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__1229\,
            I => count_9
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1226\,
            I => count_9
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1223\,
            I => count_9
        );

    \I__217\ : CascadeMux
    port map (
            O => \N__1216\,
            I => \N__1213\
        );

    \I__216\ : InMux
    port map (
            O => \N__1213\,
            I => \N__1210\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1210\,
            I => \un2_count_1_cry_8_c_RNIJHMCZ0\
        );

    \I__214\ : InMux
    port map (
            O => \N__1207\,
            I => \bfn_2_7_0_\
        );

    \I__213\ : InMux
    port map (
            O => \N__1204\,
            I => un2_count_1_cry_9
        );

    \I__212\ : CascadeMux
    port map (
            O => \N__1201\,
            I => \N__1197\
        );

    \I__211\ : InMux
    port map (
            O => \N__1200\,
            I => \N__1193\
        );

    \I__210\ : InMux
    port map (
            O => \N__1197\,
            I => \N__1190\
        );

    \I__209\ : InMux
    port map (
            O => \N__1196\,
            I => \N__1187\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1193\,
            I => count_11
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1190\,
            I => count_11
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1187\,
            I => count_11
        );

    \I__205\ : CascadeMux
    port map (
            O => \N__1180\,
            I => \N__1177\
        );

    \I__204\ : InMux
    port map (
            O => \N__1177\,
            I => \N__1174\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1174\,
            I => \un2_count_1_cry_10_c_RNISE0AZ0\
        );

    \I__202\ : InMux
    port map (
            O => \N__1171\,
            I => un2_count_1_cry_10
        );

    \I__201\ : CascadeMux
    port map (
            O => \N__1168\,
            I => \N__1165\
        );

    \I__200\ : InMux
    port map (
            O => \N__1165\,
            I => \N__1162\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1162\,
            I => \un2_count_1_cry_11_c_RNITG1AZ0\
        );

    \I__198\ : InMux
    port map (
            O => \N__1159\,
            I => un2_count_1_cry_11
        );

    \I__197\ : InMux
    port map (
            O => \N__1156\,
            I => un2_count_1_cry_12
        );

    \I__196\ : InMux
    port map (
            O => \N__1153\,
            I => \N__1150\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1150\,
            I => \N__1147\
        );

    \I__194\ : Odrv4
    port map (
            O => \N__1147\,
            I => \un2_count_1_cry_13_c_RNIVK3AZ0\
        );

    \I__193\ : InMux
    port map (
            O => \N__1144\,
            I => un2_count_1_cry_13
        );

    \I__192\ : InMux
    port map (
            O => \N__1141\,
            I => un2_count_1_cry_14
        );

    \I__191\ : InMux
    port map (
            O => \N__1138\,
            I => \N__1135\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1135\,
            I => \un2_count_1_cry_14_c_RNI0N4AZ0\
        );

    \I__189\ : InMux
    port map (
            O => \N__1132\,
            I => \N__1125\
        );

    \I__188\ : InMux
    port map (
            O => \N__1131\,
            I => \N__1125\
        );

    \I__187\ : InMux
    port map (
            O => \N__1130\,
            I => \N__1122\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1125\,
            I => count_15
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1122\,
            I => count_15
        );

    \I__184\ : CascadeMux
    port map (
            O => \N__1117\,
            I => \N__1113\
        );

    \I__183\ : InMux
    port map (
            O => \N__1116\,
            I => \N__1110\
        );

    \I__182\ : InMux
    port map (
            O => \N__1113\,
            I => \N__1107\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1110\,
            I => \N__1101\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1107\,
            I => \N__1101\
        );

    \I__179\ : InMux
    port map (
            O => \N__1106\,
            I => \N__1098\
        );

    \I__178\ : Odrv4
    port map (
            O => \N__1101\,
            I => count_14
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1098\,
            I => count_14
        );

    \I__176\ : InMux
    port map (
            O => \N__1093\,
            I => \N__1086\
        );

    \I__175\ : InMux
    port map (
            O => \N__1092\,
            I => \N__1086\
        );

    \I__174\ : InMux
    port map (
            O => \N__1091\,
            I => \N__1083\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1086\,
            I => count_12
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1083\,
            I => count_12
        );

    \I__171\ : InMux
    port map (
            O => \N__1078\,
            I => \N__1075\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1075\,
            I => un8_clk_100k_8
        );

    \I__169\ : InMux
    port map (
            O => \N__1072\,
            I => \N__1068\
        );

    \I__168\ : InMux
    port map (
            O => \N__1071\,
            I => \N__1063\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1068\,
            I => \N__1060\
        );

    \I__166\ : InMux
    port map (
            O => \N__1067\,
            I => \N__1057\
        );

    \I__165\ : InMux
    port map (
            O => \N__1066\,
            I => \N__1054\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1063\,
            I => count_1
        );

    \I__163\ : Odrv4
    port map (
            O => \N__1060\,
            I => count_1
        );

    \I__162\ : LocalMux
    port map (
            O => \N__1057\,
            I => count_1
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1054\,
            I => count_1
        );

    \I__160\ : CascadeMux
    port map (
            O => \N__1045\,
            I => \N__1041\
        );

    \I__159\ : CascadeMux
    port map (
            O => \N__1044\,
            I => \N__1037\
        );

    \I__158\ : InMux
    port map (
            O => \N__1041\,
            I => \N__1033\
        );

    \I__157\ : InMux
    port map (
            O => \N__1040\,
            I => \N__1026\
        );

    \I__156\ : InMux
    port map (
            O => \N__1037\,
            I => \N__1026\
        );

    \I__155\ : InMux
    port map (
            O => \N__1036\,
            I => \N__1026\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1033\,
            I => count_0
        );

    \I__153\ : LocalMux
    port map (
            O => \N__1026\,
            I => count_0
        );

    \I__152\ : InMux
    port map (
            O => \N__1021\,
            I => \N__1017\
        );

    \I__151\ : InMux
    port map (
            O => \N__1020\,
            I => \N__1014\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1017\,
            I => count_2
        );

    \I__149\ : LocalMux
    port map (
            O => \N__1014\,
            I => count_2
        );

    \I__148\ : InMux
    port map (
            O => \N__1009\,
            I => \N__1006\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1006\,
            I => \un2_count_1_cry_1_c_RNIC3FCZ0\
        );

    \I__146\ : InMux
    port map (
            O => \N__1003\,
            I => un2_count_1_cry_1
        );

    \I__145\ : InMux
    port map (
            O => \N__1000\,
            I => \N__995\
        );

    \I__144\ : InMux
    port map (
            O => \N__999\,
            I => \N__992\
        );

    \I__143\ : InMux
    port map (
            O => \N__998\,
            I => \N__989\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__995\,
            I => count_3
        );

    \I__141\ : LocalMux
    port map (
            O => \N__992\,
            I => count_3
        );

    \I__140\ : LocalMux
    port map (
            O => \N__989\,
            I => count_3
        );

    \I__139\ : InMux
    port map (
            O => \N__982\,
            I => \N__979\
        );

    \I__138\ : LocalMux
    port map (
            O => \N__979\,
            I => \un2_count_1_cry_2_c_RNID5GCZ0\
        );

    \I__137\ : InMux
    port map (
            O => \N__976\,
            I => un2_count_1_cry_2
        );

    \I__136\ : InMux
    port map (
            O => \N__973\,
            I => un2_count_1_cry_3
        );

    \I__135\ : InMux
    port map (
            O => \N__970\,
            I => \N__966\
        );

    \I__134\ : InMux
    port map (
            O => \N__969\,
            I => \N__963\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__966\,
            I => \N__959\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__963\,
            I => \N__956\
        );

    \I__131\ : InMux
    port map (
            O => \N__962\,
            I => \N__953\
        );

    \I__130\ : Odrv4
    port map (
            O => \N__959\,
            I => count_5
        );

    \I__129\ : Odrv4
    port map (
            O => \N__956\,
            I => count_5
        );

    \I__128\ : LocalMux
    port map (
            O => \N__953\,
            I => count_5
        );

    \I__127\ : InMux
    port map (
            O => \N__946\,
            I => \N__943\
        );

    \I__126\ : LocalMux
    port map (
            O => \N__943\,
            I => \N__940\
        );

    \I__125\ : Odrv4
    port map (
            O => \N__940\,
            I => \un2_count_1_cry_4_c_RNIF9ICZ0\
        );

    \I__124\ : InMux
    port map (
            O => \N__937\,
            I => un2_count_1_cry_4
        );

    \I__123\ : InMux
    port map (
            O => \N__934\,
            I => un2_count_1_cry_5
        );

    \I__122\ : InMux
    port map (
            O => \N__931\,
            I => \N__928\
        );

    \I__121\ : LocalMux
    port map (
            O => \N__928\,
            I => \N__923\
        );

    \I__120\ : InMux
    port map (
            O => \N__927\,
            I => \N__920\
        );

    \I__119\ : InMux
    port map (
            O => \N__926\,
            I => \N__917\
        );

    \I__118\ : Odrv4
    port map (
            O => \N__923\,
            I => count_7
        );

    \I__117\ : LocalMux
    port map (
            O => \N__920\,
            I => count_7
        );

    \I__116\ : LocalMux
    port map (
            O => \N__917\,
            I => count_7
        );

    \I__115\ : CascadeMux
    port map (
            O => \N__910\,
            I => \N__907\
        );

    \I__114\ : InMux
    port map (
            O => \N__907\,
            I => \N__904\
        );

    \I__113\ : LocalMux
    port map (
            O => \N__904\,
            I => \un2_count_1_cry_6_c_RNIHDKCZ0\
        );

    \I__112\ : InMux
    port map (
            O => \N__901\,
            I => un2_count_1_cry_6
        );

    \I__111\ : InMux
    port map (
            O => \N__898\,
            I => \N__893\
        );

    \I__110\ : InMux
    port map (
            O => \N__897\,
            I => \N__890\
        );

    \I__109\ : InMux
    port map (
            O => \N__896\,
            I => \N__887\
        );

    \I__108\ : LocalMux
    port map (
            O => \N__893\,
            I => count_8
        );

    \I__107\ : LocalMux
    port map (
            O => \N__890\,
            I => count_8
        );

    \I__106\ : LocalMux
    port map (
            O => \N__887\,
            I => count_8
        );

    \I__105\ : InMux
    port map (
            O => \N__880\,
            I => \N__877\
        );

    \I__104\ : LocalMux
    port map (
            O => \N__877\,
            I => \un2_count_1_cry_7_c_RNIIFLCZ0\
        );

    \I__103\ : InMux
    port map (
            O => \N__874\,
            I => un2_count_1_cry_7
        );

    \I__102\ : CascadeMux
    port map (
            O => \N__871\,
            I => \count_1_9_cascade_\
        );

    \I__101\ : CascadeMux
    port map (
            O => \N__868\,
            I => \count_1_11_cascade_\
        );

    \I__100\ : CascadeMux
    port map (
            O => \N__865\,
            I => \count_1_14_cascade_\
        );

    \I__99\ : InMux
    port map (
            O => \N__862\,
            I => \N__859\
        );

    \I__98\ : LocalMux
    port map (
            O => \N__859\,
            I => count_1_3
        );

    \I__97\ : CascadeMux
    port map (
            O => \N__856\,
            I => \count_1_7_cascade_\
        );

    \I__96\ : InMux
    port map (
            O => \N__853\,
            I => \N__850\
        );

    \I__95\ : LocalMux
    port map (
            O => \N__850\,
            I => un8_clk_100k_11
        );

    \I__94\ : CascadeMux
    port map (
            O => \N__847\,
            I => \un8_clk_100k_10_cascade_\
        );

    \I__93\ : CascadeMux
    port map (
            O => \N__844\,
            I => \un8_clk_100k_cascade_\
        );

    \I__92\ : CascadeMux
    port map (
            O => \N__841\,
            I => \count_1_2_cascade_\
        );

    \I__91\ : CascadeMux
    port map (
            O => \N__838\,
            I => \count_2_cascade_\
        );

    \I__90\ : InMux
    port map (
            O => \N__835\,
            I => \N__832\
        );

    \I__89\ : LocalMux
    port map (
            O => \N__832\,
            I => un8_clk_100k_9
        );

    \I__88\ : CascadeMux
    port map (
            O => \N__829\,
            I => \count_1_12_cascade_\
        );

    \I__87\ : CascadeMux
    port map (
            O => \N__826\,
            I => \count_1_5_cascade_\
        );

    \I__86\ : InMux
    port map (
            O => \N__823\,
            I => \N__814\
        );

    \I__85\ : InMux
    port map (
            O => \N__822\,
            I => \N__814\
        );

    \I__84\ : InMux
    port map (
            O => \N__821\,
            I => \N__814\
        );

    \I__83\ : LocalMux
    port map (
            O => \N__814\,
            I => curr_state_1
        );

    \I__82\ : InMux
    port map (
            O => \N__811\,
            I => \N__808\
        );

    \I__81\ : LocalMux
    port map (
            O => \N__808\,
            I => \G_23\
        );

    \I__80\ : CascadeMux
    port map (
            O => \N__805\,
            I => \count_1_0_cascade_\
        );

    \I__79\ : CascadeMux
    port map (
            O => \N__802\,
            I => \count_0_cascade_\
        );

    \I__78\ : InMux
    port map (
            O => \N__799\,
            I => \N__796\
        );

    \I__77\ : LocalMux
    port map (
            O => \N__796\,
            I => \clk_100k_ibuf_RNIZ0Z_1\
        );

    \I__76\ : CascadeMux
    port map (
            O => \N__793\,
            I => \count_1_15_cascade_\
        );

    \I__75\ : CascadeMux
    port map (
            O => \N__790\,
            I => \count_1_8_cascade_\
        );

    \I__74\ : CascadeMux
    port map (
            O => \N__787\,
            I => \curr_state_1_cascade_\
        );

    \I__73\ : CascadeMux
    port map (
            O => \N__784\,
            I => \curr_state_0_cascade_\
        );

    \I__72\ : IoInMux
    port map (
            O => \N__781\,
            I => \N__778\
        );

    \I__71\ : LocalMux
    port map (
            O => \N__778\,
            I => \N__775\
        );

    \I__70\ : IoSpan4Mux
    port map (
            O => \N__775\,
            I => \N__771\
        );

    \I__69\ : InMux
    port map (
            O => \N__774\,
            I => \N__768\
        );

    \I__68\ : Odrv4
    port map (
            O => \N__771\,
            I => pwrbtn_c
        );

    \I__67\ : LocalMux
    port map (
            O => \N__768\,
            I => pwrbtn_c
        );

    \I__66\ : CascadeMux
    port map (
            O => \N__763\,
            I => \count_1_1_cascade_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_count_1_cry_8,
            carryinitout => \bfn_2_7_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIQGTD_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__1347\,
            in1 => \N__811\,
            in2 => \_gnd_net_\,
            in3 => \N__821\,
            lcout => curr_state_1,
            ltout => \curr_state_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIQGTD_0_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010101010"
        )
    port map (
            in0 => \N__1678\,
            in1 => \N__1628\,
            in2 => \N__787\,
            in3 => \N__1345\,
            lcout => curr_state_0,
            ltout => \curr_state_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIQGTD_1_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__1346\,
            in1 => \_gnd_net_\,
            in2 => \N__784\,
            in3 => \N__774\,
            lcout => pwrbtn_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI_0_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__822\,
            in1 => \_gnd_net_\,
            in2 => \N__1711\,
            in3 => \_gnd_net_\,
            lcout => un17_clk_100k_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNITC49_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__1630\,
            in1 => \N__1685\,
            in2 => \N__1543\,
            in3 => \N__799\,
            lcout => OPEN,
            ltout => \count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNINT1N_0_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__1066\,
            in1 => \N__1396\,
            in2 => \N__763\,
            in3 => \N__1344\,
            lcout => count_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \curr_state_8_1_0__m4_0_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101001000000"
        )
    port map (
            in0 => \N__823\,
            in1 => \N__1629\,
            in2 => \N__1712\,
            in3 => \N__1536\,
            lcout => \G_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNITC49_0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__1516\,
            in1 => \N__1695\,
            in2 => \N__1627\,
            in3 => \N__1040\,
            lcout => OPEN,
            ltout => \count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNINT1N_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__1036\,
            in1 => \N__1320\,
            in2 => \N__805\,
            in3 => \N__1402\,
            lcout => count_0,
            ltout => \count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI_1_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__1067\,
            in1 => \_gnd_net_\,
            in2 => \N__802\,
            in3 => \_gnd_net_\,
            lcout => \clk_100k_ibuf_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIT39J_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__1694\,
            in1 => \N__1605\,
            in2 => \N__1535\,
            in3 => \N__1138\,
            lcout => OPEN,
            ltout => \count_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNINK611_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1319\,
            in1 => \N__1401\,
            in2 => \N__793\,
            in3 => \N__1130\,
            lcout => count_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI_4_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__969\,
            in1 => \N__1000\,
            in2 => \N__1044\,
            in3 => \N__1753\,
            lcout => un8_clk_100k_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIFSPL_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__1604\,
            in1 => \N__1693\,
            in2 => \N__1534\,
            in3 => \N__880\,
            lcout => OPEN,
            ltout => \count_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI9DN31_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1400\,
            in1 => \N__1318\,
            in2 => \N__790\,
            in3 => \N__896\,
            lcout => count_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI_3_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1233\,
            in1 => \N__897\,
            in2 => \N__1201\,
            in3 => \N__931\,
            lcout => OPEN,
            ltout => \un8_clk_100k_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI_5_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__853\,
            in1 => \N__835\,
            in2 => \N__847\,
            in3 => \N__1078\,
            lcout => un8_clk_100k,
            ltout => \un8_clk_100k_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNI9GJL_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__1511\,
            in1 => \N__1009\,
            in2 => \N__844\,
            in3 => \N__1715\,
            lcout => OPEN,
            ltout => \count_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI31H31_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1316\,
            in1 => \N__1424\,
            in2 => \N__841\,
            in3 => \N__1020\,
            lcout => count_2,
            ltout => \count_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI_2_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1072\,
            in1 => \N__1254\,
            in2 => \N__838\,
            in3 => \N__1828\,
            lcout => un8_clk_100k_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIQT5J_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__1716\,
            in1 => \N__1600\,
            in2 => \N__1168\,
            in3 => \N__1512\,
            lcout => OPEN,
            ltout => \count_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIKE311_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__1425\,
            in1 => \N__1091\,
            in2 => \N__829\,
            in3 => \N__1317\,
            lcout => count_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNICMML_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__1717\,
            in1 => \N__1601\,
            in2 => \N__1533\,
            in3 => \N__946\,
            lcout => OPEN,
            ltout => \count_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI67K31_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__962\,
            in1 => \N__1426\,
            in2 => \N__826\,
            in3 => \N__1275\,
            lcout => count_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIGUQL_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__1718\,
            in1 => \N__1602\,
            in2 => \N__1216\,
            in3 => \N__1509\,
            lcout => OPEN,
            ltout => \count_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIAFO31_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__1232\,
            in1 => \N__1427\,
            in2 => \N__871\,
            in3 => \N__1276\,
            lcout => count_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIPR4J_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__1719\,
            in1 => \N__1603\,
            in2 => \N__1180\,
            in3 => \N__1510\,
            lcout => OPEN,
            ltout => \count_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIJC211_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__1196\,
            in1 => \N__1428\,
            in2 => \N__868\,
            in3 => \N__1277\,
            lcout => count_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIS18J_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__1633\,
            in1 => \N__1153\,
            in2 => \N__1714\,
            in3 => \N__1542\,
            lcout => OPEN,
            ltout => \count_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIMI511_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1352\,
            in1 => \N__1399\,
            in2 => \N__865\,
            in3 => \N__1106\,
            lcout => count_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIAIKL_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__1631\,
            in1 => \N__982\,
            in2 => \N__1713\,
            in3 => \N__1540\,
            lcout => count_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI43I31_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__1397\,
            in1 => \N__998\,
            in2 => \N__1354\,
            in3 => \N__862\,
            lcout => count_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIEQOL_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__1541\,
            in1 => \N__1632\,
            in2 => \N__910\,
            in3 => \N__1689\,
            lcout => OPEN,
            ltout => \count_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI8BM31_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1398\,
            in1 => \N__1351\,
            in2 => \N__856\,
            in3 => \N__926\,
            lcout => count_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_1_c_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1071\,
            in2 => \N__1045\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => un2_count_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_1_c_RNIC3FC_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1021\,
            in2 => \_gnd_net_\,
            in3 => \N__1003\,
            lcout => \un2_count_1_cry_1_c_RNIC3FCZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_1,
            carryout => un2_count_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_2_c_RNID5GC_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__999\,
            in2 => \_gnd_net_\,
            in3 => \N__976\,
            lcout => \un2_count_1_cry_2_c_RNID5GCZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_2,
            carryout => un2_count_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_3_c_RNIE7HC_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1752\,
            in2 => \_gnd_net_\,
            in3 => \N__973\,
            lcout => \un2_count_1_cry_3_c_RNIE7HCZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_3,
            carryout => un2_count_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_4_c_RNIF9IC_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__970\,
            in2 => \_gnd_net_\,
            in3 => \N__937\,
            lcout => \un2_count_1_cry_4_c_RNIF9ICZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_4,
            carryout => un2_count_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_5_c_RNIGBJC_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1255\,
            in2 => \_gnd_net_\,
            in3 => \N__934\,
            lcout => \un2_count_1_cry_5_c_RNIGBJCZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_5,
            carryout => un2_count_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_6_c_RNIHDKC_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__927\,
            in2 => \_gnd_net_\,
            in3 => \N__901\,
            lcout => \un2_count_1_cry_6_c_RNIHDKCZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_6,
            carryout => un2_count_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_7_c_RNIIFLC_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__898\,
            in2 => \_gnd_net_\,
            in3 => \N__874\,
            lcout => \un2_count_1_cry_7_c_RNIIFLCZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_7,
            carryout => un2_count_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_8_c_RNIJHMC_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1234\,
            in2 => \_gnd_net_\,
            in3 => \N__1207\,
            lcout => \un2_count_1_cry_8_c_RNIJHMCZ0\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => un2_count_1_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_9_c_RNIKJNC_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1827\,
            in2 => \_gnd_net_\,
            in3 => \N__1204\,
            lcout => \un2_count_1_cry_9_c_RNIKJNCZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_9,
            carryout => un2_count_1_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_10_c_RNISE0A_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1200\,
            in2 => \_gnd_net_\,
            in3 => \N__1171\,
            lcout => \un2_count_1_cry_10_c_RNISE0AZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_10,
            carryout => un2_count_1_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_11_c_RNITG1A_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1093\,
            in2 => \_gnd_net_\,
            in3 => \N__1159\,
            lcout => \un2_count_1_cry_11_c_RNITG1AZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_11,
            carryout => un2_count_1_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_12_c_RNIUI2A_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1786\,
            in2 => \_gnd_net_\,
            in3 => \N__1156\,
            lcout => \un2_count_1_cry_12_c_RNIUI2AZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_12,
            carryout => un2_count_1_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_13_c_RNIVK3A_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1116\,
            in2 => \_gnd_net_\,
            in3 => \N__1144\,
            lcout => \un2_count_1_cry_13_c_RNIVK3AZ0\,
            ltout => OPEN,
            carryin => un2_count_1_cry_13,
            carryout => un2_count_1_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_count_1_cry_14_c_RNI0N4A_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1132\,
            in2 => \_gnd_net_\,
            in3 => \N__1141\,
            lcout => \un2_count_1_cry_14_c_RNI0N4AZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1131\,
            in1 => \N__1785\,
            in2 => \N__1117\,
            in3 => \N__1092\,
            lcout => un8_clk_100k_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNIBHP31_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__1431\,
            in1 => \N__1804\,
            in2 => \N__1353\,
            in3 => \N__1826\,
            lcout => count_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIH0SL_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__1618\,
            in1 => \N__1810\,
            in2 => \N__1532\,
            in3 => \N__1731\,
            lcout => count_1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIRV6J_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__1732\,
            in1 => \N__1619\,
            in2 => \N__1798\,
            in3 => \N__1505\,
            lcout => OPEN,
            ltout => \count_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNILG411_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__1784\,
            in1 => \N__1432\,
            in2 => \N__1789\,
            in3 => \N__1343\,
            lcout => count_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIBKLL_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__1729\,
            in1 => \N__1616\,
            in2 => \N__1768\,
            in3 => \N__1500\,
            lcout => OPEN,
            ltout => \count_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI55J31_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__1745\,
            in1 => \N__1429\,
            in2 => \N__1756\,
            in3 => \N__1338\,
            lcout => count_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rsmrst_n_ibuf_RNIDONL_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__1730\,
            in1 => \N__1617\,
            in2 => \N__1555\,
            in3 => \N__1501\,
            lcout => OPEN,
            ltout => \count_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_100k_ibuf_RNI79L31_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__1250\,
            in1 => \N__1430\,
            in2 => \N__1357\,
            in3 => \N__1339\,
            lcout => count_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
