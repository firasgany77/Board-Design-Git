-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 24 2022 21:31:32

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : in std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : in std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : in std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__37287\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \b2v_inst16.count_rst_12_cascade_\ : std_logic;
signal \b2v_inst16.count_rst_13_cascade_\ : std_logic;
signal \b2v_inst16.count_rst_14_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst16.count_4_9\ : std_logic;
signal \b2v_inst16.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst16.count_4_1\ : std_logic;
signal \b2v_inst16.count_4_11\ : std_logic;
signal \b2v_inst16.count_rst_0_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst16.count_4_8\ : std_logic;
signal \b2v_inst16.count_4_6\ : std_logic;
signal \b2v_inst16.count_4_15\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_1_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_16\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_0\ : std_logic;
signal \b2v_inst200.count_RNIZ0Z_1\ : std_logic;
signal \b2v_inst200.count_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_1_cascade_\ : std_logic;
signal \b2v_inst200.count_3_1\ : std_logic;
signal \b2v_inst200.count_3_2\ : std_logic;
signal \b2v_inst200.count_3_4\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_1\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \b2v_inst200.countZ0Z_2\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_5_cZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_16\ : std_logic;
signal \b2v_inst200.count_1_16\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_15\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.count_0_8\ : std_logic;
signal \b2v_inst11.count_0_9\ : std_logic;
signal \b2v_inst11.count_0_10\ : std_logic;
signal \b2v_inst11.count_0_11\ : std_logic;
signal \b2v_inst11.count_1_1_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_0_1\ : std_logic;
signal \b2v_inst11.count_0_2\ : std_logic;
signal \b2v_inst11.count_0_12\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \b2v_inst11.count_1_2\ : std_logic;
signal \b2v_inst11.un1_count_cry_1_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_cry_2\ : std_logic;
signal \b2v_inst11.un1_count_cry_3\ : std_logic;
signal \b2v_inst11.un1_count_cry_4\ : std_logic;
signal \b2v_inst11.un1_count_cry_5\ : std_logic;
signal \b2v_inst11.un1_count_cry_6\ : std_logic;
signal \b2v_inst11.count_1_8\ : std_logic;
signal \b2v_inst11.un1_count_cry_7\ : std_logic;
signal \b2v_inst11.un1_count_cry_8\ : std_logic;
signal \b2v_inst11.count_1_9\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \b2v_inst11.count_1_10\ : std_logic;
signal \b2v_inst11.un1_count_cry_9\ : std_logic;
signal \b2v_inst11.count_1_11\ : std_logic;
signal \b2v_inst11.un1_count_cry_10\ : std_logic;
signal \b2v_inst11.count_1_12\ : std_logic;
signal \b2v_inst11.un1_count_cry_11\ : std_logic;
signal \b2v_inst11.un1_count_cry_12\ : std_logic;
signal \b2v_inst11.un1_count_cry_13\ : std_logic;
signal \b2v_inst11.un1_count_cry_14\ : std_logic;
signal \b2v_inst16.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst16.count_4_4\ : std_logic;
signal \b2v_inst16.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst16.count_4_5\ : std_logic;
signal \b2v_inst16.count_4_7\ : std_logic;
signal \b2v_inst16.countZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst16.count_4_i_a3_8_0\ : std_logic;
signal \b2v_inst16.count_4_i_a3_9_0_cascade_\ : std_logic;
signal \b2v_inst16.count_4_i_a3_7_0\ : std_logic;
signal \b2v_inst16.count_rst_5\ : std_logic;
signal \b2v_inst16.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst16.N_414\ : std_logic;
signal \b2v_inst16.count_4_0\ : std_logic;
signal \b2v_inst16.count_4_2\ : std_logic;
signal \b2v_inst16.countZ0Z_0\ : std_logic;
signal \b2v_inst16.countZ0Z_1\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \b2v_inst16.un4_count_1_axb_2\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_1_c_RNIAGMEZ0\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_1\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_2\ : std_logic;
signal \b2v_inst16.countZ0Z_4\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_3\ : std_logic;
signal \b2v_inst16.countZ0Z_5\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_4\ : std_logic;
signal \b2v_inst16.countZ0Z_6\ : std_logic;
signal \b2v_inst16.count_rst_11\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_5\ : std_logic;
signal \b2v_inst16.countZ0Z_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_6\ : std_logic;
signal \b2v_inst16.countZ0Z_8\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_8\ : std_logic;
signal \b2v_inst16.countZ0Z_9\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_9\ : std_logic;
signal \b2v_inst16.countZ0Z_11\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_10\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_11\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_12\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_13\ : std_logic;
signal \b2v_inst16.countZ0Z_15\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_14\ : std_logic;
signal \b2v_inst16.count_rst_4\ : std_logic;
signal \b2v_inst200.count_3_14\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\ : std_logic;
signal \b2v_inst200.count_3_6\ : std_logic;
signal \b2v_inst200.count_1_6\ : std_logic;
signal \b2v_inst200.count_3_7\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\ : std_logic;
signal \b2v_inst200.count_0_17\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\ : std_logic;
signal \b2v_inst200.countZ0Z_17\ : std_logic;
signal \b2v_inst200.count_1_10\ : std_logic;
signal \b2v_inst200.count_3_10\ : std_logic;
signal \b2v_inst200.count_1_0\ : std_logic;
signal \b2v_inst200.countZ0Z_10\ : std_logic;
signal \b2v_inst200.count_1_8\ : std_logic;
signal \b2v_inst200.count_3_8\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_8\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_15\ : std_logic;
signal \b2v_inst200.count_3_15\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71\ : std_logic;
signal \b2v_inst200.countZ0Z_6\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_7\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_13\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_6_cascade_\ : std_logic;
signal \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_0\ : std_logic;
signal \b2v_inst200.count_3_0\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_9\ : std_logic;
signal \b2v_inst200.count_3_12\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\ : std_logic;
signal \b2v_inst200.countZ0Z_12\ : std_logic;
signal \b2v_inst200.count_3_9\ : std_logic;
signal \b2v_inst200.countZ0Z_12_cascade_\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_5\ : std_logic;
signal \b2v_inst200.count_3_11\ : std_logic;
signal \b2v_inst200.count_1_11\ : std_logic;
signal \b2v_inst200.countZ0Z_11\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_3\ : std_logic;
signal \b2v_inst200.countZ0Z_14\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_4\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_5_cascade_\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_14\ : std_logic;
signal \b2v_inst200.count_3_3\ : std_logic;
signal \b2v_inst200.countZ0Z_4\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_2\ : std_logic;
signal \b2v_inst200.count_3_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\ : std_logic;
signal \b2v_inst200.count_3_5\ : std_logic;
signal \b2v_inst200.countZ0Z_7\ : std_logic;
signal \b2v_inst200.count_en_g\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_3\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i_0_8\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_i_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_s_8\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_s_8\ : std_logic;
signal pwrbtn_led : std_logic;
signal \b2v_inst11.curr_state_3_0_cascade_\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_0_sqmuxa_i\ : std_logic;
signal \b2v_inst11.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \b2v_inst11.count_1_0_cascade_\ : std_logic;
signal \b2v_inst11.count_0_0\ : std_logic;
signal \b2v_inst11.pwm_outZ0\ : std_logic;
signal \b2v_inst11.g0_i_o3_0\ : std_logic;
signal \b2v_inst11.count_1_3\ : std_logic;
signal \b2v_inst11.count_0_3\ : std_logic;
signal \b2v_inst11.count_1_13\ : std_logic;
signal \b2v_inst11.count_0_13\ : std_logic;
signal \b2v_inst11.count_1_4\ : std_logic;
signal \b2v_inst11.count_0_4\ : std_logic;
signal \b2v_inst11.count_1_5\ : std_logic;
signal \b2v_inst11.count_0_5\ : std_logic;
signal \b2v_inst11.pwm_out_1_sqmuxa\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlt6_cascade_\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_3\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.N_8\ : std_logic;
signal \b2v_inst11.count_1_14\ : std_logic;
signal \b2v_inst11.count_0_14\ : std_logic;
signal \b2v_inst11.count_1_6\ : std_logic;
signal \b2v_inst11.count_0_6\ : std_logic;
signal \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\ : std_logic;
signal \b2v_inst11.count_0_15\ : std_logic;
signal \b2v_inst11.count_1_7\ : std_logic;
signal \b2v_inst11.count_0_7\ : std_logic;
signal \b2v_inst200.count_enZ0\ : std_logic;
signal pch_pwrok : std_logic;
signal vpp_en : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgd_eZ0Z_0\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgd_en\ : std_logic;
signal \b2v_inst16.N_26\ : std_logic;
signal \b2v_inst16.N_416\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst16.N_26_cascade_\ : std_logic;
signal \b2v_inst16.count_4_i_a3_10_0\ : std_logic;
signal \b2v_inst16.countZ0Z_14\ : std_logic;
signal \b2v_inst16.count_rst_3\ : std_logic;
signal \b2v_inst16.count_4_14\ : std_logic;
signal \b2v_inst16.countZ0Z_12\ : std_logic;
signal \b2v_inst16.count_rst_1\ : std_logic;
signal \b2v_inst16.count_4_12\ : std_logic;
signal \b2v_inst16.countZ0Z_13\ : std_logic;
signal \b2v_inst16.count_rst_2\ : std_logic;
signal \b2v_inst16.count_4_13\ : std_logic;
signal \b2v_inst16.N_3079_i\ : std_logic;
signal \b2v_inst16.count_4_3\ : std_logic;
signal \b2v_inst16.count_rst_8\ : std_logic;
signal \b2v_inst16.countZ0Z_3\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_7\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_3_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_7_1_cascade_\ : std_logic;
signal \b2v_inst16.curr_state_2_1\ : std_logic;
signal \b2v_inst16.curr_state_7_0_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_0_2_cascade_\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_a2_1_4\ : std_logic;
signal \b2v_inst11.N_355_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_55_1_tz\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_11_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_50_a0_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_50_a0_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_12_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_4_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_4_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_9Z0Z_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_46_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_11_1_0\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_l_fx_3\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \b2v_inst11.mult1_un54_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_s_8\ : std_logic;
signal \b2v_inst11.countZ0Z_0\ : std_logic;
signal \b2v_inst11.N_5980_i\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \b2v_inst11.countZ0Z_1\ : std_logic;
signal \b2v_inst11.N_5981_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_0\ : std_logic;
signal \b2v_inst11.countZ0Z_2\ : std_logic;
signal \b2v_inst11.N_5982_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_1\ : std_logic;
signal \b2v_inst11.countZ0Z_3\ : std_logic;
signal \b2v_inst11.N_5983_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_2\ : std_logic;
signal \b2v_inst11.countZ0Z_4\ : std_logic;
signal \b2v_inst11.N_5984_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_3\ : std_logic;
signal \b2v_inst11.countZ0Z_5\ : std_logic;
signal \b2v_inst11.N_5985_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_4\ : std_logic;
signal \b2v_inst11.countZ0Z_6\ : std_logic;
signal \b2v_inst11.N_5986_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_5\ : std_logic;
signal \b2v_inst11.countZ0Z_7\ : std_logic;
signal \b2v_inst11.N_5987_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_6\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_7\ : std_logic;
signal \b2v_inst11.countZ0Z_8\ : std_logic;
signal \b2v_inst11.N_5988_i\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \b2v_inst11.countZ0Z_9\ : std_logic;
signal \b2v_inst11.N_5989_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i_8\ : std_logic;
signal \b2v_inst11.countZ0Z_10\ : std_logic;
signal \b2v_inst11.N_5990_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_9\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i_8\ : std_logic;
signal \b2v_inst11.countZ0Z_11\ : std_logic;
signal \b2v_inst11.N_5991_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_10\ : std_logic;
signal \b2v_inst11.countZ0Z_12\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5992_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_11\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i_8\ : std_logic;
signal \b2v_inst11.countZ0Z_13\ : std_logic;
signal \b2v_inst11.N_5993_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_12\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i_8\ : std_logic;
signal \b2v_inst11.countZ0Z_14\ : std_logic;
signal \b2v_inst11.N_5994_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_13\ : std_logic;
signal \b2v_inst11.countZ0Z_15\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5995_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_14\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i_8\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_0\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2814\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_5\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0\ : std_logic;
signal \b2v_inst200.N_58_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst200.N_56\ : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \b2v_inst200.m6_i_0\ : std_logic;
signal \N_411\ : std_logic;
signal \b2v_inst200.m6_i_0_cascade_\ : std_logic;
signal \b2v_inst200.count_RNI5RUP8Z0Z_8\ : std_logic;
signal \b2v_inst200.curr_state_3_0\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_2\ : std_logic;
signal \b2v_inst200.i4_mux_cascade_\ : std_logic;
signal \b2v_inst200.curr_state_i_2_cascade_\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \b2v_inst200.N_3031_i\ : std_logic;
signal \b2v_inst200.N_205\ : std_logic;
signal \b2v_inst200.curr_state_i_2\ : std_logic;
signal \b2v_inst200.N_205_cascade_\ : std_logic;
signal \b2v_inst200.HDA_SDO_ATP_0\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst200.N_282\ : std_logic;
signal \b2v_inst200.curr_state_3_1\ : std_logic;
signal \b2v_inst16.curr_state_2_0\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \b2v_inst20.un4_counter_0\ : std_logic;
signal \b2v_inst20.un4_counter_2_and\ : std_logic;
signal \b2v_inst20.un4_counter_1\ : std_logic;
signal \b2v_inst20.un4_counter_3_and\ : std_logic;
signal \b2v_inst20.un4_counter_2\ : std_logic;
signal \b2v_inst20.un4_counter_4_and\ : std_logic;
signal \b2v_inst20.un4_counter_3\ : std_logic;
signal \b2v_inst20.un4_counter_5_and\ : std_logic;
signal \b2v_inst20.un4_counter_4\ : std_logic;
signal \b2v_inst20.un4_counter_5\ : std_logic;
signal \b2v_inst20.un4_counter_6\ : std_logic;
signal b2v_inst20_un4_counter_7 : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_11_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_39_0_1_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_7\ : std_logic;
signal \b2v_inst20.un4_counter_6_and\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_39_d_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNITSFK3Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_10\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNITSFK3Z0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_30_a1_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_5_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_6\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_9_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_8Z0Z_6\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_l_fx_6\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_i\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_12\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_8\ : std_logic;
signal \b2v_inst11.curr_state_4_0\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_s_4_sf\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_5\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_5_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_s_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_i_29\ : std_logic;
signal \b2v_inst16.count_rst\ : std_logic;
signal \b2v_inst16.count_4_10\ : std_logic;
signal \b2v_inst16.count_en\ : std_logic;
signal \b2v_inst16.countZ0Z_10\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i_8\ : std_logic;
signal vccst_en : std_logic;
signal \b2v_inst11.un85_clk_100khz_4\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i_8\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_2\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i_8\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_3\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i_8\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_s_8_cascade_\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_7_l_fx\ : std_logic;
signal \b2v_inst11.g3_0\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_axb_6\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_s_7\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_i\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_1\ : std_logic;
signal \b2v_inst20.counter_1_cry_2\ : std_logic;
signal \b2v_inst20.counter_1_cry_3\ : std_logic;
signal \b2v_inst20.counter_1_cry_4\ : std_logic;
signal \b2v_inst20.counter_1_cry_5\ : std_logic;
signal \b2v_inst20.counter_1_cry_6\ : std_logic;
signal \b2v_inst20.counterZ0Z_8\ : std_logic;
signal \b2v_inst20.counter_1_cry_7\ : std_logic;
signal \b2v_inst20.counter_1_cry_8\ : std_logic;
signal \b2v_inst20.counterZ0Z_9\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \b2v_inst20.counterZ0Z_10\ : std_logic;
signal \b2v_inst20.counter_1_cry_9\ : std_logic;
signal \b2v_inst20.counterZ0Z_11\ : std_logic;
signal \b2v_inst20.counter_1_cry_10\ : std_logic;
signal \b2v_inst20.counterZ0Z_12\ : std_logic;
signal \b2v_inst20.counter_1_cry_11\ : std_logic;
signal \b2v_inst20.counterZ0Z_13\ : std_logic;
signal \b2v_inst20.counter_1_cry_12\ : std_logic;
signal \b2v_inst20.counterZ0Z_14\ : std_logic;
signal \b2v_inst20.counter_1_cry_13\ : std_logic;
signal \b2v_inst20.counterZ0Z_15\ : std_logic;
signal \b2v_inst20.counter_1_cry_14\ : std_logic;
signal \b2v_inst20.counterZ0Z_16\ : std_logic;
signal \b2v_inst20.counter_1_cry_15\ : std_logic;
signal \b2v_inst20.counter_1_cry_16\ : std_logic;
signal \b2v_inst20.counterZ0Z_17\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \b2v_inst20.counterZ0Z_18\ : std_logic;
signal \b2v_inst20.counter_1_cry_17\ : std_logic;
signal \b2v_inst20.counterZ0Z_19\ : std_logic;
signal \b2v_inst20.counter_1_cry_18\ : std_logic;
signal \b2v_inst20.counterZ0Z_20\ : std_logic;
signal \b2v_inst20.counter_1_cry_19\ : std_logic;
signal \b2v_inst20.counterZ0Z_21\ : std_logic;
signal \b2v_inst20.counter_1_cry_20\ : std_logic;
signal \b2v_inst20.counterZ0Z_22\ : std_logic;
signal \b2v_inst20.counter_1_cry_21\ : std_logic;
signal \b2v_inst20.counterZ0Z_23\ : std_logic;
signal \b2v_inst20.counter_1_cry_22\ : std_logic;
signal \b2v_inst20.counterZ0Z_24\ : std_logic;
signal \b2v_inst20.counter_1_cry_23\ : std_logic;
signal \b2v_inst20.counter_1_cry_24\ : std_logic;
signal \b2v_inst20.counterZ0Z_25\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \b2v_inst20.counterZ0Z_26\ : std_logic;
signal \b2v_inst20.counter_1_cry_25\ : std_logic;
signal \b2v_inst20.counterZ0Z_27\ : std_logic;
signal \b2v_inst20.counter_1_cry_26\ : std_logic;
signal \b2v_inst20.counter_1_cry_27\ : std_logic;
signal \b2v_inst20.counter_1_cry_28\ : std_logic;
signal \b2v_inst20.counter_1_cry_29\ : std_logic;
signal \b2v_inst20.counter_1_cry_30\ : std_logic;
signal \b2v_inst20.counterZ0Z_28\ : std_logic;
signal \b2v_inst20.counterZ0Z_29\ : std_logic;
signal \b2v_inst20.counterZ0Z_30\ : std_logic;
signal \b2v_inst20.counterZ0Z_31\ : std_logic;
signal \b2v_inst20.un4_counter_7_and\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_9_1_1\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_5_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_8\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_3_0_tz\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.N_26_i_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_9_1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_13\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_4\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_8Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_4_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_8_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_3_1_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_3_cascade_\ : std_logic;
signal \b2v_inst11.un1_i3_mux_cascade_\ : std_logic;
signal \b2v_inst11.d_i3_mux\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_2\ : std_logic;
signal \b2v_inst11.mult1_un124_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_2\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_5\ : std_logic;
signal \b2v_inst11.mult1_un117_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_3\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_7\ : std_logic;
signal \b2v_inst11.mult1_un110_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_5\ : std_logic;
signal \b2v_inst11.mult1_un103_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_10\ : std_logic;
signal \b2v_inst11.mult1_un96_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_11\ : std_logic;
signal \b2v_inst11.mult1_un89_sum\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_12\ : std_logic;
signal \b2v_inst11.mult1_un82_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_13\ : std_logic;
signal \b2v_inst11.mult1_un75_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \b2v_inst11.mult1_un68_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_15\ : std_logic;
signal \b2v_inst11.mult1_un61_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_13\ : std_logic;
signal \b2v_inst11.mult1_un54_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_12\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \b2v_inst11.mult1_un47_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \b2v_inst11.CO2\ : std_logic;
signal \b2v_inst11.CO2_THRU_CO\ : std_logic;
signal \b2v_inst11.mult1_un131_sum\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_14\ : std_logic;
signal \b2v_inst5.count_1_6\ : std_logic;
signal vr_ready_vccinaux : std_logic;
signal vr_ready_vccin : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_4_l_fx\ : std_logic;
signal \b2v_inst11.mult1_un138_sum\ : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_2_c\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3_c\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4_c\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5_c\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6_c\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_s_8_cascade_\ : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_s_8_cascade_\ : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_axb_7\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i_0_8\ : std_logic;
signal \b2v_inst36.count_rst_3_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst36.count_2_11\ : std_logic;
signal \b2v_inst36.count_2_1\ : std_logic;
signal \b2v_inst36.count_2_15\ : std_logic;
signal \b2v_inst36.count_2_13\ : std_logic;
signal \b2v_inst36.count_2_14\ : std_logic;
signal \b2v_inst36.count_i_0\ : std_logic;
signal \b2v_inst5.count_1_7\ : std_logic;
signal \b2v_inst5.count_1_11\ : std_logic;
signal \b2v_inst5.countZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst5.count_1_12\ : std_logic;
signal \b2v_inst20.counterZ0Z_7\ : std_logic;
signal \b2v_inst20.un4_counter_1_and\ : std_logic;
signal \b2v_inst20.counter_1_cry_5_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_6\ : std_logic;
signal \b2v_inst20.counterZ0Z_1\ : std_logic;
signal \b2v_inst20.counterZ0Z_0\ : std_logic;
signal \b2v_inst20.un4_counter_0_and\ : std_logic;
signal \b2v_inst20.counter_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_5\ : std_logic;
signal \b2v_inst20.counter_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_4\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_0\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst5.count_rst_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst5.countZ0Z_7\ : std_logic;
signal \b2v_inst5.count_rst_7\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_11\ : std_logic;
signal \b2v_inst5.count_rst_3\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_14\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9JZ0Z1\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJZ0Z1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJZ0Z1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_3\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_3_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_0_3\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_40_and_i_0_0_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIT35D7Z0Z_4\ : std_logic;
signal \b2v_inst11.N_155_N\ : std_logic;
signal \b2v_inst11.dutycycle_en_11_cascade_\ : std_logic;
signal \b2v_inst11.N_158_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIT35D7Z0Z_15\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\ : std_logic;
signal \b2v_inst11.dutycycle_RNIT35D7Z0Z_15_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_15\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_14\ : std_logic;
signal \b2v_inst11.dutycycle_en_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_12\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_12_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_13\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19\ : std_logic;
signal \b2v_inst11.dutycycle_set_1_cascade_\ : std_logic;
signal \b2v_inst11.N_300\ : std_logic;
signal \b2v_inst11.N_300_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29\ : std_logic;
signal \b2v_inst11.dutycycle_set_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_set_0_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_0_6\ : std_logic;
signal \b2v_inst11.dutycycle_0_5\ : std_logic;
signal \b2v_inst11.dutycycle_set_1\ : std_logic;
signal \b2v_inst11.dutycycle_eena_13_0\ : std_logic;
signal \b2v_inst11.N_200_i_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_3\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_5\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_32_and_i_0_c\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_40_and_i_0_c\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_3\ : std_logic;
signal \b2v_inst11.mult1_un145_sum\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i\ : std_logic;
signal \b2v_inst11.N_10\ : std_logic;
signal \b2v_inst11.count_clk_0_8\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\ : std_logic;
signal \b2v_inst11.N_379\ : std_logic;
signal \b2v_inst11.N_379_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_9\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.N_190\ : std_logic;
signal \b2v_inst11.count_clk_0_5\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_1\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_15_cascade_\ : std_logic;
signal \b2v_inst11.N_175\ : std_logic;
signal \b2v_inst11.count_clk_0_14\ : std_logic;
signal \b2v_inst11.count_clk_0_15\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_3_cascade_\ : std_logic;
signal \b2v_inst36.count_rst_11\ : std_logic;
signal \b2v_inst36.count_rst_11_cascade_\ : std_logic;
signal \b2v_inst36.count_2_3\ : std_logic;
signal \b2v_inst36.count_rst_12_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst36.count_2_2\ : std_logic;
signal \b2v_inst36.count_rst_7_cascade_\ : std_logic;
signal \b2v_inst36.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst36.count_2_5\ : std_logic;
signal \b2v_inst36.count_2_7\ : std_logic;
signal \b2v_inst36.count_rst_7\ : std_logic;
signal \b2v_inst36.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst36.count_2_0\ : std_logic;
signal \b2v_inst36.count_rst_14\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_0\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_1\ : std_logic;
signal \b2v_inst36.count_rst_13\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_0\ : std_logic;
signal \b2v_inst36.countZ0Z_2\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_3\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst36.countZ0Z_5\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_7\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst36.countZ0Z_11\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst36.countZ0Z_13\ : std_logic;
signal \b2v_inst36.count_rst_1\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst36.countZ0Z_14\ : std_logic;
signal \b2v_inst36.count_rst_0\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst36.countZ0Z_15\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst36.count_rst\ : std_logic;
signal \b2v_inst20.counter_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_2\ : std_logic;
signal \b2v_inst36.curr_state_RNI3E27Z0Z_0_cascade_\ : std_logic;
signal dsw_pwrok : std_logic;
signal \b2v_inst20_un4_counter_7_THRU_CO\ : std_logic;
signal \b2v_inst20.counter_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_3\ : std_logic;
signal \b2v_inst5.countZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst5.count_1_13\ : std_logic;
signal \b2v_inst5.count_i_0_cascade_\ : std_logic;
signal \b2v_inst5.count_rst_14\ : std_logic;
signal \b2v_inst5.count_1_0\ : std_logic;
signal \b2v_inst5.count_rst_14_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_0\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2\ : std_logic;
signal \b2v_inst5.count_1_14\ : std_logic;
signal \b2v_inst5.countZ0Z_14\ : std_logic;
signal \b2v_inst5.count_i_0\ : std_logic;
signal \b2v_inst5.countZ0Z_14_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_12\ : std_logic;
signal \b2v_inst5.count_rst_6\ : std_logic;
signal \b2v_inst5.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_8_cascade_\ : std_logic;
signal \b2v_inst5.count_1_8\ : std_logic;
signal \b2v_inst5.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_4\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst5.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst5.count_1_4\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12_THRU_CO\ : std_logic;
signal \b2v_inst5.count_rst_1\ : std_logic;
signal \b2v_inst11.N_396_N_cascade_\ : std_logic;
signal \b2v_inst11.N_234_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_9\ : std_logic;
signal \b2v_inst11.dutycycle_rst_8\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_12\ : std_logic;
signal \b2v_inst11.dutycycle_eena_9_cascade_\ : std_logic;
signal \b2v_inst11.N_234_N\ : std_logic;
signal \b2v_inst11.dutycycle_eena_7\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_eena_7_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUFZ0Z1\ : std_logic;
signal \b2v_inst11.dutycycle_RNIT35D7Z0Z_13\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_11\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_5\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_6\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_9\ : std_logic;
signal \b2v_inst11.N_365_cascade_\ : std_logic;
signal \b2v_inst11.N_366_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_8\ : std_logic;
signal \b2v_inst11.N_153_N\ : std_logic;
signal \b2v_inst11.g2_i_a6_0\ : std_logic;
signal \b2v_inst11.N_363\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\ : std_logic;
signal \b2v_inst11.func_state_RNIDUQ02Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf0_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf1\ : std_logic;
signal \b2v_inst11.N_14_0_cascade_\ : std_logic;
signal \b2v_inst11.g2_i_2\ : std_logic;
signal \b2v_inst11.func_state_RNI_6Z0Z_0\ : std_logic;
signal \b2v_inst11.N_395_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.g0_4_2\ : std_logic;
signal \b2v_inst11.g0_0_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_36_and_i_o3_0_c_0\ : std_logic;
signal \b2v_inst11.g0_0_0_1\ : std_logic;
signal \b2v_inst11.func_state_RNI8H551Z0Z_0\ : std_logic;
signal \b2v_inst11.func_state_RNIDUQ02Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_eena_5_d_1_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_5_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_36_and_i_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI2IQ6CZ0Z_7\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_en_0\ : std_logic;
signal \b2v_inst11.N_328_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.count_clk_en_cascade_\ : std_logic;
signal \b2v_inst11.N_218\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_329_N_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_0\ : std_logic;
signal \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_2\ : std_logic;
signal \b2v_inst11.count_clk_0_3\ : std_logic;
signal \b2v_inst11.count_clk_0_4\ : std_logic;
signal \b2v_inst11.count_clk_0_6\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_2\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_3\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_6\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_8\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_9\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_9_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_10\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_11\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_12\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_14\ : std_logic;
signal \b2v_inst11.count_clk_1_14\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_13\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_15\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_14\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\ : std_logic;
signal \b2v_inst11.count_clk_0_11\ : std_logic;
signal \b2v_inst11.count_clk_1_11\ : std_logic;
signal \b2v_inst36.curr_state_7_0_cascade_\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.curr_state_0_0\ : std_logic;
signal \b2v_inst36.curr_state_0_1\ : std_logic;
signal \b2v_inst36.curr_state_7_1\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst36.DSW_PWROK_0\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst36.count_2_8\ : std_logic;
signal \b2v_inst36.count_rst_6\ : std_logic;
signal \b2v_inst36.countZ0Z_8\ : std_logic;
signal \b2v_inst36.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_5\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_4\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_6_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_7\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_9\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_13_cascade_\ : std_logic;
signal \b2v_inst36.N_1_i_cascade_\ : std_logic;
signal \b2v_inst36.count_rst_4\ : std_logic;
signal \b2v_inst36.count_rst_4_cascade_\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_10_cascade_\ : std_logic;
signal \b2v_inst36.N_1_i\ : std_logic;
signal \b2v_inst36.count_2_10\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_6\ : std_logic;
signal \b2v_inst36.count_rst_10\ : std_logic;
signal \b2v_inst36.count_2_4\ : std_logic;
signal \b2v_inst36.countZ0Z_4\ : std_logic;
signal \b2v_inst36.count_rst_8\ : std_logic;
signal \b2v_inst36.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst36.count_2_6\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_0\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_12\ : std_logic;
signal \b2v_inst36.count_2_12\ : std_logic;
signal \b2v_inst36.count_rst_2\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_1\ : std_logic;
signal \b2v_inst5.count_rst_13\ : std_logic;
signal \b2v_inst5.count_1_1\ : std_logic;
signal \b2v_inst5.count_rst_12\ : std_logic;
signal \b2v_inst5.count_1_2\ : std_logic;
signal \b2v_inst5.count_rst_11\ : std_logic;
signal \b2v_inst5.count_1_3\ : std_logic;
signal \b2v_inst5.countZ0Z_3\ : std_logic;
signal \b2v_inst5.countZ0Z_13\ : std_logic;
signal \b2v_inst5.countZ0Z_1\ : std_logic;
signal \b2v_inst5.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_2\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_11\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_4\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_5_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_10_cascade_\ : std_logic;
signal \b2v_inst5.count_1_10\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_1\ : std_logic;
signal \b2v_inst5.countZ0Z_5\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_9\ : std_logic;
signal \b2v_inst5.countZ0Z_6\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_12\ : std_logic;
signal \b2v_inst5.countZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst5.count_1_9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_10\ : std_logic;
signal \b2v_inst5.count_rst_4\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst5.curr_state_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_15\ : std_logic;
signal \b2v_inst5.count_rst\ : std_logic;
signal \b2v_inst5.count_1_15\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst5.countZ0Z_9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst5.N_1_i\ : std_logic;
signal \b2v_inst5.count_rst_5\ : std_logic;
signal \b2v_inst5.count_rst_9\ : std_logic;
signal \b2v_inst5.count_1_5\ : std_logic;
signal \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst5.m4_0\ : std_logic;
signal \b2v_inst5.N_2898_i_cascade_\ : std_logic;
signal \N_413\ : std_logic;
signal \b2v_inst5.curr_state_0_0\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst5.curr_state_RNIZ0Z_1\ : std_logic;
signal \b2v_inst5.N_2898_i\ : std_logic;
signal \b2v_inst5.count_0_sqmuxa\ : std_logic;
signal \b2v_inst11.N_172_i\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_2_i_o3_out\ : std_logic;
signal \b2v_inst11.N_19_cascade_\ : std_logic;
signal \rsmrstn_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3_fast\ : std_logic;
signal \b2v_inst11.N_168_cascade_\ : std_logic;
signal \curr_state_RNID8DP1_0_0\ : std_logic;
signal \RSMRSTn_0\ : std_logic;
signal \b2v_inst11.count_clk_RNIDQ4A1Z0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_\ : std_logic;
signal \b2v_inst11.N_186_i_cascade_\ : std_logic;
signal \b2v_inst11.N_115_f0_cascade_\ : std_logic;
signal \b2v_inst11.N_381\ : std_logic;
signal \b2v_inst11.g0_i_a7_1_2\ : std_logic;
signal \b2v_inst16.curr_state_RNIUCAD1Z0Z_0\ : std_logic;
signal \b2v_inst16.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst16.N_268\ : std_logic;
signal \b2v_inst11.N_395\ : std_logic;
signal \b2v_inst11.N_159\ : std_logic;
signal \b2v_inst11.N_159_cascade_\ : std_logic;
signal \b2v_inst11.N_425\ : std_logic;
signal \b2v_inst11.g2\ : std_logic;
signal \b2v_inst11.N_366\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.N_406_cascade_\ : std_logic;
signal \b2v_inst11.func_stateZ1Z_0\ : std_logic;
signal \b2v_inst11.func_state_enZ0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_cascade_\ : std_logic;
signal \b2v_inst11.N_428\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_0\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\ : std_logic;
signal \b2v_inst11.N_369\ : std_logic;
signal \b2v_inst11.func_state_1_m2_ns_1_1_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_1_m2_ns_1_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_1_m2_0\ : std_logic;
signal \b2v_inst11.N_327\ : std_logic;
signal \b2v_inst11.func_state_1_m2_ns_1_1_1\ : std_logic;
signal \b2v_inst11.N_382_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_2\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_0\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_a3_1\ : std_logic;
signal \b2v_inst11.N_406\ : std_logic;
signal \b2v_inst11.func_state_1_m2_ns_1_1\ : std_logic;
signal \b2v_inst11.func_state_1_m2_1_cascade_\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.N_337\ : std_logic;
signal \b2v_inst11.N_338_cascade_\ : std_logic;
signal \b2v_inst11.N_76\ : std_logic;
signal \b2v_inst11.func_state_enZ0\ : std_logic;
signal \b2v_inst11.func_state_1_m2_1\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_5\ : std_logic;
signal \b2v_inst11.func_state_1_m2s2_i_0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_1\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_0\ : std_logic;
signal \b2v_inst11.func_state_RNINIV94_0_0\ : std_logic;
signal \b2v_inst11.count_clk_0_0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_7\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_7\ : std_logic;
signal \b2v_inst11.count_clk_0_10\ : std_logic;
signal \b2v_inst11.count_clk_1_10\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_13\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_11\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_10\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o2_4\ : std_logic;
signal \b2v_inst11.count_clk_1_12\ : std_logic;
signal \b2v_inst11.count_clk_0_12\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_12\ : std_logic;
signal \b2v_inst11.count_clk_1_13\ : std_logic;
signal \b2v_inst11.count_clk_0_13\ : std_logic;
signal \b2v_inst11.count_clk_en\ : std_logic;
signal \bfn_11_1_0_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst6.count_0_15\ : std_logic;
signal \b2v_inst6.count_rst\ : std_logic;
signal \b2v_inst6.countZ0Z_15\ : std_logic;
signal \b2v_inst6.countZ0Z_15_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_7\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_7_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_7\ : std_logic;
signal \b2v_inst6.count_0_7\ : std_logic;
signal \b2v_inst6.count_rst_7_cascade_\ : std_logic;
signal \b2v_inst6.count_en_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_6\ : std_logic;
signal \b2v_inst6.countZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_0_0_cascade_\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0\ : std_logic;
signal v33dsw_ok : std_logic;
signal \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_9\ : std_logic;
signal \b2v_inst36.count_rst_5\ : std_logic;
signal \b2v_inst36.count_2_9\ : std_logic;
signal \b2v_inst36.curr_state_RNINSDSZ0Z_0\ : std_logic;
signal \b2v_inst36.count_0_sqmuxa\ : std_logic;
signal \b2v_inst6.count_0_10\ : std_logic;
signal \b2v_inst6.count_rst_4\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_10\ : std_logic;
signal v33a_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal v1p8a_ok : std_logic;
signal v5a_ok : std_logic;
signal \b2v_inst6.count_rst_5_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_9_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst6.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst6.count_0_8\ : std_logic;
signal \b2v_inst6.curr_state_1_0\ : std_logic;
signal \b2v_inst6.curr_state_7_0_cascade_\ : std_logic;
signal \b2v_inst6.N_42\ : std_logic;
signal \b2v_inst6.curr_state_1_1\ : std_logic;
signal \b2v_inst6.N_42_cascade_\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst6.N_3053_i_cascade_\ : std_logic;
signal \b2v_inst6.N_3034_i\ : std_logic;
signal \b2v_inst6.N_3034_i_cascade_\ : std_logic;
signal \b2v_inst6.curr_state_RNIUP4B1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\ : std_logic;
signal \N_222\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst6.N_3053_i\ : std_logic;
signal \b2v_inst6.N_192\ : std_logic;
signal \N_241\ : std_logic;
signal \b2v_inst6.N_276_0\ : std_logic;
signal \b2v_inst6.curr_state_RNIUP4B1Z0Z_0\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_ok_0\ : std_logic;
signal \b2v_inst11.N_9\ : std_logic;
signal \b2v_inst11.N_172_cascade_\ : std_logic;
signal \b2v_inst11.g0_i_a7_1_3\ : std_logic;
signal \b2v_inst11.g0_i_0_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3_rep1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8\ : std_logic;
signal \b2v_inst11.N_295_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3_out\ : std_logic;
signal \b2v_inst11.N_355\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_0_2\ : std_logic;
signal \b2v_inst11.N_168\ : std_logic;
signal \b2v_inst11.dutycycle_RNIAEUL3Z0Z_2\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_2\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_6\ : std_logic;
signal \b2v_inst11.N_365\ : std_logic;
signal \b2v_inst11.func_state_RNI_2Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.N_186_i\ : std_logic;
signal \b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2\ : std_logic;
signal \b2v_inst11.func_state_1_ss0_i_0_o3_0_cascade_\ : std_logic;
signal \b2v_inst11.N_430\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3\ : std_logic;
signal \b2v_inst11.N_161\ : std_logic;
signal \b2v_inst11.N_339\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_eena_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_0\ : std_logic;
signal \b2v_inst11.N_119_f0_1\ : std_logic;
signal \b2v_inst11.dutycycle\ : std_logic;
signal \b2v_inst11.dutycycle_eena_0\ : std_logic;
signal \G_146\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_1\ : std_logic;
signal \b2v_inst11.dutycycle_eena_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_1\ : std_logic;
signal \b2v_inst11.N_224_iZ0\ : std_logic;
signal \b2v_inst11.count_off_1_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_330_N\ : std_logic;
signal \b2v_inst11.func_state\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.N_382\ : std_logic;
signal \b2v_inst11.count_clk_RNI_0Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.N_315_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7\ : std_logic;
signal \b2v_inst11.N_125_cascade_\ : std_logic;
signal \b2v_inst11.N_382_N\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_1\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_3\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_4\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_7\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_8\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_9\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_10\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_11\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_12\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_13\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14\ : std_logic;
signal \b2v_inst11.count_off_1_14\ : std_logic;
signal \b2v_inst11.count_off_0_14\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DTZ0Z63\ : std_logic;
signal \b2v_inst11.count_off_0_15\ : std_logic;
signal \b2v_inst11.count_off_1_6\ : std_logic;
signal \b2v_inst11.count_off_0_6\ : std_logic;
signal \b2v_inst11.count_off_1_7\ : std_logic;
signal \b2v_inst11.count_off_0_7\ : std_logic;
signal \b2v_inst11.count_off_1_8\ : std_logic;
signal \b2v_inst11.count_off_0_8\ : std_logic;
signal \b2v_inst6.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_4\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_4_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_10\ : std_logic;
signal \b2v_inst6.count_0_4\ : std_logic;
signal \b2v_inst6.count_rst_11_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst6.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst6.count_0_3\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_2\ : std_logic;
signal \b2v_inst6.count_0_14\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_13_c_RNI06SPZ0Z1\ : std_logic;
signal \b2v_inst6.countZ0Z_14\ : std_logic;
signal \b2v_inst6.count_0_2\ : std_logic;
signal \b2v_inst6.countZ0Z_14_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_12\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_12\ : std_logic;
signal \b2v_inst6.count_rst_2\ : std_logic;
signal \b2v_inst6.count_0_12\ : std_logic;
signal \b2v_inst6.count_rst_1\ : std_logic;
signal \b2v_inst6.count_0_13\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_13\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\ : std_logic;
signal \b2v_inst6.count_0_6\ : std_logic;
signal \b2v_inst6.N_394_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_5\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst6.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst6.count_0_5\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst6.N_394\ : std_logic;
signal \b2v_inst6.count_rst_3_cascade_\ : std_logic;
signal \b2v_inst6.count_0_11\ : std_logic;
signal \b2v_inst6.count_RNIM6FE1Z0Z_0\ : std_logic;
signal \b2v_inst6.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_11\ : std_logic;
signal \b2v_inst6.count_rst_13_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_5_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_6_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_3_0_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_7_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_1_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_12_0_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_2_0\ : std_logic;
signal \b2v_inst6.N_389\ : std_logic;
signal \b2v_inst6.N_389_cascade_\ : std_logic;
signal \b2v_inst6.count_0_0\ : std_logic;
signal \b2v_inst6.count_rst_13\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_1\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_1_cascade_\ : std_logic;
signal \b2v_inst6.count_0_1\ : std_logic;
signal \b2v_inst6.curr_state_RNIM6FE1Z0Z_1\ : std_logic;
signal \b2v_inst6.count_rst_5\ : std_logic;
signal \b2v_inst6.count_0_9\ : std_logic;
signal \b2v_inst6.countZ0Z_8\ : std_logic;
signal \b2v_inst6.count_en\ : std_logic;
signal \b2v_inst6.count_1_i_a3_4_0\ : std_logic;
signal \b2v_inst5.N_51\ : std_logic;
signal \b2v_inst5.curr_state_0_1\ : std_logic;
signal \N_606_g\ : std_logic;
signal \b2v_inst6.countZ0Z_0\ : std_logic;
signal \b2v_inst6.N_3036_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal v5s_ok : std_logic;
signal v33s_ok : std_logic;
signal \SYNTHESIZED_WIRE_8\ : std_logic;
signal vccinaux_en : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_0_cascade_\ : std_logic;
signal slp_s4n : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m1_ns_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m1\ : std_logic;
signal \b2v_inst11.g0_i_2\ : std_logic;
signal \b2v_inst11.g0_0_0Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.g0_13_1_cascade_\ : std_logic;
signal \b2v_inst11.N_4690_0_0_cascade_\ : std_logic;
signal \b2v_inst11.N_19_0\ : std_logic;
signal \b2v_inst11.N_19_1\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m0\ : std_logic;
signal \b2v_inst11.g3_3\ : std_logic;
signal \b2v_inst11.N_172\ : std_logic;
signal \b2v_inst11.N_200_i\ : std_logic;
signal \b2v_inst11.N_3099_0_0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_2\ : std_logic;
signal \b2v_inst11.N_237\ : std_logic;
signal \b2v_inst11.N_293_0_0\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_6\ : std_logic;
signal \b2v_inst11.g2_1_0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_5\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_0\ : std_logic;
signal \G_6_i_a3_1\ : std_logic;
signal \N_5_cascade_\ : std_logic;
signal v5s_enn : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_rn_1\ : std_logic;
signal \b2v_inst11_un1_clk_100khz_52_and_i_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_sn\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_0_cascade_\ : std_logic;
signal \b2v_inst11.N_6063_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_eena_14_0_0\ : std_logic;
signal slp_s3n : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal rsmrstn : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0\ : std_logic;
signal \b2v_inst11.N_2946_i\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_5\ : std_logic;
signal \b2v_inst11.g0_1_1\ : std_logic;
signal vddq_ok : std_logic;
signal \VCCST_EN_i_0_o3_0\ : std_logic;
signal \b2v_inst16.N_208_0\ : std_logic;
signal \b2v_inst11.count_off_1_1\ : std_logic;
signal \b2v_inst11.count_offZ0Z_6\ : std_logic;
signal \b2v_inst11.count_offZ0Z_5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_offZ0Z_2\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_9_cascade_\ : std_logic;
signal \b2v_inst11.count_off_RNI_0Z0Z_1\ : std_logic;
signal \b2v_inst11.count_offZ0Z_15\ : std_logic;
signal \b2v_inst11.count_offZ0Z_13\ : std_logic;
signal \b2v_inst11.count_offZ0Z_14\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_10\ : std_logic;
signal \b2v_inst11.count_offZ0Z_7\ : std_logic;
signal \b2v_inst11.count_offZ0Z_8\ : std_logic;
signal \b2v_inst11.count_offZ0Z_3\ : std_logic;
signal \b2v_inst11.count_offZ0Z_4\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_8\ : std_logic;
signal \b2v_inst11.count_offZ0Z_1\ : std_logic;
signal \b2v_inst11.count_off_0_1\ : std_logic;
signal \b2v_inst11.count_offZ0Z_0\ : std_logic;
signal \b2v_inst11.N_125\ : std_logic;
signal \b2v_inst11.count_off_0_0\ : std_logic;
signal \b2v_inst11.count_off_0_9\ : std_logic;
signal \b2v_inst11.count_off_1_9\ : std_logic;
signal \b2v_inst11.count_offZ0Z_9\ : std_logic;
signal \b2v_inst11.count_offZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_11\ : std_logic;
signal \b2v_inst11.count_offZ0Z_10\ : std_logic;
signal \b2v_inst11.count_off_1_10\ : std_logic;
signal \b2v_inst11.count_off_0_10\ : std_logic;
signal \b2v_inst11.count_offZ0Z_11\ : std_logic;
signal \b2v_inst11.count_off_1_11\ : std_logic;
signal \b2v_inst11.count_off_0_11\ : std_logic;
signal \b2v_inst11.count_offZ0Z_12\ : std_logic;
signal \b2v_inst11.count_off_1_12\ : std_logic;
signal \b2v_inst11.count_off_0_12\ : std_logic;
signal \b2v_inst11.count_off_1_13\ : std_logic;
signal \b2v_inst11.count_off_0_13\ : std_logic;
signal \b2v_inst11.count_off_1_2\ : std_logic;
signal \b2v_inst11.count_off_0_2\ : std_logic;
signal \b2v_inst11.count_off_1_3\ : std_logic;
signal \b2v_inst11.count_off_0_3\ : std_logic;
signal \b2v_inst11.count_off_1_4\ : std_logic;
signal \b2v_inst11.count_off_0_4\ : std_logic;
signal \b2v_inst11.count_off_1_5\ : std_logic;
signal \b2v_inst11.count_off_0_5\ : std_logic;
signal fpga_osc : std_logic;
signal \b2v_inst11.dutycycle_RNIHJNV7Z0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    \SUSWARN_N_wire\ <= SUSWARN_N;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    \VCCINAUX_VR_PE_wire\ <= VCCINAUX_VR_PE;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    \VCCIN_VR_PE_wire\ <= VCCIN_VR_PE;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37287\,
            DIN => \N__37286\,
            DOUT => \N__37285\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37287\,
            PADOUT => \N__37286\,
            PADIN => \N__37285\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccinaux,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37278\,
            DIN => \N__37277\,
            DOUT => \N__37276\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37278\,
            PADOUT => \N__37277\,
            PADIN => \N__37276\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37269\,
            DIN => \N__37268\,
            DOUT => \N__37267\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37269\,
            PADOUT => \N__37268\,
            PADIN => \N__37267\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37260\,
            DIN => \N__37259\,
            DOUT => \N__37258\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37260\,
            PADOUT => \N__37259\,
            PADIN => \N__37258\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18191\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37251\,
            DIN => \N__37250\,
            DOUT => \N__37249\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37251\,
            PADOUT => \N__37250\,
            PADIN => \N__37249\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37242\,
            DIN => \N__37241\,
            DOUT => \N__37240\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37242\,
            PADOUT => \N__37241\,
            PADIN => \N__37240\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37233\,
            DIN => \N__37232\,
            DOUT => \N__37231\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37233\,
            PADOUT => \N__37232\,
            PADIN => \N__37231\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37224\,
            DIN => \N__37223\,
            DOUT => \N__37222\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37224\,
            PADOUT => \N__37223\,
            PADIN => \N__37222\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37215\,
            DIN => \N__37214\,
            DOUT => \N__37213\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37215\,
            PADOUT => \N__37214\,
            PADIN => \N__37213\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34945\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37206\,
            DIN => \N__37205\,
            DOUT => \N__37204\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37206\,
            PADOUT => \N__37205\,
            PADIN => \N__37204\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37197\,
            DIN => \N__37196\,
            DOUT => \N__37195\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37197\,
            PADOUT => \N__37196\,
            PADIN => \N__37195\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37188\,
            DIN => \N__37187\,
            DOUT => \N__37186\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37188\,
            PADOUT => \N__37187\,
            PADIN => \N__37186\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17168\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37179\,
            DIN => \N__37178\,
            DOUT => \N__37177\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37179\,
            PADOUT => \N__37178\,
            PADIN => \N__37177\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37170\,
            DIN => \N__37169\,
            DOUT => \N__37168\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37170\,
            PADOUT => \N__37169\,
            PADIN => \N__37168\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37161\,
            DIN => \N__37160\,
            DOUT => \N__37159\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37161\,
            PADOUT => \N__37160\,
            PADIN => \N__37159\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37152\,
            DIN => \N__37151\,
            DOUT => \N__37150\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37152\,
            PADOUT => \N__37151\,
            PADIN => \N__37150\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37143\,
            DIN => \N__37142\,
            DOUT => \N__37141\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37143\,
            PADOUT => \N__37142\,
            PADIN => \N__37141\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19916\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37134\,
            DIN => \N__37133\,
            DOUT => \N__37132\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37134\,
            PADOUT => \N__37133\,
            PADIN => \N__37132\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33dsw_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37125\,
            DIN => \N__37124\,
            DOUT => \N__37123\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37125\,
            PADOUT => \N__37124\,
            PADIN => \N__37123\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37116\,
            DIN => \N__37115\,
            DOUT => \N__37114\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37116\,
            PADOUT => \N__37115\,
            PADIN => \N__37114\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37107\,
            DIN => \N__37106\,
            DOUT => \N__37105\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37107\,
            PADOUT => \N__37106\,
            PADIN => \N__37105\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37098\,
            DIN => \N__37097\,
            DOUT => \N__37096\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37098\,
            PADOUT => \N__37097\,
            PADIN => \N__37096\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37089\,
            DIN => \N__37088\,
            DOUT => \N__37087\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37089\,
            PADOUT => \N__37088\,
            PADIN => \N__37087\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37080\,
            DIN => \N__37079\,
            DOUT => \N__37078\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37080\,
            PADOUT => \N__37079\,
            PADIN => \N__37078\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37071\,
            DIN => \N__37070\,
            DOUT => \N__37069\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37071\,
            PADOUT => \N__37070\,
            PADIN => \N__37069\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34319\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37062\,
            DIN => \N__37061\,
            DOUT => \N__37060\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37062\,
            PADOUT => \N__37061\,
            PADIN => \N__37060\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37053\,
            DIN => \N__37052\,
            DOUT => \N__37051\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37053\,
            PADOUT => \N__37052\,
            PADIN => \N__37051\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17344\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37044\,
            DIN => \N__37043\,
            DOUT => \N__37042\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37044\,
            PADOUT => \N__37043\,
            PADIN => \N__37042\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17354\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37035\,
            DIN => \N__37034\,
            DOUT => \N__37033\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37035\,
            PADOUT => \N__37034\,
            PADIN => \N__37033\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37026\,
            DIN => \N__37025\,
            DOUT => \N__37024\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37026\,
            PADOUT => \N__37025\,
            PADIN => \N__37024\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37017\,
            DIN => \N__37016\,
            DOUT => \N__37015\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37017\,
            PADOUT => \N__37016\,
            PADIN => \N__37015\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37008\,
            DIN => \N__37007\,
            DOUT => \N__37006\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37008\,
            PADOUT => \N__37007\,
            PADIN => \N__37006\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36999\,
            DIN => \N__36998\,
            DOUT => \N__36997\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36999\,
            PADOUT => \N__36998\,
            PADIN => \N__36997\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36990\,
            DIN => \N__36989\,
            DOUT => \N__36988\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36990\,
            PADOUT => \N__36989\,
            PADIN => \N__36988\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19379\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36981\,
            DIN => \N__36980\,
            DOUT => \N__36979\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36981\,
            PADOUT => \N__36980\,
            PADIN => \N__36979\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36972\,
            DIN => \N__36971\,
            DOUT => \N__36970\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36972\,
            PADOUT => \N__36971\,
            PADIN => \N__36970\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17771\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36963\,
            DIN => \N__36962\,
            DOUT => \N__36961\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36963\,
            PADOUT => \N__36962\,
            PADIN => \N__36961\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36954\,
            DIN => \N__36953\,
            DOUT => \N__36952\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36954\,
            PADOUT => \N__36953\,
            PADIN => \N__36952\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36945\,
            DIN => \N__36944\,
            DOUT => \N__36943\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36945\,
            PADOUT => \N__36944\,
            PADIN => \N__36943\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36936\,
            DIN => \N__36935\,
            DOUT => \N__36934\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36936\,
            PADOUT => \N__36935\,
            PADIN => \N__36934\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36927\,
            DIN => \N__36926\,
            DOUT => \N__36925\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36927\,
            PADOUT => \N__36926\,
            PADIN => \N__36925\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32938\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36918\,
            DIN => \N__36917\,
            DOUT => \N__36916\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36918\,
            PADOUT => \N__36917\,
            PADIN => \N__36916\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36909\,
            DIN => \N__36908\,
            DOUT => \N__36907\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36909\,
            PADOUT => \N__36908\,
            PADIN => \N__36907\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34946\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36900\,
            DIN => \N__36899\,
            DOUT => \N__36898\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36900\,
            PADOUT => \N__36899\,
            PADIN => \N__36898\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36891\,
            DIN => \N__36890\,
            DOUT => \N__36889\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36891\,
            PADOUT => \N__36890\,
            PADIN => \N__36889\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24212\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36882\,
            DIN => \N__36881\,
            DOUT => \N__36880\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36882\,
            PADOUT => \N__36881\,
            PADIN => \N__36880\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32060\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36873\,
            DIN => \N__36872\,
            DOUT => \N__36871\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36873\,
            PADOUT => \N__36872\,
            PADIN => \N__36871\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36864\,
            DIN => \N__36863\,
            DOUT => \N__36862\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36864\,
            PADOUT => \N__36863\,
            PADIN => \N__36862\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36855\,
            DIN => \N__36854\,
            DOUT => \N__36853\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36855\,
            PADOUT => \N__36854\,
            PADIN => \N__36853\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36846\,
            DIN => \N__36845\,
            DOUT => \N__36844\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36846\,
            PADOUT => \N__36845\,
            PADIN => \N__36844\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36837\,
            DIN => \N__36836\,
            DOUT => \N__36835\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36837\,
            PADOUT => \N__36836\,
            PADIN => \N__36835\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32951\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36828\,
            DIN => \N__36827\,
            DOUT => \N__36826\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36828\,
            PADOUT => \N__36827\,
            PADIN => \N__36826\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36819\,
            DIN => \N__36818\,
            DOUT => \N__36817\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36819\,
            PADOUT => \N__36818\,
            PADIN => \N__36817\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36810\,
            DIN => \N__36809\,
            DOUT => \N__36808\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36810\,
            PADOUT => \N__36809\,
            PADIN => \N__36808\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36801\,
            DIN => \N__36800\,
            DOUT => \N__36799\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36801\,
            PADOUT => \N__36800\,
            PADIN => \N__36799\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36792\,
            DIN => \N__36791\,
            DOUT => \N__36790\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36792\,
            PADOUT => \N__36791\,
            PADIN => \N__36790\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36783\,
            DIN => \N__36782\,
            DOUT => \N__36781\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36783\,
            PADOUT => \N__36782\,
            PADIN => \N__36781\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36774\,
            DIN => \N__36773\,
            DOUT => \N__36772\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36774\,
            PADOUT => \N__36773\,
            PADIN => \N__36772\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17337\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36765\,
            DIN => \N__36764\,
            DOUT => \N__36763\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36765\,
            PADOUT => \N__36764\,
            PADIN => \N__36763\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__8563\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__36743\,
            I => \N__36739\
        );

    \I__8561\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36736\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__36739\,
            I => \N__36733\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__36736\,
            I => \b2v_inst11.count_off_1_3\
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__36733\,
            I => \b2v_inst11.count_off_1_3\
        );

    \I__8557\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__36722\,
            I => \b2v_inst11.count_off_0_3\
        );

    \I__8554\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36716\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__36716\,
            I => \N__36712\
        );

    \I__8552\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36709\
        );

    \I__8551\ : Span4Mux_h
    port map (
            O => \N__36712\,
            I => \N__36706\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__36709\,
            I => \b2v_inst11.count_off_1_4\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__36706\,
            I => \b2v_inst11.count_off_1_4\
        );

    \I__8548\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36698\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36695\
        );

    \I__8546\ : Odrv4
    port map (
            O => \N__36695\,
            I => \b2v_inst11.count_off_0_4\
        );

    \I__8545\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36689\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36685\
        );

    \I__8543\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36682\
        );

    \I__8542\ : Span4Mux_s3_v
    port map (
            O => \N__36685\,
            I => \N__36679\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__36682\,
            I => \b2v_inst11.count_off_1_5\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__36679\,
            I => \b2v_inst11.count_off_1_5\
        );

    \I__8539\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36671\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36668\
        );

    \I__8537\ : Odrv4
    port map (
            O => \N__36668\,
            I => \b2v_inst11.count_off_0_5\
        );

    \I__8536\ : ClkMux
    port map (
            O => \N__36665\,
            I => \N__36662\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__36662\,
            I => \N__36658\
        );

    \I__8534\ : ClkMux
    port map (
            O => \N__36661\,
            I => \N__36653\
        );

    \I__8533\ : Span4Mux_s3_h
    port map (
            O => \N__36658\,
            I => \N__36649\
        );

    \I__8532\ : ClkMux
    port map (
            O => \N__36657\,
            I => \N__36646\
        );

    \I__8531\ : ClkMux
    port map (
            O => \N__36656\,
            I => \N__36643\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__36653\,
            I => \N__36640\
        );

    \I__8529\ : ClkMux
    port map (
            O => \N__36652\,
            I => \N__36637\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__36649\,
            I => \N__36628\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__36646\,
            I => \N__36628\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__36643\,
            I => \N__36628\
        );

    \I__8525\ : Span4Mux_v
    port map (
            O => \N__36640\,
            I => \N__36623\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__36637\,
            I => \N__36623\
        );

    \I__8523\ : ClkMux
    port map (
            O => \N__36636\,
            I => \N__36620\
        );

    \I__8522\ : ClkMux
    port map (
            O => \N__36635\,
            I => \N__36615\
        );

    \I__8521\ : Span4Mux_v
    port map (
            O => \N__36628\,
            I => \N__36608\
        );

    \I__8520\ : Span4Mux_h
    port map (
            O => \N__36623\,
            I => \N__36608\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__36620\,
            I => \N__36608\
        );

    \I__8518\ : ClkMux
    port map (
            O => \N__36619\,
            I => \N__36605\
        );

    \I__8517\ : ClkMux
    port map (
            O => \N__36618\,
            I => \N__36599\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__36615\,
            I => \N__36593\
        );

    \I__8515\ : Span4Mux_v
    port map (
            O => \N__36608\,
            I => \N__36593\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36590\
        );

    \I__8513\ : ClkMux
    port map (
            O => \N__36604\,
            I => \N__36587\
        );

    \I__8512\ : ClkMux
    port map (
            O => \N__36603\,
            I => \N__36583\
        );

    \I__8511\ : ClkMux
    port map (
            O => \N__36602\,
            I => \N__36576\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__36599\,
            I => \N__36572\
        );

    \I__8509\ : ClkMux
    port map (
            O => \N__36598\,
            I => \N__36569\
        );

    \I__8508\ : IoSpan4Mux
    port map (
            O => \N__36593\,
            I => \N__36565\
        );

    \I__8507\ : Span4Mux_v
    port map (
            O => \N__36590\,
            I => \N__36560\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__36587\,
            I => \N__36560\
        );

    \I__8505\ : ClkMux
    port map (
            O => \N__36586\,
            I => \N__36557\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__36583\,
            I => \N__36553\
        );

    \I__8503\ : ClkMux
    port map (
            O => \N__36582\,
            I => \N__36549\
        );

    \I__8502\ : ClkMux
    port map (
            O => \N__36581\,
            I => \N__36546\
        );

    \I__8501\ : ClkMux
    port map (
            O => \N__36580\,
            I => \N__36543\
        );

    \I__8500\ : ClkMux
    port map (
            O => \N__36579\,
            I => \N__36538\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__36576\,
            I => \N__36535\
        );

    \I__8498\ : ClkMux
    port map (
            O => \N__36575\,
            I => \N__36532\
        );

    \I__8497\ : Span4Mux_v
    port map (
            O => \N__36572\,
            I => \N__36527\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__36569\,
            I => \N__36524\
        );

    \I__8495\ : ClkMux
    port map (
            O => \N__36568\,
            I => \N__36521\
        );

    \I__8494\ : Span4Mux_s1_h
    port map (
            O => \N__36565\,
            I => \N__36514\
        );

    \I__8493\ : Span4Mux_h
    port map (
            O => \N__36560\,
            I => \N__36514\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__36557\,
            I => \N__36514\
        );

    \I__8491\ : ClkMux
    port map (
            O => \N__36556\,
            I => \N__36511\
        );

    \I__8490\ : IoSpan4Mux
    port map (
            O => \N__36553\,
            I => \N__36507\
        );

    \I__8489\ : ClkMux
    port map (
            O => \N__36552\,
            I => \N__36504\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__36549\,
            I => \N__36498\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__36546\,
            I => \N__36498\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__36543\,
            I => \N__36495\
        );

    \I__8485\ : ClkMux
    port map (
            O => \N__36542\,
            I => \N__36492\
        );

    \I__8484\ : ClkMux
    port map (
            O => \N__36541\,
            I => \N__36486\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__36538\,
            I => \N__36482\
        );

    \I__8482\ : Span4Mux_s2_v
    port map (
            O => \N__36535\,
            I => \N__36474\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36474\
        );

    \I__8480\ : ClkMux
    port map (
            O => \N__36531\,
            I => \N__36471\
        );

    \I__8479\ : ClkMux
    port map (
            O => \N__36530\,
            I => \N__36465\
        );

    \I__8478\ : Span4Mux_v
    port map (
            O => \N__36527\,
            I => \N__36454\
        );

    \I__8477\ : Span4Mux_s1_h
    port map (
            O => \N__36524\,
            I => \N__36454\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__36521\,
            I => \N__36454\
        );

    \I__8475\ : Span4Mux_h
    port map (
            O => \N__36514\,
            I => \N__36454\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__36511\,
            I => \N__36454\
        );

    \I__8473\ : ClkMux
    port map (
            O => \N__36510\,
            I => \N__36451\
        );

    \I__8472\ : Span4Mux_s2_h
    port map (
            O => \N__36507\,
            I => \N__36442\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__36504\,
            I => \N__36442\
        );

    \I__8470\ : ClkMux
    port map (
            O => \N__36503\,
            I => \N__36439\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__36498\,
            I => \N__36429\
        );

    \I__8468\ : Span4Mux_v
    port map (
            O => \N__36495\,
            I => \N__36429\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__36492\,
            I => \N__36429\
        );

    \I__8466\ : ClkMux
    port map (
            O => \N__36491\,
            I => \N__36426\
        );

    \I__8465\ : ClkMux
    port map (
            O => \N__36490\,
            I => \N__36423\
        );

    \I__8464\ : ClkMux
    port map (
            O => \N__36489\,
            I => \N__36417\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36413\
        );

    \I__8462\ : ClkMux
    port map (
            O => \N__36485\,
            I => \N__36410\
        );

    \I__8461\ : Span4Mux_s1_h
    port map (
            O => \N__36482\,
            I => \N__36407\
        );

    \I__8460\ : ClkMux
    port map (
            O => \N__36481\,
            I => \N__36404\
        );

    \I__8459\ : ClkMux
    port map (
            O => \N__36480\,
            I => \N__36398\
        );

    \I__8458\ : ClkMux
    port map (
            O => \N__36479\,
            I => \N__36395\
        );

    \I__8457\ : Span4Mux_v
    port map (
            O => \N__36474\,
            I => \N__36389\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__36471\,
            I => \N__36389\
        );

    \I__8455\ : ClkMux
    port map (
            O => \N__36470\,
            I => \N__36386\
        );

    \I__8454\ : ClkMux
    port map (
            O => \N__36469\,
            I => \N__36383\
        );

    \I__8453\ : ClkMux
    port map (
            O => \N__36468\,
            I => \N__36380\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__36465\,
            I => \N__36377\
        );

    \I__8451\ : Span4Mux_v
    port map (
            O => \N__36454\,
            I => \N__36372\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36372\
        );

    \I__8449\ : ClkMux
    port map (
            O => \N__36450\,
            I => \N__36369\
        );

    \I__8448\ : ClkMux
    port map (
            O => \N__36449\,
            I => \N__36364\
        );

    \I__8447\ : ClkMux
    port map (
            O => \N__36448\,
            I => \N__36361\
        );

    \I__8446\ : ClkMux
    port map (
            O => \N__36447\,
            I => \N__36357\
        );

    \I__8445\ : Span4Mux_s3_v
    port map (
            O => \N__36442\,
            I => \N__36351\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__36439\,
            I => \N__36351\
        );

    \I__8443\ : ClkMux
    port map (
            O => \N__36438\,
            I => \N__36346\
        );

    \I__8442\ : ClkMux
    port map (
            O => \N__36437\,
            I => \N__36343\
        );

    \I__8441\ : ClkMux
    port map (
            O => \N__36436\,
            I => \N__36340\
        );

    \I__8440\ : Span4Mux_v
    port map (
            O => \N__36429\,
            I => \N__36332\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__36426\,
            I => \N__36332\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__36423\,
            I => \N__36332\
        );

    \I__8437\ : ClkMux
    port map (
            O => \N__36422\,
            I => \N__36329\
        );

    \I__8436\ : ClkMux
    port map (
            O => \N__36421\,
            I => \N__36326\
        );

    \I__8435\ : ClkMux
    port map (
            O => \N__36420\,
            I => \N__36323\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__36417\,
            I => \N__36319\
        );

    \I__8433\ : ClkMux
    port map (
            O => \N__36416\,
            I => \N__36316\
        );

    \I__8432\ : Span4Mux_h
    port map (
            O => \N__36413\,
            I => \N__36309\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__36410\,
            I => \N__36309\
        );

    \I__8430\ : Span4Mux_h
    port map (
            O => \N__36407\,
            I => \N__36304\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__36404\,
            I => \N__36304\
        );

    \I__8428\ : ClkMux
    port map (
            O => \N__36403\,
            I => \N__36301\
        );

    \I__8427\ : ClkMux
    port map (
            O => \N__36402\,
            I => \N__36298\
        );

    \I__8426\ : ClkMux
    port map (
            O => \N__36401\,
            I => \N__36295\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__36398\,
            I => \N__36292\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__36395\,
            I => \N__36288\
        );

    \I__8423\ : ClkMux
    port map (
            O => \N__36394\,
            I => \N__36285\
        );

    \I__8422\ : Span4Mux_v
    port map (
            O => \N__36389\,
            I => \N__36280\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__36386\,
            I => \N__36280\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__36383\,
            I => \N__36277\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__36380\,
            I => \N__36274\
        );

    \I__8418\ : Span4Mux_s1_h
    port map (
            O => \N__36377\,
            I => \N__36267\
        );

    \I__8417\ : Span4Mux_s1_v
    port map (
            O => \N__36372\,
            I => \N__36267\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__36369\,
            I => \N__36267\
        );

    \I__8415\ : ClkMux
    port map (
            O => \N__36368\,
            I => \N__36264\
        );

    \I__8414\ : ClkMux
    port map (
            O => \N__36367\,
            I => \N__36260\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__36364\,
            I => \N__36257\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__36361\,
            I => \N__36254\
        );

    \I__8411\ : ClkMux
    port map (
            O => \N__36360\,
            I => \N__36251\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__36357\,
            I => \N__36248\
        );

    \I__8409\ : ClkMux
    port map (
            O => \N__36356\,
            I => \N__36245\
        );

    \I__8408\ : Span4Mux_v
    port map (
            O => \N__36351\,
            I => \N__36241\
        );

    \I__8407\ : ClkMux
    port map (
            O => \N__36350\,
            I => \N__36238\
        );

    \I__8406\ : ClkMux
    port map (
            O => \N__36349\,
            I => \N__36235\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__36346\,
            I => \N__36231\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__36343\,
            I => \N__36228\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__36340\,
            I => \N__36225\
        );

    \I__8402\ : ClkMux
    port map (
            O => \N__36339\,
            I => \N__36222\
        );

    \I__8401\ : Span4Mux_v
    port map (
            O => \N__36332\,
            I => \N__36213\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__36329\,
            I => \N__36213\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__36326\,
            I => \N__36213\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__36323\,
            I => \N__36213\
        );

    \I__8397\ : ClkMux
    port map (
            O => \N__36322\,
            I => \N__36210\
        );

    \I__8396\ : Span4Mux_s3_v
    port map (
            O => \N__36319\,
            I => \N__36202\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__36316\,
            I => \N__36202\
        );

    \I__8394\ : ClkMux
    port map (
            O => \N__36315\,
            I => \N__36199\
        );

    \I__8393\ : ClkMux
    port map (
            O => \N__36314\,
            I => \N__36195\
        );

    \I__8392\ : Span4Mux_v
    port map (
            O => \N__36309\,
            I => \N__36185\
        );

    \I__8391\ : Span4Mux_v
    port map (
            O => \N__36304\,
            I => \N__36185\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__36301\,
            I => \N__36185\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__36298\,
            I => \N__36182\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__36295\,
            I => \N__36179\
        );

    \I__8387\ : Span4Mux_s1_h
    port map (
            O => \N__36292\,
            I => \N__36176\
        );

    \I__8386\ : ClkMux
    port map (
            O => \N__36291\,
            I => \N__36173\
        );

    \I__8385\ : Span4Mux_v
    port map (
            O => \N__36288\,
            I => \N__36168\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__36285\,
            I => \N__36168\
        );

    \I__8383\ : Span4Mux_v
    port map (
            O => \N__36280\,
            I => \N__36156\
        );

    \I__8382\ : Span4Mux_s2_h
    port map (
            O => \N__36277\,
            I => \N__36156\
        );

    \I__8381\ : Span4Mux_s2_h
    port map (
            O => \N__36274\,
            I => \N__36156\
        );

    \I__8380\ : Span4Mux_h
    port map (
            O => \N__36267\,
            I => \N__36156\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__36264\,
            I => \N__36156\
        );

    \I__8378\ : ClkMux
    port map (
            O => \N__36263\,
            I => \N__36153\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__36260\,
            I => \N__36150\
        );

    \I__8376\ : Span4Mux_s2_h
    port map (
            O => \N__36257\,
            I => \N__36139\
        );

    \I__8375\ : Span4Mux_h
    port map (
            O => \N__36254\,
            I => \N__36139\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__36251\,
            I => \N__36139\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__36248\,
            I => \N__36139\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__36245\,
            I => \N__36139\
        );

    \I__8371\ : ClkMux
    port map (
            O => \N__36244\,
            I => \N__36136\
        );

    \I__8370\ : Span4Mux_v
    port map (
            O => \N__36241\,
            I => \N__36131\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__36238\,
            I => \N__36131\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__36235\,
            I => \N__36128\
        );

    \I__8367\ : ClkMux
    port map (
            O => \N__36234\,
            I => \N__36125\
        );

    \I__8366\ : Span4Mux_h
    port map (
            O => \N__36231\,
            I => \N__36116\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__36228\,
            I => \N__36116\
        );

    \I__8364\ : Span4Mux_h
    port map (
            O => \N__36225\,
            I => \N__36116\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__36222\,
            I => \N__36116\
        );

    \I__8362\ : IoSpan4Mux
    port map (
            O => \N__36213\,
            I => \N__36113\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__36210\,
            I => \N__36110\
        );

    \I__8360\ : ClkMux
    port map (
            O => \N__36209\,
            I => \N__36107\
        );

    \I__8359\ : ClkMux
    port map (
            O => \N__36208\,
            I => \N__36104\
        );

    \I__8358\ : ClkMux
    port map (
            O => \N__36207\,
            I => \N__36100\
        );

    \I__8357\ : Span4Mux_v
    port map (
            O => \N__36202\,
            I => \N__36096\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__36199\,
            I => \N__36093\
        );

    \I__8355\ : ClkMux
    port map (
            O => \N__36198\,
            I => \N__36090\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__36195\,
            I => \N__36087\
        );

    \I__8353\ : ClkMux
    port map (
            O => \N__36194\,
            I => \N__36084\
        );

    \I__8352\ : ClkMux
    port map (
            O => \N__36193\,
            I => \N__36081\
        );

    \I__8351\ : ClkMux
    port map (
            O => \N__36192\,
            I => \N__36078\
        );

    \I__8350\ : Span4Mux_v
    port map (
            O => \N__36185\,
            I => \N__36075\
        );

    \I__8349\ : Span4Mux_s1_h
    port map (
            O => \N__36182\,
            I => \N__36072\
        );

    \I__8348\ : Span4Mux_s2_h
    port map (
            O => \N__36179\,
            I => \N__36065\
        );

    \I__8347\ : Span4Mux_h
    port map (
            O => \N__36176\,
            I => \N__36065\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__36173\,
            I => \N__36065\
        );

    \I__8345\ : Span4Mux_v
    port map (
            O => \N__36168\,
            I => \N__36062\
        );

    \I__8344\ : ClkMux
    port map (
            O => \N__36167\,
            I => \N__36059\
        );

    \I__8343\ : Span4Mux_h
    port map (
            O => \N__36156\,
            I => \N__36054\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__36153\,
            I => \N__36054\
        );

    \I__8341\ : Span4Mux_s2_h
    port map (
            O => \N__36150\,
            I => \N__36047\
        );

    \I__8340\ : Span4Mux_v
    port map (
            O => \N__36139\,
            I => \N__36047\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__36136\,
            I => \N__36047\
        );

    \I__8338\ : Span4Mux_v
    port map (
            O => \N__36131\,
            I => \N__36040\
        );

    \I__8337\ : Span4Mux_s2_h
    port map (
            O => \N__36128\,
            I => \N__36040\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__36125\,
            I => \N__36040\
        );

    \I__8335\ : Span4Mux_v
    port map (
            O => \N__36116\,
            I => \N__36031\
        );

    \I__8334\ : IoSpan4Mux
    port map (
            O => \N__36113\,
            I => \N__36031\
        );

    \I__8333\ : Span4Mux_v
    port map (
            O => \N__36110\,
            I => \N__36031\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__36107\,
            I => \N__36031\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__36104\,
            I => \N__36028\
        );

    \I__8330\ : ClkMux
    port map (
            O => \N__36103\,
            I => \N__36025\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__36100\,
            I => \N__36021\
        );

    \I__8328\ : ClkMux
    port map (
            O => \N__36099\,
            I => \N__36018\
        );

    \I__8327\ : Span4Mux_h
    port map (
            O => \N__36096\,
            I => \N__36011\
        );

    \I__8326\ : Span4Mux_v
    port map (
            O => \N__36093\,
            I => \N__36011\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__36090\,
            I => \N__36011\
        );

    \I__8324\ : Span4Mux_h
    port map (
            O => \N__36087\,
            I => \N__36002\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__36084\,
            I => \N__36002\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__36081\,
            I => \N__36002\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__36078\,
            I => \N__36002\
        );

    \I__8320\ : Span4Mux_v
    port map (
            O => \N__36075\,
            I => \N__35994\
        );

    \I__8319\ : Span4Mux_h
    port map (
            O => \N__36072\,
            I => \N__35994\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__36065\,
            I => \N__35994\
        );

    \I__8317\ : Span4Mux_v
    port map (
            O => \N__36062\,
            I => \N__35989\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__36059\,
            I => \N__35989\
        );

    \I__8315\ : Span4Mux_h
    port map (
            O => \N__36054\,
            I => \N__35986\
        );

    \I__8314\ : IoSpan4Mux
    port map (
            O => \N__36047\,
            I => \N__35979\
        );

    \I__8313\ : IoSpan4Mux
    port map (
            O => \N__36040\,
            I => \N__35979\
        );

    \I__8312\ : IoSpan4Mux
    port map (
            O => \N__36031\,
            I => \N__35979\
        );

    \I__8311\ : Span4Mux_h
    port map (
            O => \N__36028\,
            I => \N__35974\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__36025\,
            I => \N__35974\
        );

    \I__8309\ : ClkMux
    port map (
            O => \N__36024\,
            I => \N__35971\
        );

    \I__8308\ : Span12Mux_s5_h
    port map (
            O => \N__36021\,
            I => \N__35962\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__36018\,
            I => \N__35962\
        );

    \I__8306\ : Sp12to4
    port map (
            O => \N__36011\,
            I => \N__35962\
        );

    \I__8305\ : Sp12to4
    port map (
            O => \N__36002\,
            I => \N__35962\
        );

    \I__8304\ : ClkMux
    port map (
            O => \N__36001\,
            I => \N__35959\
        );

    \I__8303\ : Odrv4
    port map (
            O => \N__35994\,
            I => fpga_osc
        );

    \I__8302\ : Odrv4
    port map (
            O => \N__35989\,
            I => fpga_osc
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__35986\,
            I => fpga_osc
        );

    \I__8300\ : Odrv4
    port map (
            O => \N__35979\,
            I => fpga_osc
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__35974\,
            I => fpga_osc
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__35971\,
            I => fpga_osc
        );

    \I__8297\ : Odrv12
    port map (
            O => \N__35962\,
            I => fpga_osc
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__35959\,
            I => fpga_osc
        );

    \I__8295\ : CEMux
    port map (
            O => \N__35942\,
            I => \N__35931\
        );

    \I__8294\ : CEMux
    port map (
            O => \N__35941\,
            I => \N__35926\
        );

    \I__8293\ : CEMux
    port map (
            O => \N__35940\,
            I => \N__35923\
        );

    \I__8292\ : CEMux
    port map (
            O => \N__35939\,
            I => \N__35920\
        );

    \I__8291\ : CEMux
    port map (
            O => \N__35938\,
            I => \N__35917\
        );

    \I__8290\ : InMux
    port map (
            O => \N__35937\,
            I => \N__35908\
        );

    \I__8289\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35908\
        );

    \I__8288\ : InMux
    port map (
            O => \N__35935\,
            I => \N__35908\
        );

    \I__8287\ : InMux
    port map (
            O => \N__35934\,
            I => \N__35908\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__35931\,
            I => \N__35905\
        );

    \I__8285\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35902\
        );

    \I__8284\ : InMux
    port map (
            O => \N__35929\,
            I => \N__35899\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__35926\,
            I => \N__35892\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__35923\,
            I => \N__35883\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__35920\,
            I => \N__35880\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__35917\,
            I => \N__35875\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__35908\,
            I => \N__35875\
        );

    \I__8278\ : Span4Mux_s3_v
    port map (
            O => \N__35905\,
            I => \N__35868\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__35902\,
            I => \N__35868\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__35899\,
            I => \N__35868\
        );

    \I__8275\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35859\
        );

    \I__8274\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35859\
        );

    \I__8273\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35859\
        );

    \I__8272\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35859\
        );

    \I__8271\ : Span4Mux_s2_h
    port map (
            O => \N__35892\,
            I => \N__35856\
        );

    \I__8270\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35843\
        );

    \I__8269\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35843\
        );

    \I__8268\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35843\
        );

    \I__8267\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35843\
        );

    \I__8266\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35843\
        );

    \I__8265\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35843\
        );

    \I__8264\ : Span4Mux_s0_h
    port map (
            O => \N__35883\,
            I => \N__35834\
        );

    \I__8263\ : Span4Mux_v
    port map (
            O => \N__35880\,
            I => \N__35834\
        );

    \I__8262\ : Span4Mux_s3_v
    port map (
            O => \N__35875\,
            I => \N__35834\
        );

    \I__8261\ : Span4Mux_v
    port map (
            O => \N__35868\,
            I => \N__35834\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__35859\,
            I => \N__35831\
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__35856\,
            I => \b2v_inst11.dutycycle_RNIHJNV7Z0Z_0\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__35843\,
            I => \b2v_inst11.dutycycle_RNIHJNV7Z0Z_0\
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__35834\,
            I => \b2v_inst11.dutycycle_RNIHJNV7Z0Z_0\
        );

    \I__8256\ : Odrv4
    port map (
            O => \N__35831\,
            I => \b2v_inst11.dutycycle_RNIHJNV7Z0Z_0\
        );

    \I__8255\ : CascadeMux
    port map (
            O => \N__35822\,
            I => \b2v_inst11.count_offZ0Z_9_cascade_\
        );

    \I__8254\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35816\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__35816\,
            I => \b2v_inst11.un34_clk_100khz_11\
        );

    \I__8252\ : CascadeMux
    port map (
            O => \N__35813\,
            I => \N__35809\
        );

    \I__8251\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35806\
        );

    \I__8250\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35803\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__35806\,
            I => \b2v_inst11.count_offZ0Z_10\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__35803\,
            I => \b2v_inst11.count_offZ0Z_10\
        );

    \I__8247\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35792\
        );

    \I__8246\ : InMux
    port map (
            O => \N__35797\,
            I => \N__35792\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__35792\,
            I => \b2v_inst11.count_off_1_10\
        );

    \I__8244\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35786\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__35786\,
            I => \b2v_inst11.count_off_0_10\
        );

    \I__8242\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35779\
        );

    \I__8241\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35776\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__35779\,
            I => \b2v_inst11.count_offZ0Z_11\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__35776\,
            I => \b2v_inst11.count_offZ0Z_11\
        );

    \I__8238\ : InMux
    port map (
            O => \N__35771\,
            I => \N__35765\
        );

    \I__8237\ : InMux
    port map (
            O => \N__35770\,
            I => \N__35765\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__35765\,
            I => \b2v_inst11.count_off_1_11\
        );

    \I__8235\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35759\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__35759\,
            I => \b2v_inst11.count_off_0_11\
        );

    \I__8233\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35752\
        );

    \I__8232\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35749\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__35752\,
            I => \b2v_inst11.count_offZ0Z_12\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__35749\,
            I => \b2v_inst11.count_offZ0Z_12\
        );

    \I__8229\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35740\
        );

    \I__8228\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35737\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__35740\,
            I => \b2v_inst11.count_off_1_12\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__35737\,
            I => \b2v_inst11.count_off_1_12\
        );

    \I__8225\ : InMux
    port map (
            O => \N__35732\,
            I => \N__35729\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__35729\,
            I => \b2v_inst11.count_off_0_12\
        );

    \I__8223\ : InMux
    port map (
            O => \N__35726\,
            I => \N__35722\
        );

    \I__8222\ : InMux
    port map (
            O => \N__35725\,
            I => \N__35719\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__35722\,
            I => \N__35716\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__35719\,
            I => \b2v_inst11.count_off_1_13\
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__35716\,
            I => \b2v_inst11.count_off_1_13\
        );

    \I__8218\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35708\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__35708\,
            I => \N__35705\
        );

    \I__8216\ : Span4Mux_h
    port map (
            O => \N__35705\,
            I => \N__35702\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__35702\,
            I => \b2v_inst11.count_off_0_13\
        );

    \I__8214\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35696\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__35696\,
            I => \N__35692\
        );

    \I__8212\ : InMux
    port map (
            O => \N__35695\,
            I => \N__35689\
        );

    \I__8211\ : Span4Mux_h
    port map (
            O => \N__35692\,
            I => \N__35686\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__35689\,
            I => \b2v_inst11.count_off_1_2\
        );

    \I__8209\ : Odrv4
    port map (
            O => \N__35686\,
            I => \b2v_inst11.count_off_1_2\
        );

    \I__8208\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35678\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__35675\,
            I => \b2v_inst11.count_off_0_2\
        );

    \I__8205\ : InMux
    port map (
            O => \N__35672\,
            I => \N__35668\
        );

    \I__8204\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35665\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__35668\,
            I => \N__35662\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35659\
        );

    \I__8201\ : Odrv4
    port map (
            O => \N__35662\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__35659\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__8199\ : InMux
    port map (
            O => \N__35654\,
            I => \N__35650\
        );

    \I__8198\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35647\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__35650\,
            I => \N__35644\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__35647\,
            I => \N__35641\
        );

    \I__8195\ : Span4Mux_v
    port map (
            O => \N__35644\,
            I => \N__35638\
        );

    \I__8194\ : Span4Mux_s2_h
    port map (
            O => \N__35641\,
            I => \N__35635\
        );

    \I__8193\ : Odrv4
    port map (
            O => \N__35638\,
            I => \b2v_inst11.count_offZ0Z_5\
        );

    \I__8192\ : Odrv4
    port map (
            O => \N__35635\,
            I => \b2v_inst11.count_offZ0Z_5\
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__35630\,
            I => \b2v_inst11.count_offZ0Z_1_cascade_\
        );

    \I__8190\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35623\
        );

    \I__8189\ : InMux
    port map (
            O => \N__35626\,
            I => \N__35620\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__35623\,
            I => \N__35617\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__35620\,
            I => \N__35614\
        );

    \I__8186\ : Span4Mux_v
    port map (
            O => \N__35617\,
            I => \N__35611\
        );

    \I__8185\ : Span4Mux_s2_h
    port map (
            O => \N__35614\,
            I => \N__35608\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__35611\,
            I => \b2v_inst11.count_offZ0Z_2\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__35608\,
            I => \b2v_inst11.count_offZ0Z_2\
        );

    \I__8182\ : CascadeMux
    port map (
            O => \N__35603\,
            I => \b2v_inst11.un34_clk_100khz_9_cascade_\
        );

    \I__8181\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35596\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__35599\,
            I => \N__35591\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__35596\,
            I => \N__35588\
        );

    \I__8178\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35578\
        );

    \I__8177\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35578\
        );

    \I__8176\ : InMux
    port map (
            O => \N__35591\,
            I => \N__35574\
        );

    \I__8175\ : Span4Mux_v
    port map (
            O => \N__35588\,
            I => \N__35571\
        );

    \I__8174\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35568\
        );

    \I__8173\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35561\
        );

    \I__8172\ : InMux
    port map (
            O => \N__35585\,
            I => \N__35561\
        );

    \I__8171\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35561\
        );

    \I__8170\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35558\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__35578\,
            I => \N__35555\
        );

    \I__8168\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35552\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__35574\,
            I => \N__35549\
        );

    \I__8166\ : Span4Mux_v
    port map (
            O => \N__35571\,
            I => \N__35542\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35542\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35542\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__35558\,
            I => \N__35537\
        );

    \I__8162\ : Span4Mux_h
    port map (
            O => \N__35555\,
            I => \N__35537\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__35552\,
            I => \b2v_inst11.count_off_RNI_0Z0Z_1\
        );

    \I__8160\ : Odrv12
    port map (
            O => \N__35549\,
            I => \b2v_inst11.count_off_RNI_0Z0Z_1\
        );

    \I__8159\ : Odrv4
    port map (
            O => \N__35542\,
            I => \b2v_inst11.count_off_RNI_0Z0Z_1\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__35537\,
            I => \b2v_inst11.count_off_RNI_0Z0Z_1\
        );

    \I__8157\ : InMux
    port map (
            O => \N__35528\,
            I => \N__35525\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__35525\,
            I => \N__35521\
        );

    \I__8155\ : InMux
    port map (
            O => \N__35524\,
            I => \N__35518\
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__35521\,
            I => \b2v_inst11.count_offZ0Z_15\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__35518\,
            I => \b2v_inst11.count_offZ0Z_15\
        );

    \I__8152\ : InMux
    port map (
            O => \N__35513\,
            I => \N__35510\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__35510\,
            I => \N__35507\
        );

    \I__8150\ : Span4Mux_s2_h
    port map (
            O => \N__35507\,
            I => \N__35503\
        );

    \I__8149\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35500\
        );

    \I__8148\ : Span4Mux_h
    port map (
            O => \N__35503\,
            I => \N__35497\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35494\
        );

    \I__8146\ : Odrv4
    port map (
            O => \N__35497\,
            I => \b2v_inst11.count_offZ0Z_13\
        );

    \I__8145\ : Odrv4
    port map (
            O => \N__35494\,
            I => \b2v_inst11.count_offZ0Z_13\
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__35489\,
            I => \N__35486\
        );

    \I__8143\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35483\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__35483\,
            I => \N__35479\
        );

    \I__8141\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35476\
        );

    \I__8140\ : Span4Mux_v
    port map (
            O => \N__35479\,
            I => \N__35471\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__35476\,
            I => \N__35471\
        );

    \I__8138\ : Odrv4
    port map (
            O => \N__35471\,
            I => \b2v_inst11.count_offZ0Z_14\
        );

    \I__8137\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__35465\,
            I => \b2v_inst11.un34_clk_100khz_10\
        );

    \I__8135\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35459\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__35459\,
            I => \N__35455\
        );

    \I__8133\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35452\
        );

    \I__8132\ : Span4Mux_v
    port map (
            O => \N__35455\,
            I => \N__35449\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__35452\,
            I => \N__35446\
        );

    \I__8130\ : Odrv4
    port map (
            O => \N__35449\,
            I => \b2v_inst11.count_offZ0Z_7\
        );

    \I__8129\ : Odrv4
    port map (
            O => \N__35446\,
            I => \b2v_inst11.count_offZ0Z_7\
        );

    \I__8128\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35438\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__35438\,
            I => \N__35434\
        );

    \I__8126\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35431\
        );

    \I__8125\ : Span4Mux_s1_h
    port map (
            O => \N__35434\,
            I => \N__35428\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__35431\,
            I => \N__35425\
        );

    \I__8123\ : Odrv4
    port map (
            O => \N__35428\,
            I => \b2v_inst11.count_offZ0Z_8\
        );

    \I__8122\ : Odrv12
    port map (
            O => \N__35425\,
            I => \b2v_inst11.count_offZ0Z_8\
        );

    \I__8121\ : CascadeMux
    port map (
            O => \N__35420\,
            I => \N__35417\
        );

    \I__8120\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35413\
        );

    \I__8119\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35410\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__35413\,
            I => \N__35407\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__35410\,
            I => \N__35404\
        );

    \I__8116\ : Span4Mux_v
    port map (
            O => \N__35407\,
            I => \N__35401\
        );

    \I__8115\ : Span4Mux_s2_h
    port map (
            O => \N__35404\,
            I => \N__35398\
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__35401\,
            I => \b2v_inst11.count_offZ0Z_3\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__35398\,
            I => \b2v_inst11.count_offZ0Z_3\
        );

    \I__8112\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35389\
        );

    \I__8111\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35386\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__35389\,
            I => \N__35383\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__35386\,
            I => \N__35380\
        );

    \I__8108\ : Span4Mux_s3_h
    port map (
            O => \N__35383\,
            I => \N__35377\
        );

    \I__8107\ : Span4Mux_s2_h
    port map (
            O => \N__35380\,
            I => \N__35374\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__35377\,
            I => \b2v_inst11.count_offZ0Z_4\
        );

    \I__8105\ : Odrv4
    port map (
            O => \N__35374\,
            I => \b2v_inst11.count_offZ0Z_4\
        );

    \I__8104\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__35366\,
            I => \b2v_inst11.un34_clk_100khz_8\
        );

    \I__8102\ : CascadeMux
    port map (
            O => \N__35363\,
            I => \N__35359\
        );

    \I__8101\ : InMux
    port map (
            O => \N__35362\,
            I => \N__35355\
        );

    \I__8100\ : InMux
    port map (
            O => \N__35359\,
            I => \N__35352\
        );

    \I__8099\ : InMux
    port map (
            O => \N__35358\,
            I => \N__35349\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__35355\,
            I => \N__35344\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__35352\,
            I => \N__35344\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__35349\,
            I => \b2v_inst11.count_offZ0Z_1\
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__35344\,
            I => \b2v_inst11.count_offZ0Z_1\
        );

    \I__8094\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__35336\,
            I => \b2v_inst11.count_off_0_1\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__35333\,
            I => \N__35329\
        );

    \I__8091\ : InMux
    port map (
            O => \N__35332\,
            I => \N__35318\
        );

    \I__8090\ : InMux
    port map (
            O => \N__35329\,
            I => \N__35318\
        );

    \I__8089\ : InMux
    port map (
            O => \N__35328\,
            I => \N__35318\
        );

    \I__8088\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35315\
        );

    \I__8087\ : InMux
    port map (
            O => \N__35326\,
            I => \N__35310\
        );

    \I__8086\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35310\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__35318\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__35315\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__35310\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__8082\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35288\
        );

    \I__8081\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35288\
        );

    \I__8080\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35288\
        );

    \I__8079\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35279\
        );

    \I__8078\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35279\
        );

    \I__8077\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35279\
        );

    \I__8076\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35279\
        );

    \I__8075\ : InMux
    port map (
            O => \N__35296\,
            I => \N__35266\
        );

    \I__8074\ : InMux
    port map (
            O => \N__35295\,
            I => \N__35266\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__35288\,
            I => \N__35261\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__35279\,
            I => \N__35261\
        );

    \I__8071\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35254\
        );

    \I__8070\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35254\
        );

    \I__8069\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35254\
        );

    \I__8068\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35245\
        );

    \I__8067\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35245\
        );

    \I__8066\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35245\
        );

    \I__8065\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35245\
        );

    \I__8064\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35242\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__35266\,
            I => \b2v_inst11.N_125\
        );

    \I__8062\ : Odrv4
    port map (
            O => \N__35261\,
            I => \b2v_inst11.N_125\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__35254\,
            I => \b2v_inst11.N_125\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__35245\,
            I => \b2v_inst11.N_125\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__35242\,
            I => \b2v_inst11.N_125\
        );

    \I__8058\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35228\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__35228\,
            I => \b2v_inst11.count_off_0_0\
        );

    \I__8056\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35222\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__35222\,
            I => \b2v_inst11.count_off_0_9\
        );

    \I__8054\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35213\
        );

    \I__8053\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35213\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__35213\,
            I => \b2v_inst11.count_off_1_9\
        );

    \I__8051\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35207\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__35207\,
            I => \b2v_inst11.count_offZ0Z_9\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__35204\,
            I => \N__35201\
        );

    \I__8048\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35193\
        );

    \I__8047\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35193\
        );

    \I__8046\ : InMux
    port map (
            O => \N__35199\,
            I => \N__35189\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__35198\,
            I => \N__35185\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__35193\,
            I => \N__35179\
        );

    \I__8043\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35176\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__35189\,
            I => \N__35172\
        );

    \I__8041\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35167\
        );

    \I__8040\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35167\
        );

    \I__8039\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35164\
        );

    \I__8038\ : InMux
    port map (
            O => \N__35183\,
            I => \N__35161\
        );

    \I__8037\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35158\
        );

    \I__8036\ : Span4Mux_v
    port map (
            O => \N__35179\,
            I => \N__35155\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__35176\,
            I => \N__35152\
        );

    \I__8034\ : InMux
    port map (
            O => \N__35175\,
            I => \N__35149\
        );

    \I__8033\ : Span4Mux_s1_h
    port map (
            O => \N__35172\,
            I => \N__35146\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__35167\,
            I => \N__35139\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__35164\,
            I => \N__35139\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__35161\,
            I => \N__35139\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__35158\,
            I => \N__35136\
        );

    \I__8028\ : Span4Mux_h
    port map (
            O => \N__35155\,
            I => \N__35128\
        );

    \I__8027\ : Span4Mux_h
    port map (
            O => \N__35152\,
            I => \N__35128\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__35149\,
            I => \N__35128\
        );

    \I__8025\ : Span4Mux_h
    port map (
            O => \N__35146\,
            I => \N__35121\
        );

    \I__8024\ : Span4Mux_v
    port map (
            O => \N__35139\,
            I => \N__35121\
        );

    \I__8023\ : Span4Mux_h
    port map (
            O => \N__35136\,
            I => \N__35121\
        );

    \I__8022\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35118\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__35128\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__35121\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__35118\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__8018\ : InMux
    port map (
            O => \N__35111\,
            I => \N__35097\
        );

    \I__8017\ : InMux
    port map (
            O => \N__35110\,
            I => \N__35097\
        );

    \I__8016\ : InMux
    port map (
            O => \N__35109\,
            I => \N__35097\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__35108\,
            I => \N__35085\
        );

    \I__8014\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35078\
        );

    \I__8013\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35078\
        );

    \I__8012\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35073\
        );

    \I__8011\ : InMux
    port map (
            O => \N__35104\,
            I => \N__35073\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__35097\,
            I => \N__35069\
        );

    \I__8009\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35066\
        );

    \I__8008\ : CascadeMux
    port map (
            O => \N__35095\,
            I => \N__35063\
        );

    \I__8007\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35059\
        );

    \I__8006\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35052\
        );

    \I__8005\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35052\
        );

    \I__8004\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35052\
        );

    \I__8003\ : InMux
    port map (
            O => \N__35090\,
            I => \N__35045\
        );

    \I__8002\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35045\
        );

    \I__8001\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35045\
        );

    \I__8000\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35040\
        );

    \I__7999\ : InMux
    port map (
            O => \N__35084\,
            I => \N__35040\
        );

    \I__7998\ : InMux
    port map (
            O => \N__35083\,
            I => \N__35037\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__35078\,
            I => \N__35032\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__35073\,
            I => \N__35032\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__35072\,
            I => \N__35027\
        );

    \I__7994\ : Span4Mux_s2_h
    port map (
            O => \N__35069\,
            I => \N__35022\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__35066\,
            I => \N__35019\
        );

    \I__7992\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35014\
        );

    \I__7991\ : InMux
    port map (
            O => \N__35062\,
            I => \N__35014\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__35059\,
            I => \N__35007\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__35052\,
            I => \N__35007\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__35045\,
            I => \N__35007\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__35040\,
            I => \N__35004\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__35037\,
            I => \N__34999\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__35032\,
            I => \N__34999\
        );

    \I__7984\ : InMux
    port map (
            O => \N__35031\,
            I => \N__34996\
        );

    \I__7983\ : InMux
    port map (
            O => \N__35030\,
            I => \N__34991\
        );

    \I__7982\ : InMux
    port map (
            O => \N__35027\,
            I => \N__34991\
        );

    \I__7981\ : InMux
    port map (
            O => \N__35026\,
            I => \N__34986\
        );

    \I__7980\ : InMux
    port map (
            O => \N__35025\,
            I => \N__34986\
        );

    \I__7979\ : Span4Mux_v
    port map (
            O => \N__35022\,
            I => \N__34983\
        );

    \I__7978\ : Span4Mux_v
    port map (
            O => \N__35019\,
            I => \N__34976\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__35014\,
            I => \N__34976\
        );

    \I__7976\ : Span4Mux_s3_h
    port map (
            O => \N__35007\,
            I => \N__34976\
        );

    \I__7975\ : Odrv12
    port map (
            O => \N__35004\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__34999\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__34996\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__34991\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__34986\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__34983\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__34976\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__7968\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34958\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__34958\,
            I => \N__34955\
        );

    \I__7966\ : Span4Mux_v
    port map (
            O => \N__34955\,
            I => \N__34952\
        );

    \I__7965\ : Odrv4
    port map (
            O => \N__34952\,
            I => \G_6_i_a3_1\
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__34949\,
            I => \N_5_cascade_\
        );

    \I__7963\ : IoInMux
    port map (
            O => \N__34946\,
            I => \N__34942\
        );

    \I__7962\ : IoInMux
    port map (
            O => \N__34945\,
            I => \N__34939\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__34942\,
            I => \N__34933\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__34939\,
            I => \N__34933\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__34938\,
            I => \N__34923\
        );

    \I__7958\ : IoSpan4Mux
    port map (
            O => \N__34933\,
            I => \N__34920\
        );

    \I__7957\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34916\
        );

    \I__7956\ : InMux
    port map (
            O => \N__34931\,
            I => \N__34913\
        );

    \I__7955\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34910\
        );

    \I__7954\ : InMux
    port map (
            O => \N__34929\,
            I => \N__34907\
        );

    \I__7953\ : InMux
    port map (
            O => \N__34928\,
            I => \N__34904\
        );

    \I__7952\ : InMux
    port map (
            O => \N__34927\,
            I => \N__34901\
        );

    \I__7951\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34898\
        );

    \I__7950\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34895\
        );

    \I__7949\ : Span4Mux_s3_h
    port map (
            O => \N__34920\,
            I => \N__34891\
        );

    \I__7948\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34888\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__34916\,
            I => \N__34885\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34878\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__34910\,
            I => \N__34878\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__34907\,
            I => \N__34875\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__34904\,
            I => \N__34870\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__34901\,
            I => \N__34870\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__34898\,
            I => \N__34865\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__34895\,
            I => \N__34865\
        );

    \I__7939\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34862\
        );

    \I__7938\ : Span4Mux_h
    port map (
            O => \N__34891\,
            I => \N__34857\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__34888\,
            I => \N__34857\
        );

    \I__7936\ : Span4Mux_v
    port map (
            O => \N__34885\,
            I => \N__34854\
        );

    \I__7935\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34849\
        );

    \I__7934\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34849\
        );

    \I__7933\ : Span12Mux_s3_h
    port map (
            O => \N__34878\,
            I => \N__34846\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__34875\,
            I => \N__34837\
        );

    \I__7931\ : Span4Mux_s3_h
    port map (
            O => \N__34870\,
            I => \N__34837\
        );

    \I__7930\ : Span4Mux_s3_h
    port map (
            O => \N__34865\,
            I => \N__34837\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__34862\,
            I => \N__34837\
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__34857\,
            I => v5s_enn
        );

    \I__7927\ : Odrv4
    port map (
            O => \N__34854\,
            I => v5s_enn
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__34849\,
            I => v5s_enn
        );

    \I__7925\ : Odrv12
    port map (
            O => \N__34846\,
            I => v5s_enn
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__34837\,
            I => v5s_enn
        );

    \I__7923\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34823\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__34823\,
            I => \N__34820\
        );

    \I__7921\ : Odrv12
    port map (
            O => \N__34820\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_rn_1\
        );

    \I__7920\ : CascadeMux
    port map (
            O => \N__34817\,
            I => \b2v_inst11_un1_clk_100khz_52_and_i_0_cascade_\
        );

    \I__7919\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34801\
        );

    \I__7918\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34792\
        );

    \I__7917\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34787\
        );

    \I__7916\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34787\
        );

    \I__7915\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34784\
        );

    \I__7914\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34779\
        );

    \I__7913\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34779\
        );

    \I__7912\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34776\
        );

    \I__7911\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34773\
        );

    \I__7910\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34770\
        );

    \I__7909\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34767\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__34801\,
            I => \N__34764\
        );

    \I__7907\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34757\
        );

    \I__7906\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34757\
        );

    \I__7905\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34757\
        );

    \I__7904\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34752\
        );

    \I__7903\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34752\
        );

    \I__7902\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34749\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__34792\,
            I => \N__34744\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__34787\,
            I => \N__34740\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__34784\,
            I => \N__34732\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__34779\,
            I => \N__34732\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__34776\,
            I => \N__34717\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__34773\,
            I => \N__34717\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__34770\,
            I => \N__34717\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__34767\,
            I => \N__34717\
        );

    \I__7893\ : Span4Mux_h
    port map (
            O => \N__34764\,
            I => \N__34717\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__34757\,
            I => \N__34717\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__34752\,
            I => \N__34717\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__34749\,
            I => \N__34714\
        );

    \I__7889\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34711\
        );

    \I__7888\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34708\
        );

    \I__7887\ : Span4Mux_s3_h
    port map (
            O => \N__34744\,
            I => \N__34705\
        );

    \I__7886\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34702\
        );

    \I__7885\ : Span4Mux_h
    port map (
            O => \N__34740\,
            I => \N__34699\
        );

    \I__7884\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34694\
        );

    \I__7883\ : InMux
    port map (
            O => \N__34738\,
            I => \N__34694\
        );

    \I__7882\ : InMux
    port map (
            O => \N__34737\,
            I => \N__34691\
        );

    \I__7881\ : Span4Mux_v
    port map (
            O => \N__34732\,
            I => \N__34686\
        );

    \I__7880\ : Span4Mux_v
    port map (
            O => \N__34717\,
            I => \N__34686\
        );

    \I__7879\ : Span4Mux_s2_h
    port map (
            O => \N__34714\,
            I => \N__34683\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__34711\,
            I => \N__34678\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__34708\,
            I => \N__34678\
        );

    \I__7876\ : Odrv4
    port map (
            O => \N__34705\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__34702\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7874\ : Odrv4
    port map (
            O => \N__34699\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__34694\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__34691\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7871\ : Odrv4
    port map (
            O => \N__34686\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__34683\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7869\ : Odrv12
    port map (
            O => \N__34678\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__7868\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34658\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__34658\,
            I => \N__34655\
        );

    \I__7866\ : Odrv12
    port map (
            O => \N__34655\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_sn\
        );

    \I__7865\ : CascadeMux
    port map (
            O => \N__34652\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_0_cascade_\
        );

    \I__7864\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__34646\,
            I => \b2v_inst11.N_6063_0_0\
        );

    \I__7862\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34637\
        );

    \I__7861\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34637\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__34637\,
            I => \N__34634\
        );

    \I__7859\ : Span4Mux_h
    port map (
            O => \N__34634\,
            I => \N__34631\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__34631\,
            I => \N__34628\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__34628\,
            I => \b2v_inst11.dutycycle_eena_14_0_0\
        );

    \I__7856\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34616\
        );

    \I__7855\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34611\
        );

    \I__7854\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34608\
        );

    \I__7853\ : CascadeMux
    port map (
            O => \N__34622\,
            I => \N__34605\
        );

    \I__7852\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34596\
        );

    \I__7851\ : InMux
    port map (
            O => \N__34620\,
            I => \N__34593\
        );

    \I__7850\ : InMux
    port map (
            O => \N__34619\,
            I => \N__34590\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__34616\,
            I => \N__34587\
        );

    \I__7848\ : InMux
    port map (
            O => \N__34615\,
            I => \N__34584\
        );

    \I__7847\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34581\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__34611\,
            I => \N__34578\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__34608\,
            I => \N__34575\
        );

    \I__7844\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34572\
        );

    \I__7843\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34569\
        );

    \I__7842\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34566\
        );

    \I__7841\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34563\
        );

    \I__7840\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34556\
        );

    \I__7839\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34556\
        );

    \I__7838\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34556\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__34596\,
            I => \N__34550\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__34593\,
            I => \N__34550\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__34590\,
            I => \N__34547\
        );

    \I__7834\ : Span4Mux_v
    port map (
            O => \N__34587\,
            I => \N__34544\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__34584\,
            I => \N__34539\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__34581\,
            I => \N__34539\
        );

    \I__7831\ : Span4Mux_v
    port map (
            O => \N__34578\,
            I => \N__34536\
        );

    \I__7830\ : Span4Mux_v
    port map (
            O => \N__34575\,
            I => \N__34531\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__34572\,
            I => \N__34531\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__34569\,
            I => \N__34526\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__34566\,
            I => \N__34526\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__34563\,
            I => \N__34521\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__34556\,
            I => \N__34521\
        );

    \I__7824\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34518\
        );

    \I__7823\ : Span4Mux_v
    port map (
            O => \N__34550\,
            I => \N__34515\
        );

    \I__7822\ : Span4Mux_v
    port map (
            O => \N__34547\,
            I => \N__34508\
        );

    \I__7821\ : Span4Mux_s2_h
    port map (
            O => \N__34544\,
            I => \N__34508\
        );

    \I__7820\ : Span4Mux_v
    port map (
            O => \N__34539\,
            I => \N__34508\
        );

    \I__7819\ : Span4Mux_s2_v
    port map (
            O => \N__34536\,
            I => \N__34503\
        );

    \I__7818\ : Span4Mux_v
    port map (
            O => \N__34531\,
            I => \N__34503\
        );

    \I__7817\ : Span4Mux_v
    port map (
            O => \N__34526\,
            I => \N__34496\
        );

    \I__7816\ : Span4Mux_h
    port map (
            O => \N__34521\,
            I => \N__34496\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__34518\,
            I => \N__34496\
        );

    \I__7814\ : Span4Mux_h
    port map (
            O => \N__34515\,
            I => \N__34488\
        );

    \I__7813\ : Span4Mux_v
    port map (
            O => \N__34508\,
            I => \N__34488\
        );

    \I__7812\ : Span4Mux_h
    port map (
            O => \N__34503\,
            I => \N__34483\
        );

    \I__7811\ : Span4Mux_v
    port map (
            O => \N__34496\,
            I => \N__34483\
        );

    \I__7810\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34480\
        );

    \I__7809\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34477\
        );

    \I__7808\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34474\
        );

    \I__7807\ : IoSpan4Mux
    port map (
            O => \N__34488\,
            I => \N__34469\
        );

    \I__7806\ : IoSpan4Mux
    port map (
            O => \N__34483\,
            I => \N__34469\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__34480\,
            I => \N__34462\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__34477\,
            I => \N__34462\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__34474\,
            I => \N__34462\
        );

    \I__7802\ : Odrv4
    port map (
            O => \N__34469\,
            I => slp_s3n
        );

    \I__7801\ : Odrv12
    port map (
            O => \N__34462\,
            I => slp_s3n
        );

    \I__7800\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34449\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__34456\,
            I => \N__34446\
        );

    \I__7798\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34442\
        );

    \I__7797\ : CascadeMux
    port map (
            O => \N__34454\,
            I => \N__34439\
        );

    \I__7796\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34434\
        );

    \I__7795\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34434\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__34449\,
            I => \N__34429\
        );

    \I__7793\ : InMux
    port map (
            O => \N__34446\,
            I => \N__34426\
        );

    \I__7792\ : CascadeMux
    port map (
            O => \N__34445\,
            I => \N__34423\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__34442\,
            I => \N__34418\
        );

    \I__7790\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34415\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34412\
        );

    \I__7788\ : InMux
    port map (
            O => \N__34433\,
            I => \N__34409\
        );

    \I__7787\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34406\
        );

    \I__7786\ : Span4Mux_v
    port map (
            O => \N__34429\,
            I => \N__34400\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__34426\,
            I => \N__34400\
        );

    \I__7784\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34397\
        );

    \I__7783\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34392\
        );

    \I__7782\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34389\
        );

    \I__7781\ : Span4Mux_v
    port map (
            O => \N__34418\,
            I => \N__34385\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__34415\,
            I => \N__34382\
        );

    \I__7779\ : Span4Mux_h
    port map (
            O => \N__34412\,
            I => \N__34375\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__34409\,
            I => \N__34375\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__34406\,
            I => \N__34375\
        );

    \I__7776\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34372\
        );

    \I__7775\ : Span4Mux_h
    port map (
            O => \N__34400\,
            I => \N__34369\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__34397\,
            I => \N__34366\
        );

    \I__7773\ : InMux
    port map (
            O => \N__34396\,
            I => \N__34363\
        );

    \I__7772\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34360\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34355\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__34389\,
            I => \N__34355\
        );

    \I__7769\ : InMux
    port map (
            O => \N__34388\,
            I => \N__34352\
        );

    \I__7768\ : Span4Mux_h
    port map (
            O => \N__34385\,
            I => \N__34343\
        );

    \I__7767\ : Span4Mux_v
    port map (
            O => \N__34382\,
            I => \N__34343\
        );

    \I__7766\ : Span4Mux_v
    port map (
            O => \N__34375\,
            I => \N__34343\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__34372\,
            I => \N__34343\
        );

    \I__7764\ : Sp12to4
    port map (
            O => \N__34369\,
            I => \N__34330\
        );

    \I__7763\ : Sp12to4
    port map (
            O => \N__34366\,
            I => \N__34330\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__34363\,
            I => \N__34330\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__34360\,
            I => \N__34330\
        );

    \I__7760\ : Sp12to4
    port map (
            O => \N__34355\,
            I => \N__34330\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34330\
        );

    \I__7758\ : Span4Mux_v
    port map (
            O => \N__34343\,
            I => \N__34327\
        );

    \I__7757\ : Span12Mux_v
    port map (
            O => \N__34330\,
            I => \N__34324\
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__34327\,
            I => gpio_fpga_soc_4
        );

    \I__7755\ : Odrv12
    port map (
            O => \N__34324\,
            I => gpio_fpga_soc_4
        );

    \I__7754\ : IoInMux
    port map (
            O => \N__34319\,
            I => \N__34316\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__34316\,
            I => \N__34313\
        );

    \I__7752\ : IoSpan4Mux
    port map (
            O => \N__34313\,
            I => \N__34308\
        );

    \I__7751\ : CascadeMux
    port map (
            O => \N__34312\,
            I => \N__34305\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__34311\,
            I => \N__34302\
        );

    \I__7749\ : IoSpan4Mux
    port map (
            O => \N__34308\,
            I => \N__34297\
        );

    \I__7748\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34294\
        );

    \I__7747\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34291\
        );

    \I__7746\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34281\
        );

    \I__7745\ : CascadeMux
    port map (
            O => \N__34300\,
            I => \N__34278\
        );

    \I__7744\ : Span4Mux_s3_v
    port map (
            O => \N__34297\,
            I => \N__34270\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__34294\,
            I => \N__34270\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__34291\,
            I => \N__34270\
        );

    \I__7741\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34265\
        );

    \I__7740\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34265\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__34288\,
            I => \N__34262\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__34287\,
            I => \N__34259\
        );

    \I__7737\ : CascadeMux
    port map (
            O => \N__34286\,
            I => \N__34256\
        );

    \I__7736\ : CascadeMux
    port map (
            O => \N__34285\,
            I => \N__34253\
        );

    \I__7735\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34245\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__34281\,
            I => \N__34242\
        );

    \I__7733\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34238\
        );

    \I__7732\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34235\
        );

    \I__7731\ : Span4Mux_v
    port map (
            O => \N__34270\,
            I => \N__34230\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__34265\,
            I => \N__34230\
        );

    \I__7729\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34225\
        );

    \I__7728\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34225\
        );

    \I__7727\ : InMux
    port map (
            O => \N__34256\,
            I => \N__34222\
        );

    \I__7726\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34216\
        );

    \I__7725\ : InMux
    port map (
            O => \N__34252\,
            I => \N__34211\
        );

    \I__7724\ : InMux
    port map (
            O => \N__34251\,
            I => \N__34211\
        );

    \I__7723\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34208\
        );

    \I__7722\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34205\
        );

    \I__7721\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34202\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__34245\,
            I => \N__34197\
        );

    \I__7719\ : Span4Mux_v
    port map (
            O => \N__34242\,
            I => \N__34194\
        );

    \I__7718\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34191\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__34238\,
            I => \N__34186\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__34235\,
            I => \N__34186\
        );

    \I__7715\ : Sp12to4
    port map (
            O => \N__34230\,
            I => \N__34183\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__34225\,
            I => \N__34178\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__34222\,
            I => \N__34175\
        );

    \I__7712\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34172\
        );

    \I__7711\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34169\
        );

    \I__7710\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34166\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__34216\,
            I => \N__34163\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__34211\,
            I => \N__34160\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__34208\,
            I => \N__34155\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__34205\,
            I => \N__34155\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34152\
        );

    \I__7704\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34149\
        );

    \I__7703\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34146\
        );

    \I__7702\ : Span12Mux_s8_v
    port map (
            O => \N__34197\,
            I => \N__34143\
        );

    \I__7701\ : Sp12to4
    port map (
            O => \N__34194\,
            I => \N__34134\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__34191\,
            I => \N__34134\
        );

    \I__7699\ : Span12Mux_s8_v
    port map (
            O => \N__34186\,
            I => \N__34134\
        );

    \I__7698\ : Span12Mux_s7_v
    port map (
            O => \N__34183\,
            I => \N__34134\
        );

    \I__7697\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34131\
        );

    \I__7696\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34128\
        );

    \I__7695\ : Span4Mux_h
    port map (
            O => \N__34178\,
            I => \N__34117\
        );

    \I__7694\ : Span4Mux_h
    port map (
            O => \N__34175\,
            I => \N__34117\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__34172\,
            I => \N__34117\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__34169\,
            I => \N__34117\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__34166\,
            I => \N__34117\
        );

    \I__7690\ : Span4Mux_h
    port map (
            O => \N__34163\,
            I => \N__34110\
        );

    \I__7689\ : Span4Mux_h
    port map (
            O => \N__34160\,
            I => \N__34110\
        );

    \I__7688\ : Span4Mux_s3_h
    port map (
            O => \N__34155\,
            I => \N__34110\
        );

    \I__7687\ : Span4Mux_s2_h
    port map (
            O => \N__34152\,
            I => \N__34107\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__34149\,
            I => \N__34102\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__34146\,
            I => \N__34102\
        );

    \I__7684\ : Odrv12
    port map (
            O => \N__34143\,
            I => rsmrstn
        );

    \I__7683\ : Odrv12
    port map (
            O => \N__34134\,
            I => rsmrstn
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__34131\,
            I => rsmrstn
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__34128\,
            I => rsmrstn
        );

    \I__7680\ : Odrv4
    port map (
            O => \N__34117\,
            I => rsmrstn
        );

    \I__7679\ : Odrv4
    port map (
            O => \N__34110\,
            I => rsmrstn
        );

    \I__7678\ : Odrv4
    port map (
            O => \N__34107\,
            I => rsmrstn
        );

    \I__7677\ : Odrv12
    port map (
            O => \N__34102\,
            I => rsmrstn
        );

    \I__7676\ : InMux
    port map (
            O => \N__34085\,
            I => \N__34082\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__34082\,
            I => \N__34079\
        );

    \I__7674\ : Span4Mux_v
    port map (
            O => \N__34079\,
            I => \N__34075\
        );

    \I__7673\ : InMux
    port map (
            O => \N__34078\,
            I => \N__34072\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__34075\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__34072\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0\
        );

    \I__7670\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34053\
        );

    \I__7669\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34049\
        );

    \I__7668\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34045\
        );

    \I__7667\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34042\
        );

    \I__7666\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34035\
        );

    \I__7665\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34035\
        );

    \I__7664\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34032\
        );

    \I__7663\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34027\
        );

    \I__7662\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34027\
        );

    \I__7661\ : InMux
    port map (
            O => \N__34058\,
            I => \N__34020\
        );

    \I__7660\ : InMux
    port map (
            O => \N__34057\,
            I => \N__34020\
        );

    \I__7659\ : InMux
    port map (
            O => \N__34056\,
            I => \N__34020\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__34053\,
            I => \N__34017\
        );

    \I__7657\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34011\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__34049\,
            I => \N__34008\
        );

    \I__7655\ : InMux
    port map (
            O => \N__34048\,
            I => \N__34005\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__34045\,
            I => \N__34000\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__34042\,
            I => \N__34000\
        );

    \I__7652\ : InMux
    port map (
            O => \N__34041\,
            I => \N__33995\
        );

    \I__7651\ : InMux
    port map (
            O => \N__34040\,
            I => \N__33995\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__34035\,
            I => \N__33990\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__34032\,
            I => \N__33990\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__33985\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__33985\
        );

    \I__7646\ : Span12Mux_s2_h
    port map (
            O => \N__34017\,
            I => \N__33982\
        );

    \I__7645\ : InMux
    port map (
            O => \N__34016\,
            I => \N__33979\
        );

    \I__7644\ : InMux
    port map (
            O => \N__34015\,
            I => \N__33976\
        );

    \I__7643\ : InMux
    port map (
            O => \N__34014\,
            I => \N__33973\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__34011\,
            I => \N__33970\
        );

    \I__7641\ : Span4Mux_h
    port map (
            O => \N__34008\,
            I => \N__33961\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__34005\,
            I => \N__33961\
        );

    \I__7639\ : Span4Mux_s3_h
    port map (
            O => \N__34000\,
            I => \N__33961\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__33995\,
            I => \N__33961\
        );

    \I__7637\ : Span4Mux_s2_h
    port map (
            O => \N__33990\,
            I => \N__33958\
        );

    \I__7636\ : Span4Mux_s2_h
    port map (
            O => \N__33985\,
            I => \N__33955\
        );

    \I__7635\ : Odrv12
    port map (
            O => \N__33982\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__33979\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__33976\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__33973\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7631\ : Odrv12
    port map (
            O => \N__33970\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__33961\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7629\ : Odrv4
    port map (
            O => \N__33958\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7628\ : Odrv4
    port map (
            O => \N__33955\,
            I => \b2v_inst11.N_2946_i\
        );

    \I__7627\ : CascadeMux
    port map (
            O => \N__33938\,
            I => \N__33934\
        );

    \I__7626\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33930\
        );

    \I__7625\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33925\
        );

    \I__7624\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33922\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33914\
        );

    \I__7622\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33909\
        );

    \I__7621\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33909\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33904\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__33922\,
            I => \N__33904\
        );

    \I__7618\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33899\
        );

    \I__7617\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33899\
        );

    \I__7616\ : InMux
    port map (
            O => \N__33919\,
            I => \N__33895\
        );

    \I__7615\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33892\
        );

    \I__7614\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33888\
        );

    \I__7613\ : Span4Mux_h
    port map (
            O => \N__33914\,
            I => \N__33874\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__33909\,
            I => \N__33874\
        );

    \I__7611\ : Span4Mux_h
    port map (
            O => \N__33904\,
            I => \N__33874\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33871\
        );

    \I__7609\ : InMux
    port map (
            O => \N__33898\,
            I => \N__33868\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__33895\,
            I => \N__33861\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__33892\,
            I => \N__33861\
        );

    \I__7606\ : InMux
    port map (
            O => \N__33891\,
            I => \N__33858\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__33888\,
            I => \N__33855\
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__33887\,
            I => \N__33851\
        );

    \I__7603\ : InMux
    port map (
            O => \N__33886\,
            I => \N__33837\
        );

    \I__7602\ : InMux
    port map (
            O => \N__33885\,
            I => \N__33837\
        );

    \I__7601\ : InMux
    port map (
            O => \N__33884\,
            I => \N__33832\
        );

    \I__7600\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33832\
        );

    \I__7599\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33827\
        );

    \I__7598\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33827\
        );

    \I__7597\ : Span4Mux_v
    port map (
            O => \N__33874\,
            I => \N__33824\
        );

    \I__7596\ : Span4Mux_v
    port map (
            O => \N__33871\,
            I => \N__33819\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__33868\,
            I => \N__33819\
        );

    \I__7594\ : InMux
    port map (
            O => \N__33867\,
            I => \N__33814\
        );

    \I__7593\ : InMux
    port map (
            O => \N__33866\,
            I => \N__33814\
        );

    \I__7592\ : Span4Mux_v
    port map (
            O => \N__33861\,
            I => \N__33811\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__33858\,
            I => \N__33808\
        );

    \I__7590\ : Span4Mux_v
    port map (
            O => \N__33855\,
            I => \N__33805\
        );

    \I__7589\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33796\
        );

    \I__7588\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33796\
        );

    \I__7587\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33796\
        );

    \I__7586\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33796\
        );

    \I__7585\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33793\
        );

    \I__7584\ : InMux
    port map (
            O => \N__33847\,
            I => \N__33786\
        );

    \I__7583\ : InMux
    port map (
            O => \N__33846\,
            I => \N__33786\
        );

    \I__7582\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33786\
        );

    \I__7581\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33779\
        );

    \I__7580\ : InMux
    port map (
            O => \N__33843\,
            I => \N__33779\
        );

    \I__7579\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33779\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33776\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__33832\,
            I => \N__33773\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33764\
        );

    \I__7575\ : Span4Mux_h
    port map (
            O => \N__33824\,
            I => \N__33764\
        );

    \I__7574\ : Span4Mux_h
    port map (
            O => \N__33819\,
            I => \N__33764\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__33814\,
            I => \N__33764\
        );

    \I__7572\ : Span4Mux_h
    port map (
            O => \N__33811\,
            I => \N__33759\
        );

    \I__7571\ : Span4Mux_v
    port map (
            O => \N__33808\,
            I => \N__33759\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__33805\,
            I => \N__33754\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__33796\,
            I => \N__33754\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33745\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__33786\,
            I => \N__33745\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__33779\,
            I => \N__33745\
        );

    \I__7565\ : Span12Mux_s5_v
    port map (
            O => \N__33776\,
            I => \N__33745\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__33773\,
            I => \N__33740\
        );

    \I__7563\ : Span4Mux_v
    port map (
            O => \N__33764\,
            I => \N__33740\
        );

    \I__7562\ : Odrv4
    port map (
            O => \N__33759\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\
        );

    \I__7561\ : Odrv4
    port map (
            O => \N__33754\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\
        );

    \I__7560\ : Odrv12
    port map (
            O => \N__33745\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\
        );

    \I__7559\ : Odrv4
    port map (
            O => \N__33740\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\
        );

    \I__7558\ : CascadeMux
    port map (
            O => \N__33731\,
            I => \N__33727\
        );

    \I__7557\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33723\
        );

    \I__7556\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33720\
        );

    \I__7555\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33717\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__33723\,
            I => \N__33711\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__33720\,
            I => \N__33711\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__33717\,
            I => \N__33708\
        );

    \I__7551\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33704\
        );

    \I__7550\ : Span4Mux_s0_h
    port map (
            O => \N__33711\,
            I => \N__33699\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__33708\,
            I => \N__33699\
        );

    \I__7548\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33696\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__33704\,
            I => \N__33693\
        );

    \I__7546\ : Span4Mux_h
    port map (
            O => \N__33699\,
            I => \N__33688\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__33696\,
            I => \N__33688\
        );

    \I__7544\ : Span4Mux_v
    port map (
            O => \N__33693\,
            I => \N__33685\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__33688\,
            I => \N__33682\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__33685\,
            I => \N__33679\
        );

    \I__7541\ : Odrv4
    port map (
            O => \N__33682\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_5\
        );

    \I__7540\ : Odrv4
    port map (
            O => \N__33679\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_5\
        );

    \I__7539\ : InMux
    port map (
            O => \N__33674\,
            I => \N__33671\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__33668\,
            I => \b2v_inst11.g0_1_1\
        );

    \I__7536\ : InMux
    port map (
            O => \N__33665\,
            I => \N__33662\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__33662\,
            I => \N__33659\
        );

    \I__7534\ : Span4Mux_v
    port map (
            O => \N__33659\,
            I => \N__33656\
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__33656\,
            I => vddq_ok
        );

    \I__7532\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33650\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33647\
        );

    \I__7530\ : Span4Mux_h
    port map (
            O => \N__33647\,
            I => \N__33643\
        );

    \I__7529\ : InMux
    port map (
            O => \N__33646\,
            I => \N__33640\
        );

    \I__7528\ : Span4Mux_v
    port map (
            O => \N__33643\,
            I => \N__33634\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__33640\,
            I => \N__33634\
        );

    \I__7526\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33629\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__33634\,
            I => \N__33626\
        );

    \I__7524\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33623\
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__33632\,
            I => \N__33619\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33614\
        );

    \I__7521\ : Span4Mux_h
    port map (
            O => \N__33626\,
            I => \N__33609\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__33623\,
            I => \N__33609\
        );

    \I__7519\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33606\
        );

    \I__7518\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33603\
        );

    \I__7517\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33600\
        );

    \I__7516\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33597\
        );

    \I__7515\ : Span12Mux_s3_h
    port map (
            O => \N__33614\,
            I => \N__33594\
        );

    \I__7514\ : Sp12to4
    port map (
            O => \N__33609\,
            I => \N__33583\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__33606\,
            I => \N__33583\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__33603\,
            I => \N__33583\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__33600\,
            I => \N__33583\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__33597\,
            I => \N__33583\
        );

    \I__7509\ : Odrv12
    port map (
            O => \N__33594\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__7508\ : Odrv12
    port map (
            O => \N__33583\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__7507\ : InMux
    port map (
            O => \N__33578\,
            I => \N__33573\
        );

    \I__7506\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33570\
        );

    \I__7505\ : InMux
    port map (
            O => \N__33576\,
            I => \N__33567\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__33573\,
            I => \N__33562\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__33570\,
            I => \N__33562\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__33567\,
            I => \N__33559\
        );

    \I__7501\ : Span4Mux_h
    port map (
            O => \N__33562\,
            I => \N__33556\
        );

    \I__7500\ : Sp12to4
    port map (
            O => \N__33559\,
            I => \N__33553\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__33556\,
            I => \N__33550\
        );

    \I__7498\ : Span12Mux_s10_v
    port map (
            O => \N__33553\,
            I => \N__33547\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__33550\,
            I => \N__33544\
        );

    \I__7496\ : Odrv12
    port map (
            O => \N__33547\,
            I => \b2v_inst16.N_208_0\
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__33544\,
            I => \b2v_inst16.N_208_0\
        );

    \I__7494\ : InMux
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__33536\,
            I => \b2v_inst11.count_off_1_1\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__33533\,
            I => \b2v_inst11.g0_13_1_cascade_\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__33530\,
            I => \b2v_inst11.N_4690_0_0_cascade_\
        );

    \I__7490\ : InMux
    port map (
            O => \N__33527\,
            I => \N__33524\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__33524\,
            I => \b2v_inst11.N_19_0\
        );

    \I__7488\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33518\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__33518\,
            I => \b2v_inst11.N_19_1\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__33515\,
            I => \N__33510\
        );

    \I__7485\ : CascadeMux
    port map (
            O => \N__33514\,
            I => \N__33505\
        );

    \I__7484\ : CascadeMux
    port map (
            O => \N__33513\,
            I => \N__33502\
        );

    \I__7483\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33495\
        );

    \I__7482\ : InMux
    port map (
            O => \N__33509\,
            I => \N__33495\
        );

    \I__7481\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33492\
        );

    \I__7480\ : InMux
    port map (
            O => \N__33505\,
            I => \N__33489\
        );

    \I__7479\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33484\
        );

    \I__7478\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33484\
        );

    \I__7477\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33481\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33478\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__33492\,
            I => \N__33474\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__33489\,
            I => \N__33471\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__33484\,
            I => \N__33468\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__33481\,
            I => \N__33464\
        );

    \I__7471\ : Span4Mux_s2_h
    port map (
            O => \N__33478\,
            I => \N__33461\
        );

    \I__7470\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33458\
        );

    \I__7469\ : Span4Mux_s3_h
    port map (
            O => \N__33474\,
            I => \N__33451\
        );

    \I__7468\ : Span4Mux_s3_h
    port map (
            O => \N__33471\,
            I => \N__33451\
        );

    \I__7467\ : Span4Mux_v
    port map (
            O => \N__33468\,
            I => \N__33451\
        );

    \I__7466\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33448\
        );

    \I__7465\ : Odrv12
    port map (
            O => \N__33464\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__33461\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__33458\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__33451\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__33448\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__7460\ : InMux
    port map (
            O => \N__33437\,
            I => \N__33434\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__33434\,
            I => \b2v_inst11.un1_dutycycle_172_m0\
        );

    \I__7458\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33428\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__33428\,
            I => \N__33425\
        );

    \I__7456\ : Span12Mux_s10_v
    port map (
            O => \N__33425\,
            I => \N__33422\
        );

    \I__7455\ : Odrv12
    port map (
            O => \N__33422\,
            I => \b2v_inst11.g3_3\
        );

    \I__7454\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33412\
        );

    \I__7453\ : InMux
    port map (
            O => \N__33418\,
            I => \N__33408\
        );

    \I__7452\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33403\
        );

    \I__7451\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33398\
        );

    \I__7450\ : InMux
    port map (
            O => \N__33415\,
            I => \N__33398\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__33412\,
            I => \N__33395\
        );

    \I__7448\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33392\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__33408\,
            I => \N__33389\
        );

    \I__7446\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33386\
        );

    \I__7445\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33381\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__33403\,
            I => \N__33372\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__33398\,
            I => \N__33372\
        );

    \I__7442\ : Span4Mux_v
    port map (
            O => \N__33395\,
            I => \N__33369\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__33392\,
            I => \N__33366\
        );

    \I__7440\ : Span4Mux_v
    port map (
            O => \N__33389\,
            I => \N__33361\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__33386\,
            I => \N__33361\
        );

    \I__7438\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33356\
        );

    \I__7437\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33356\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__33381\,
            I => \N__33353\
        );

    \I__7435\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33348\
        );

    \I__7434\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33348\
        );

    \I__7433\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33345\
        );

    \I__7432\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33342\
        );

    \I__7431\ : Span12Mux_s8_v
    port map (
            O => \N__33372\,
            I => \N__33339\
        );

    \I__7430\ : Span4Mux_v
    port map (
            O => \N__33369\,
            I => \N__33330\
        );

    \I__7429\ : Span4Mux_h
    port map (
            O => \N__33366\,
            I => \N__33330\
        );

    \I__7428\ : Span4Mux_v
    port map (
            O => \N__33361\,
            I => \N__33330\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33330\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__33353\,
            I => \N__33327\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__33348\,
            I => \b2v_inst11.N_172\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__33345\,
            I => \b2v_inst11.N_172\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__33342\,
            I => \b2v_inst11.N_172\
        );

    \I__7422\ : Odrv12
    port map (
            O => \N__33339\,
            I => \b2v_inst11.N_172\
        );

    \I__7421\ : Odrv4
    port map (
            O => \N__33330\,
            I => \b2v_inst11.N_172\
        );

    \I__7420\ : Odrv4
    port map (
            O => \N__33327\,
            I => \b2v_inst11.N_172\
        );

    \I__7419\ : CascadeMux
    port map (
            O => \N__33314\,
            I => \N__33308\
        );

    \I__7418\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33299\
        );

    \I__7417\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33299\
        );

    \I__7416\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33294\
        );

    \I__7415\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33294\
        );

    \I__7414\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33288\
        );

    \I__7413\ : InMux
    port map (
            O => \N__33306\,
            I => \N__33288\
        );

    \I__7412\ : InMux
    port map (
            O => \N__33305\,
            I => \N__33285\
        );

    \I__7411\ : InMux
    port map (
            O => \N__33304\,
            I => \N__33282\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__33299\,
            I => \N__33276\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__33294\,
            I => \N__33273\
        );

    \I__7408\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33270\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__33288\,
            I => \N__33267\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__33285\,
            I => \N__33264\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33261\
        );

    \I__7404\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33253\
        );

    \I__7403\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33253\
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__33279\,
            I => \N__33250\
        );

    \I__7401\ : Span4Mux_s1_h
    port map (
            O => \N__33276\,
            I => \N__33243\
        );

    \I__7400\ : Span4Mux_s1_h
    port map (
            O => \N__33273\,
            I => \N__33243\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__33270\,
            I => \N__33243\
        );

    \I__7398\ : Span12Mux_s5_h
    port map (
            O => \N__33267\,
            I => \N__33240\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__33264\,
            I => \N__33235\
        );

    \I__7396\ : Span4Mux_v
    port map (
            O => \N__33261\,
            I => \N__33235\
        );

    \I__7395\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33228\
        );

    \I__7394\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33228\
        );

    \I__7393\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33228\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__33253\,
            I => \N__33225\
        );

    \I__7391\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33222\
        );

    \I__7390\ : Span4Mux_h
    port map (
            O => \N__33243\,
            I => \N__33219\
        );

    \I__7389\ : Odrv12
    port map (
            O => \N__33240\,
            I => \b2v_inst11.N_200_i\
        );

    \I__7388\ : Odrv4
    port map (
            O => \N__33235\,
            I => \b2v_inst11.N_200_i\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__33228\,
            I => \b2v_inst11.N_200_i\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__33225\,
            I => \b2v_inst11.N_200_i\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__33222\,
            I => \b2v_inst11.N_200_i\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__33219\,
            I => \b2v_inst11.N_200_i\
        );

    \I__7383\ : InMux
    port map (
            O => \N__33206\,
            I => \N__33200\
        );

    \I__7382\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33200\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__33200\,
            I => \b2v_inst11.N_3099_0_0\
        );

    \I__7380\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33193\
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__33196\,
            I => \N__33188\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__33193\,
            I => \N__33183\
        );

    \I__7377\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33178\
        );

    \I__7376\ : InMux
    port map (
            O => \N__33191\,
            I => \N__33178\
        );

    \I__7375\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33175\
        );

    \I__7374\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33171\
        );

    \I__7373\ : CascadeMux
    port map (
            O => \N__33186\,
            I => \N__33167\
        );

    \I__7372\ : Span4Mux_s2_v
    port map (
            O => \N__33183\,
            I => \N__33162\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__33178\,
            I => \N__33157\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__33175\,
            I => \N__33157\
        );

    \I__7369\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33154\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__33171\,
            I => \N__33151\
        );

    \I__7367\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33147\
        );

    \I__7366\ : InMux
    port map (
            O => \N__33167\,
            I => \N__33141\
        );

    \I__7365\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33141\
        );

    \I__7364\ : InMux
    port map (
            O => \N__33165\,
            I => \N__33138\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__33162\,
            I => \N__33131\
        );

    \I__7362\ : Span4Mux_v
    port map (
            O => \N__33157\,
            I => \N__33131\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__33154\,
            I => \N__33131\
        );

    \I__7360\ : Span4Mux_h
    port map (
            O => \N__33151\,
            I => \N__33128\
        );

    \I__7359\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33125\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__33147\,
            I => \N__33122\
        );

    \I__7357\ : InMux
    port map (
            O => \N__33146\,
            I => \N__33119\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__33141\,
            I => \N__33114\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__33138\,
            I => \N__33114\
        );

    \I__7354\ : Span4Mux_h
    port map (
            O => \N__33131\,
            I => \N__33111\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__33128\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__33125\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__7351\ : Odrv4
    port map (
            O => \N__33122\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__33119\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__7349\ : Odrv12
    port map (
            O => \N__33114\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__7348\ : Odrv4
    port map (
            O => \N__33111\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__7347\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33095\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__7345\ : Span4Mux_v
    port map (
            O => \N__33092\,
            I => \N__33089\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__33089\,
            I => \b2v_inst11.N_237\
        );

    \I__7343\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33083\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__33083\,
            I => \b2v_inst11.N_293_0_0\
        );

    \I__7341\ : CascadeMux
    port map (
            O => \N__33080\,
            I => \N__33075\
        );

    \I__7340\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33071\
        );

    \I__7339\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33068\
        );

    \I__7338\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33065\
        );

    \I__7337\ : CascadeMux
    port map (
            O => \N__33074\,
            I => \N__33062\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__33071\,
            I => \N__33059\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__33068\,
            I => \N__33056\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__33065\,
            I => \N__33053\
        );

    \I__7333\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33050\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__33059\,
            I => \N__33046\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__33056\,
            I => \N__33039\
        );

    \I__7330\ : Span4Mux_s1_h
    port map (
            O => \N__33053\,
            I => \N__33039\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__33050\,
            I => \N__33039\
        );

    \I__7328\ : InMux
    port map (
            O => \N__33049\,
            I => \N__33036\
        );

    \I__7327\ : Span4Mux_v
    port map (
            O => \N__33046\,
            I => \N__33033\
        );

    \I__7326\ : Span4Mux_h
    port map (
            O => \N__33039\,
            I => \N__33028\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__33036\,
            I => \N__33028\
        );

    \I__7324\ : Odrv4
    port map (
            O => \N__33033\,
            I => \b2v_inst11.count_clk_RNIZ0Z_6\
        );

    \I__7323\ : Odrv4
    port map (
            O => \N__33028\,
            I => \b2v_inst11.count_clk_RNIZ0Z_6\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__33023\,
            I => \N__33020\
        );

    \I__7321\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33014\
        );

    \I__7320\ : InMux
    port map (
            O => \N__33019\,
            I => \N__33014\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__33014\,
            I => \b2v_inst11.g2_1_0\
        );

    \I__7318\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33008\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__33008\,
            I => v5s_ok
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__33005\,
            I => \N__33002\
        );

    \I__7315\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32999\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__32999\,
            I => \N__32996\
        );

    \I__7313\ : Span12Mux_v
    port map (
            O => \N__32996\,
            I => \N__32993\
        );

    \I__7312\ : Odrv12
    port map (
            O => \N__32993\,
            I => v33s_ok
        );

    \I__7311\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32983\
        );

    \I__7310\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32976\
        );

    \I__7309\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32976\
        );

    \I__7308\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32976\
        );

    \I__7307\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32973\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__32983\,
            I => \N__32965\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__32976\,
            I => \N__32965\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__32973\,
            I => \N__32965\
        );

    \I__7303\ : InMux
    port map (
            O => \N__32972\,
            I => \N__32962\
        );

    \I__7302\ : Span4Mux_v
    port map (
            O => \N__32965\,
            I => \N__32959\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__32962\,
            I => \N__32956\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__32959\,
            I => \SYNTHESIZED_WIRE_8\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__32956\,
            I => \SYNTHESIZED_WIRE_8\
        );

    \I__7298\ : IoInMux
    port map (
            O => \N__32951\,
            I => \N__32948\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__32948\,
            I => \N__32945\
        );

    \I__7296\ : Span4Mux_s2_v
    port map (
            O => \N__32945\,
            I => \N__32942\
        );

    \I__7295\ : Sp12to4
    port map (
            O => \N__32942\,
            I => \N__32939\
        );

    \I__7294\ : Span12Mux_s11_h
    port map (
            O => \N__32939\,
            I => \N__32935\
        );

    \I__7293\ : IoInMux
    port map (
            O => \N__32938\,
            I => \N__32932\
        );

    \I__7292\ : Odrv12
    port map (
            O => \N__32935\,
            I => vccinaux_en
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__32932\,
            I => vccinaux_en
        );

    \I__7290\ : InMux
    port map (
            O => \N__32927\,
            I => \N__32924\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__32924\,
            I => \N__32921\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__32921\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_0\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__32918\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_0_cascade_\
        );

    \I__7286\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32912\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__32912\,
            I => \N__32901\
        );

    \I__7284\ : CascadeMux
    port map (
            O => \N__32911\,
            I => \N__32898\
        );

    \I__7283\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32891\
        );

    \I__7282\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32888\
        );

    \I__7281\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32881\
        );

    \I__7280\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32881\
        );

    \I__7279\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32881\
        );

    \I__7278\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32876\
        );

    \I__7277\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32876\
        );

    \I__7276\ : Span4Mux_v
    port map (
            O => \N__32901\,
            I => \N__32870\
        );

    \I__7275\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32865\
        );

    \I__7274\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32865\
        );

    \I__7273\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32862\
        );

    \I__7272\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32859\
        );

    \I__7271\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32856\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__32891\,
            I => \N__32847\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32847\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32847\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32847\
        );

    \I__7266\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32842\
        );

    \I__7265\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32842\
        );

    \I__7264\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32839\
        );

    \I__7263\ : Span4Mux_v
    port map (
            O => \N__32870\,
            I => \N__32836\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32833\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__32862\,
            I => \N__32828\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__32859\,
            I => \N__32828\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__32856\,
            I => \N__32825\
        );

    \I__7258\ : Span4Mux_v
    port map (
            O => \N__32847\,
            I => \N__32820\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__32842\,
            I => \N__32817\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__32839\,
            I => \N__32814\
        );

    \I__7255\ : Span4Mux_h
    port map (
            O => \N__32836\,
            I => \N__32808\
        );

    \I__7254\ : Span4Mux_v
    port map (
            O => \N__32833\,
            I => \N__32808\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__32828\,
            I => \N__32803\
        );

    \I__7252\ : Span4Mux_v
    port map (
            O => \N__32825\,
            I => \N__32803\
        );

    \I__7251\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32800\
        );

    \I__7250\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32797\
        );

    \I__7249\ : Span4Mux_v
    port map (
            O => \N__32820\,
            I => \N__32792\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__32817\,
            I => \N__32792\
        );

    \I__7247\ : Span4Mux_v
    port map (
            O => \N__32814\,
            I => \N__32789\
        );

    \I__7246\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32786\
        );

    \I__7245\ : Span4Mux_h
    port map (
            O => \N__32808\,
            I => \N__32783\
        );

    \I__7244\ : Sp12to4
    port map (
            O => \N__32803\,
            I => \N__32770\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__32800\,
            I => \N__32770\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__32797\,
            I => \N__32770\
        );

    \I__7241\ : Sp12to4
    port map (
            O => \N__32792\,
            I => \N__32770\
        );

    \I__7240\ : Sp12to4
    port map (
            O => \N__32789\,
            I => \N__32770\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__32786\,
            I => \N__32770\
        );

    \I__7238\ : Sp12to4
    port map (
            O => \N__32783\,
            I => \N__32765\
        );

    \I__7237\ : Span12Mux_s8_h
    port map (
            O => \N__32770\,
            I => \N__32765\
        );

    \I__7236\ : Odrv12
    port map (
            O => \N__32765\,
            I => slp_s4n
        );

    \I__7235\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32756\
        );

    \I__7234\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32756\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__32756\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_0\
        );

    \I__7232\ : CascadeMux
    port map (
            O => \N__32753\,
            I => \b2v_inst11.un1_dutycycle_172_m1_ns_1_cascade_\
        );

    \I__7231\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32747\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__32747\,
            I => \b2v_inst11.un1_dutycycle_172_m1\
        );

    \I__7229\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32741\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__32741\,
            I => \b2v_inst11.g0_i_2\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__32738\,
            I => \b2v_inst11.g0_0_0Z0Z_0_cascade_\
        );

    \I__7226\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32732\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__32732\,
            I => \b2v_inst6.count_1_i_a3_7_0\
        );

    \I__7224\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__32726\,
            I => \N__32723\
        );

    \I__7222\ : Odrv12
    port map (
            O => \N__32723\,
            I => \b2v_inst6.count_1_i_a3_1_0\
        );

    \I__7221\ : CascadeMux
    port map (
            O => \N__32720\,
            I => \b2v_inst6.count_1_i_a3_12_0_cascade_\
        );

    \I__7220\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32714\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__32714\,
            I => \b2v_inst6.count_1_i_a3_2_0\
        );

    \I__7218\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32705\
        );

    \I__7217\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32705\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__32705\,
            I => \b2v_inst6.N_389\
        );

    \I__7215\ : CascadeMux
    port map (
            O => \N__32702\,
            I => \b2v_inst6.N_389_cascade_\
        );

    \I__7214\ : InMux
    port map (
            O => \N__32699\,
            I => \N__32696\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__32696\,
            I => \b2v_inst6.count_0_0\
        );

    \I__7212\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__32690\,
            I => \b2v_inst6.count_rst_13\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__32687\,
            I => \N__32684\
        );

    \I__7209\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32677\
        );

    \I__7207\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32674\
        );

    \I__7206\ : Span4Mux_s0_v
    port map (
            O => \N__32677\,
            I => \N__32671\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__32674\,
            I => \b2v_inst6.un2_count_1_axb_1\
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__32671\,
            I => \b2v_inst6.un2_count_1_axb_1\
        );

    \I__7203\ : CascadeMux
    port map (
            O => \N__32666\,
            I => \b2v_inst6.un2_count_1_axb_1_cascade_\
        );

    \I__7202\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32659\
        );

    \I__7201\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32656\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__32659\,
            I => \b2v_inst6.count_0_1\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__32656\,
            I => \b2v_inst6.count_0_1\
        );

    \I__7198\ : SRMux
    port map (
            O => \N__32651\,
            I => \N__32645\
        );

    \I__7197\ : SRMux
    port map (
            O => \N__32650\,
            I => \N__32642\
        );

    \I__7196\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32636\
        );

    \I__7195\ : SRMux
    port map (
            O => \N__32648\,
            I => \N__32636\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__32645\,
            I => \N__32630\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__32642\,
            I => \N__32630\
        );

    \I__7192\ : SRMux
    port map (
            O => \N__32641\,
            I => \N__32627\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__32636\,
            I => \N__32604\
        );

    \I__7190\ : SRMux
    port map (
            O => \N__32635\,
            I => \N__32601\
        );

    \I__7189\ : Span4Mux_s2_v
    port map (
            O => \N__32630\,
            I => \N__32596\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__32627\,
            I => \N__32596\
        );

    \I__7187\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32585\
        );

    \I__7186\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32585\
        );

    \I__7185\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32585\
        );

    \I__7184\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32585\
        );

    \I__7183\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32585\
        );

    \I__7182\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32577\
        );

    \I__7181\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32577\
        );

    \I__7180\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32570\
        );

    \I__7179\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32570\
        );

    \I__7178\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32570\
        );

    \I__7177\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32567\
        );

    \I__7176\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32562\
        );

    \I__7175\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32562\
        );

    \I__7174\ : SRMux
    port map (
            O => \N__32613\,
            I => \N__32549\
        );

    \I__7173\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32549\
        );

    \I__7172\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32549\
        );

    \I__7171\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32549\
        );

    \I__7170\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32549\
        );

    \I__7169\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32549\
        );

    \I__7168\ : SRMux
    port map (
            O => \N__32607\,
            I => \N__32544\
        );

    \I__7167\ : Span4Mux_v
    port map (
            O => \N__32604\,
            I => \N__32536\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__32601\,
            I => \N__32536\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__32596\,
            I => \N__32531\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__32585\,
            I => \N__32531\
        );

    \I__7163\ : InMux
    port map (
            O => \N__32584\,
            I => \N__32524\
        );

    \I__7162\ : InMux
    port map (
            O => \N__32583\,
            I => \N__32524\
        );

    \I__7161\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32524\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__32577\,
            I => \N__32517\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32517\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__32567\,
            I => \N__32517\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__32562\,
            I => \N__32512\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32512\
        );

    \I__7155\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32507\
        );

    \I__7154\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32507\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__32544\,
            I => \N__32504\
        );

    \I__7152\ : InMux
    port map (
            O => \N__32543\,
            I => \N__32497\
        );

    \I__7151\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32497\
        );

    \I__7150\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32497\
        );

    \I__7149\ : Span4Mux_s2_v
    port map (
            O => \N__32536\,
            I => \N__32490\
        );

    \I__7148\ : Span4Mux_s2_v
    port map (
            O => \N__32531\,
            I => \N__32490\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__32524\,
            I => \N__32490\
        );

    \I__7146\ : Span4Mux_s2_v
    port map (
            O => \N__32517\,
            I => \N__32483\
        );

    \I__7145\ : Span4Mux_s1_h
    port map (
            O => \N__32512\,
            I => \N__32483\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__32507\,
            I => \N__32483\
        );

    \I__7143\ : Odrv12
    port map (
            O => \N__32504\,
            I => \b2v_inst6.curr_state_RNIM6FE1Z0Z_1\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__32497\,
            I => \b2v_inst6.curr_state_RNIM6FE1Z0Z_1\
        );

    \I__7141\ : Odrv4
    port map (
            O => \N__32490\,
            I => \b2v_inst6.curr_state_RNIM6FE1Z0Z_1\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__32483\,
            I => \b2v_inst6.curr_state_RNIM6FE1Z0Z_1\
        );

    \I__7139\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32471\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__32471\,
            I => \b2v_inst6.count_rst_5\
        );

    \I__7137\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32464\
        );

    \I__7136\ : InMux
    port map (
            O => \N__32467\,
            I => \N__32461\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__32464\,
            I => \b2v_inst6.count_0_9\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__32461\,
            I => \b2v_inst6.count_0_9\
        );

    \I__7133\ : CascadeMux
    port map (
            O => \N__32456\,
            I => \N__32452\
        );

    \I__7132\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32448\
        );

    \I__7131\ : InMux
    port map (
            O => \N__32452\,
            I => \N__32445\
        );

    \I__7130\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32442\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32439\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__32445\,
            I => \b2v_inst6.countZ0Z_8\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__32442\,
            I => \b2v_inst6.countZ0Z_8\
        );

    \I__7126\ : Odrv12
    port map (
            O => \N__32439\,
            I => \b2v_inst6.countZ0Z_8\
        );

    \I__7125\ : CEMux
    port map (
            O => \N__32432\,
            I => \N__32424\
        );

    \I__7124\ : CascadeMux
    port map (
            O => \N__32431\,
            I => \N__32419\
        );

    \I__7123\ : CEMux
    port map (
            O => \N__32430\,
            I => \N__32416\
        );

    \I__7122\ : CEMux
    port map (
            O => \N__32429\,
            I => \N__32413\
        );

    \I__7121\ : CEMux
    port map (
            O => \N__32428\,
            I => \N__32410\
        );

    \I__7120\ : CEMux
    port map (
            O => \N__32427\,
            I => \N__32407\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__32424\,
            I => \N__32404\
        );

    \I__7118\ : CEMux
    port map (
            O => \N__32423\,
            I => \N__32401\
        );

    \I__7117\ : CEMux
    port map (
            O => \N__32422\,
            I => \N__32398\
        );

    \I__7116\ : InMux
    port map (
            O => \N__32419\,
            I => \N__32393\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__32416\,
            I => \N__32390\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__32413\,
            I => \N__32383\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__32410\,
            I => \N__32383\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32383\
        );

    \I__7111\ : Span4Mux_s0_v
    port map (
            O => \N__32404\,
            I => \N__32378\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__32401\,
            I => \N__32378\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__32398\,
            I => \N__32369\
        );

    \I__7108\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32353\
        );

    \I__7107\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32353\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__32393\,
            I => \N__32344\
        );

    \I__7105\ : IoSpan4Mux
    port map (
            O => \N__32390\,
            I => \N__32344\
        );

    \I__7104\ : Span4Mux_v
    port map (
            O => \N__32383\,
            I => \N__32344\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__32378\,
            I => \N__32344\
        );

    \I__7102\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32333\
        );

    \I__7101\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32333\
        );

    \I__7100\ : InMux
    port map (
            O => \N__32375\,
            I => \N__32333\
        );

    \I__7099\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32333\
        );

    \I__7098\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32333\
        );

    \I__7097\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32327\
        );

    \I__7096\ : Span4Mux_s1_v
    port map (
            O => \N__32369\,
            I => \N__32324\
        );

    \I__7095\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32317\
        );

    \I__7094\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32317\
        );

    \I__7093\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32317\
        );

    \I__7092\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32312\
        );

    \I__7091\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32312\
        );

    \I__7090\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32303\
        );

    \I__7089\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32303\
        );

    \I__7088\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32303\
        );

    \I__7087\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32303\
        );

    \I__7086\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32298\
        );

    \I__7085\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32298\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__32353\,
            I => \N__32295\
        );

    \I__7083\ : Span4Mux_s0_v
    port map (
            O => \N__32344\,
            I => \N__32290\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__32333\,
            I => \N__32290\
        );

    \I__7081\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32283\
        );

    \I__7080\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32283\
        );

    \I__7079\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32283\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__32327\,
            I => \b2v_inst6.count_en\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__32324\,
            I => \b2v_inst6.count_en\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__32317\,
            I => \b2v_inst6.count_en\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__32312\,
            I => \b2v_inst6.count_en\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__32303\,
            I => \b2v_inst6.count_en\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__32298\,
            I => \b2v_inst6.count_en\
        );

    \I__7072\ : Odrv4
    port map (
            O => \N__32295\,
            I => \b2v_inst6.count_en\
        );

    \I__7071\ : Odrv4
    port map (
            O => \N__32290\,
            I => \b2v_inst6.count_en\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__32283\,
            I => \b2v_inst6.count_en\
        );

    \I__7069\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__32261\,
            I => \N__32258\
        );

    \I__7067\ : Odrv4
    port map (
            O => \N__32258\,
            I => \b2v_inst6.count_1_i_a3_4_0\
        );

    \I__7066\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32252\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__32252\,
            I => \N__32249\
        );

    \I__7064\ : Span4Mux_v
    port map (
            O => \N__32249\,
            I => \N__32245\
        );

    \I__7063\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32242\
        );

    \I__7062\ : Odrv4
    port map (
            O => \N__32245\,
            I => \b2v_inst5.N_51\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__32242\,
            I => \b2v_inst5.N_51\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__32237\,
            I => \N__32234\
        );

    \I__7059\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32231\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__32231\,
            I => \N__32228\
        );

    \I__7057\ : Odrv12
    port map (
            O => \N__32228\,
            I => \b2v_inst5.curr_state_0_1\
        );

    \I__7056\ : CascadeMux
    port map (
            O => \N__32225\,
            I => \N__32216\
        );

    \I__7055\ : CascadeMux
    port map (
            O => \N__32224\,
            I => \N__32211\
        );

    \I__7054\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32208\
        );

    \I__7053\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32205\
        );

    \I__7052\ : InMux
    port map (
            O => \N__32221\,
            I => \N__32202\
        );

    \I__7051\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32199\
        );

    \I__7050\ : InMux
    port map (
            O => \N__32219\,
            I => \N__32196\
        );

    \I__7049\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32191\
        );

    \I__7048\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32191\
        );

    \I__7047\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32188\
        );

    \I__7046\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32185\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32170\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32167\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__32202\,
            I => \N__32164\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__32199\,
            I => \N__32161\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__32196\,
            I => \N__32158\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32155\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__32188\,
            I => \N__32152\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__32185\,
            I => \N__32149\
        );

    \I__7037\ : CEMux
    port map (
            O => \N__32184\,
            I => \N__32108\
        );

    \I__7036\ : CEMux
    port map (
            O => \N__32183\,
            I => \N__32108\
        );

    \I__7035\ : CEMux
    port map (
            O => \N__32182\,
            I => \N__32108\
        );

    \I__7034\ : CEMux
    port map (
            O => \N__32181\,
            I => \N__32108\
        );

    \I__7033\ : CEMux
    port map (
            O => \N__32180\,
            I => \N__32108\
        );

    \I__7032\ : CEMux
    port map (
            O => \N__32179\,
            I => \N__32108\
        );

    \I__7031\ : CEMux
    port map (
            O => \N__32178\,
            I => \N__32108\
        );

    \I__7030\ : CEMux
    port map (
            O => \N__32177\,
            I => \N__32108\
        );

    \I__7029\ : CEMux
    port map (
            O => \N__32176\,
            I => \N__32108\
        );

    \I__7028\ : CEMux
    port map (
            O => \N__32175\,
            I => \N__32108\
        );

    \I__7027\ : CEMux
    port map (
            O => \N__32174\,
            I => \N__32108\
        );

    \I__7026\ : CEMux
    port map (
            O => \N__32173\,
            I => \N__32108\
        );

    \I__7025\ : Glb2LocalMux
    port map (
            O => \N__32170\,
            I => \N__32108\
        );

    \I__7024\ : Glb2LocalMux
    port map (
            O => \N__32167\,
            I => \N__32108\
        );

    \I__7023\ : Glb2LocalMux
    port map (
            O => \N__32164\,
            I => \N__32108\
        );

    \I__7022\ : Glb2LocalMux
    port map (
            O => \N__32161\,
            I => \N__32108\
        );

    \I__7021\ : Glb2LocalMux
    port map (
            O => \N__32158\,
            I => \N__32108\
        );

    \I__7020\ : Glb2LocalMux
    port map (
            O => \N__32155\,
            I => \N__32108\
        );

    \I__7019\ : Glb2LocalMux
    port map (
            O => \N__32152\,
            I => \N__32108\
        );

    \I__7018\ : Glb2LocalMux
    port map (
            O => \N__32149\,
            I => \N__32108\
        );

    \I__7017\ : GlobalMux
    port map (
            O => \N__32108\,
            I => \N__32105\
        );

    \I__7016\ : gio2CtrlBuf
    port map (
            O => \N__32105\,
            I => \N_606_g\
        );

    \I__7015\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32097\
        );

    \I__7014\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32094\
        );

    \I__7013\ : InMux
    port map (
            O => \N__32100\,
            I => \N__32091\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__32097\,
            I => \N__32088\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__32094\,
            I => \N__32085\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__32091\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7009\ : Odrv4
    port map (
            O => \N__32088\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7008\ : Odrv4
    port map (
            O => \N__32085\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7007\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32073\
        );

    \I__7006\ : InMux
    port map (
            O => \N__32077\,
            I => \N__32068\
        );

    \I__7005\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32068\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__32073\,
            I => \N__32063\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__32068\,
            I => \N__32063\
        );

    \I__7002\ : Odrv4
    port map (
            O => \N__32063\,
            I => \b2v_inst6.N_3036_i\
        );

    \I__7001\ : IoInMux
    port map (
            O => \N__32060\,
            I => \N__32056\
        );

    \I__7000\ : CascadeMux
    port map (
            O => \N__32059\,
            I => \N__32053\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__32056\,
            I => \N__32049\
        );

    \I__6998\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32043\
        );

    \I__6997\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32043\
        );

    \I__6996\ : Span4Mux_s3_h
    port map (
            O => \N__32049\,
            I => \N__32040\
        );

    \I__6995\ : InMux
    port map (
            O => \N__32048\,
            I => \N__32037\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__32034\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__32040\,
            I => \N__32029\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__32029\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__32034\,
            I => \N__32024\
        );

    \I__6990\ : Span4Mux_h
    port map (
            O => \N__32029\,
            I => \N__32024\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__32024\,
            I => \N__32021\
        );

    \I__6988\ : Odrv4
    port map (
            O => \N__32021\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__32018\,
            I => \b2v_inst6.count_rst_9_cascade_\
        );

    \I__6986\ : InMux
    port map (
            O => \N__32015\,
            I => \N__32010\
        );

    \I__6985\ : InMux
    port map (
            O => \N__32014\,
            I => \N__32007\
        );

    \I__6984\ : InMux
    port map (
            O => \N__32013\,
            I => \N__32004\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__32010\,
            I => \N__32001\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__32007\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__32004\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__32001\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__6979\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31988\
        );

    \I__6978\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31988\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31985\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__31985\,
            I => \b2v_inst6.un2_count_1_cry_4_THRU_CO\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__31982\,
            I => \b2v_inst6.countZ0Z_5_cascade_\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31976\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__31976\,
            I => \b2v_inst6.count_0_5\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__31973\,
            I => \N__31970\
        );

    \I__6971\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31967\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__31967\,
            I => \N__31963\
        );

    \I__6969\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31960\
        );

    \I__6968\ : Odrv4
    port map (
            O => \N__31963\,
            I => \b2v_inst6.un2_count_1_cry_10_THRU_CO\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__31960\,
            I => \b2v_inst6.un2_count_1_cry_10_THRU_CO\
        );

    \I__6966\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31936\
        );

    \I__6965\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31936\
        );

    \I__6964\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31931\
        );

    \I__6963\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31931\
        );

    \I__6962\ : InMux
    port map (
            O => \N__31951\,
            I => \N__31924\
        );

    \I__6961\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31924\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31924\
        );

    \I__6959\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31912\
        );

    \I__6958\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31912\
        );

    \I__6957\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31912\
        );

    \I__6956\ : InMux
    port map (
            O => \N__31945\,
            I => \N__31912\
        );

    \I__6955\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31912\
        );

    \I__6954\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31909\
        );

    \I__6953\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31904\
        );

    \I__6952\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31904\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__31936\,
            I => \N__31897\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31897\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__31924\,
            I => \N__31897\
        );

    \I__6948\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31894\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__31912\,
            I => \N__31891\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__31909\,
            I => \N__31884\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__31904\,
            I => \N__31884\
        );

    \I__6944\ : Span4Mux_v
    port map (
            O => \N__31897\,
            I => \N__31884\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__31894\,
            I => \b2v_inst6.N_394\
        );

    \I__6942\ : Odrv4
    port map (
            O => \N__31891\,
            I => \b2v_inst6.N_394\
        );

    \I__6941\ : Odrv4
    port map (
            O => \N__31884\,
            I => \b2v_inst6.N_394\
        );

    \I__6940\ : CascadeMux
    port map (
            O => \N__31877\,
            I => \b2v_inst6.count_rst_3_cascade_\
        );

    \I__6939\ : InMux
    port map (
            O => \N__31874\,
            I => \N__31871\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__31871\,
            I => \N__31868\
        );

    \I__6937\ : Odrv4
    port map (
            O => \N__31868\,
            I => \b2v_inst6.count_0_11\
        );

    \I__6936\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31862\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__31862\,
            I => \b2v_inst6.count_RNIM6FE1Z0Z_0\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__31859\,
            I => \b2v_inst6.countZ0Z_0_cascade_\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__31856\,
            I => \N__31851\
        );

    \I__6932\ : InMux
    port map (
            O => \N__31855\,
            I => \N__31848\
        );

    \I__6931\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31844\
        );

    \I__6930\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31841\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__31848\,
            I => \N__31838\
        );

    \I__6928\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31835\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__31844\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__31841\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6925\ : Odrv12
    port map (
            O => \N__31838\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__31835\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6923\ : CascadeMux
    port map (
            O => \N__31826\,
            I => \b2v_inst6.count_rst_13_cascade_\
        );

    \I__6922\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31820\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31817\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__31817\,
            I => \b2v_inst6.count_1_i_a3_5_0\
        );

    \I__6919\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31808\
        );

    \I__6917\ : Odrv12
    port map (
            O => \N__31808\,
            I => \b2v_inst6.count_1_i_a3_6_0\
        );

    \I__6916\ : CascadeMux
    port map (
            O => \N__31805\,
            I => \b2v_inst6.count_1_i_a3_3_0_cascade_\
        );

    \I__6915\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31799\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__31799\,
            I => \b2v_inst6.count_0_14\
        );

    \I__6913\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31790\
        );

    \I__6912\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31790\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__31790\,
            I => \b2v_inst6.un2_count_1_cry_13_c_RNI06SPZ0Z1\
        );

    \I__6910\ : InMux
    port map (
            O => \N__31787\,
            I => \N__31784\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__31784\,
            I => \b2v_inst6.countZ0Z_14\
        );

    \I__6908\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31777\
        );

    \I__6907\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31774\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__31777\,
            I => \b2v_inst6.count_0_2\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__31774\,
            I => \b2v_inst6.count_0_2\
        );

    \I__6904\ : CascadeMux
    port map (
            O => \N__31769\,
            I => \b2v_inst6.countZ0Z_14_cascade_\
        );

    \I__6903\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31757\
        );

    \I__6902\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31757\
        );

    \I__6901\ : InMux
    port map (
            O => \N__31764\,
            I => \N__31757\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__31757\,
            I => \b2v_inst6.count_rst_12\
        );

    \I__6899\ : InMux
    port map (
            O => \N__31754\,
            I => \N__31751\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__31751\,
            I => \b2v_inst6.un2_count_1_axb_12\
        );

    \I__6897\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31745\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__31745\,
            I => \N__31740\
        );

    \I__6895\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31735\
        );

    \I__6894\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31735\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__31740\,
            I => \b2v_inst6.count_rst_2\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__31735\,
            I => \b2v_inst6.count_rst_2\
        );

    \I__6891\ : InMux
    port map (
            O => \N__31730\,
            I => \N__31727\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__31727\,
            I => \N__31724\
        );

    \I__6889\ : Span4Mux_v
    port map (
            O => \N__31724\,
            I => \N__31720\
        );

    \I__6888\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31717\
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__31720\,
            I => \b2v_inst6.count_0_12\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__31717\,
            I => \b2v_inst6.count_0_12\
        );

    \I__6885\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31705\
        );

    \I__6884\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31705\
        );

    \I__6883\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31702\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__31705\,
            I => \b2v_inst6.count_rst_1\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__31702\,
            I => \b2v_inst6.count_rst_1\
        );

    \I__6880\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31693\
        );

    \I__6879\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31690\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__31693\,
            I => \N__31687\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__31690\,
            I => \b2v_inst6.count_0_13\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__31687\,
            I => \b2v_inst6.count_0_13\
        );

    \I__6875\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31679\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__31679\,
            I => \b2v_inst6.un2_count_1_axb_13\
        );

    \I__6873\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31673\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31669\
        );

    \I__6871\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31666\
        );

    \I__6870\ : Span4Mux_s1_h
    port map (
            O => \N__31669\,
            I => \N__31663\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__31666\,
            I => \N__31660\
        );

    \I__6868\ : Odrv4
    port map (
            O => \N__31663\,
            I => \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__31660\,
            I => \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\
        );

    \I__6866\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31652\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__31652\,
            I => \b2v_inst6.count_0_6\
        );

    \I__6864\ : CascadeMux
    port map (
            O => \N__31649\,
            I => \b2v_inst6.N_394_cascade_\
        );

    \I__6863\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31640\
        );

    \I__6862\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31640\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__31640\,
            I => \b2v_inst6.un2_count_1_cry_3_THRU_CO\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__31637\,
            I => \b2v_inst6.un2_count_1_axb_4_cascade_\
        );

    \I__6859\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31631\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__31631\,
            I => \b2v_inst6.count_rst_10\
        );

    \I__6857\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31622\
        );

    \I__6856\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31622\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__31622\,
            I => \b2v_inst6.count_0_4\
        );

    \I__6854\ : CascadeMux
    port map (
            O => \N__31619\,
            I => \b2v_inst6.count_rst_11_cascade_\
        );

    \I__6853\ : CascadeMux
    port map (
            O => \N__31616\,
            I => \N__31612\
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__31615\,
            I => \N__31608\
        );

    \I__6851\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31605\
        );

    \I__6850\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31602\
        );

    \I__6849\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31599\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__31605\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__31602\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__31599\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__6845\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31586\
        );

    \I__6844\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31586\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__31586\,
            I => \b2v_inst6.un2_count_1_cry_2_THRU_CO\
        );

    \I__6842\ : CascadeMux
    port map (
            O => \N__31583\,
            I => \b2v_inst6.countZ0Z_3_cascade_\
        );

    \I__6841\ : InMux
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__31577\,
            I => \b2v_inst6.count_0_3\
        );

    \I__6839\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31571\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__31571\,
            I => \b2v_inst6.un2_count_1_axb_2\
        );

    \I__6837\ : InMux
    port map (
            O => \N__31568\,
            I => \N__31562\
        );

    \I__6836\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31562\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__31562\,
            I => \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DTZ0Z63\
        );

    \I__6834\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31556\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__31556\,
            I => \b2v_inst11.count_off_0_15\
        );

    \I__6832\ : InMux
    port map (
            O => \N__31553\,
            I => \N__31547\
        );

    \I__6831\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31547\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__31544\,
            I => \b2v_inst11.count_off_1_6\
        );

    \I__6828\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31538\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__31538\,
            I => \b2v_inst11.count_off_0_6\
        );

    \I__6826\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31529\
        );

    \I__6825\ : InMux
    port map (
            O => \N__31534\,
            I => \N__31529\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__31526\,
            I => \b2v_inst11.count_off_1_7\
        );

    \I__6822\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31520\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__31520\,
            I => \b2v_inst11.count_off_0_7\
        );

    \I__6820\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31511\
        );

    \I__6819\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31511\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31508\
        );

    \I__6817\ : Odrv4
    port map (
            O => \N__31508\,
            I => \b2v_inst11.count_off_1_8\
        );

    \I__6816\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31502\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__31502\,
            I => \b2v_inst11.count_off_0_8\
        );

    \I__6814\ : CascadeMux
    port map (
            O => \N__31499\,
            I => \b2v_inst6.count_rst_10_cascade_\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__31496\,
            I => \N__31492\
        );

    \I__6812\ : CascadeMux
    port map (
            O => \N__31495\,
            I => \N__31489\
        );

    \I__6811\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31486\
        );

    \I__6810\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31483\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__31486\,
            I => \b2v_inst6.un2_count_1_axb_4\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__31483\,
            I => \b2v_inst6.un2_count_1_axb_4\
        );

    \I__6807\ : InMux
    port map (
            O => \N__31478\,
            I => \b2v_inst11.un3_count_off_1_cry_7\
        );

    \I__6806\ : InMux
    port map (
            O => \N__31475\,
            I => \bfn_11_14_0_\
        );

    \I__6805\ : InMux
    port map (
            O => \N__31472\,
            I => \b2v_inst11.un3_count_off_1_cry_9\
        );

    \I__6804\ : InMux
    port map (
            O => \N__31469\,
            I => \b2v_inst11.un3_count_off_1_cry_10\
        );

    \I__6803\ : InMux
    port map (
            O => \N__31466\,
            I => \b2v_inst11.un3_count_off_1_cry_11\
        );

    \I__6802\ : InMux
    port map (
            O => \N__31463\,
            I => \b2v_inst11.un3_count_off_1_cry_12\
        );

    \I__6801\ : InMux
    port map (
            O => \N__31460\,
            I => \b2v_inst11.un3_count_off_1_cry_13\
        );

    \I__6800\ : InMux
    port map (
            O => \N__31457\,
            I => \b2v_inst11.un3_count_off_1_cry_14\
        );

    \I__6799\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31450\
        );

    \I__6798\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31447\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__31450\,
            I => \N__31444\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__31447\,
            I => \b2v_inst11.count_off_1_14\
        );

    \I__6795\ : Odrv4
    port map (
            O => \N__31444\,
            I => \b2v_inst11.count_off_1_14\
        );

    \I__6794\ : InMux
    port map (
            O => \N__31439\,
            I => \N__31436\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__31436\,
            I => \N__31433\
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__31433\,
            I => \b2v_inst11.count_off_0_14\
        );

    \I__6791\ : CascadeMux
    port map (
            O => \N__31430\,
            I => \b2v_inst11.N_125_cascade_\
        );

    \I__6790\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31424\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__31424\,
            I => \N__31421\
        );

    \I__6788\ : Span4Mux_v
    port map (
            O => \N__31421\,
            I => \N__31417\
        );

    \I__6787\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31414\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__31417\,
            I => \b2v_inst11.N_382_N\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__31414\,
            I => \b2v_inst11.N_382_N\
        );

    \I__6784\ : InMux
    port map (
            O => \N__31409\,
            I => \b2v_inst11.un3_count_off_1_cry_1\
        );

    \I__6783\ : InMux
    port map (
            O => \N__31406\,
            I => \b2v_inst11.un3_count_off_1_cry_2\
        );

    \I__6782\ : InMux
    port map (
            O => \N__31403\,
            I => \b2v_inst11.un3_count_off_1_cry_3\
        );

    \I__6781\ : InMux
    port map (
            O => \N__31400\,
            I => \b2v_inst11.un3_count_off_1_cry_4\
        );

    \I__6780\ : InMux
    port map (
            O => \N__31397\,
            I => \b2v_inst11.un3_count_off_1_cry_5\
        );

    \I__6779\ : InMux
    port map (
            O => \N__31394\,
            I => \b2v_inst11.un3_count_off_1_cry_6\
        );

    \I__6778\ : CascadeMux
    port map (
            O => \N__31391\,
            I => \N__31388\
        );

    \I__6777\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31382\
        );

    \I__6776\ : InMux
    port map (
            O => \N__31387\,
            I => \N__31382\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__31382\,
            I => \b2v_inst11.N_119_f0_1\
        );

    \I__6774\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31370\
        );

    \I__6773\ : CascadeMux
    port map (
            O => \N__31378\,
            I => \N__31366\
        );

    \I__6772\ : CascadeMux
    port map (
            O => \N__31377\,
            I => \N__31361\
        );

    \I__6771\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31358\
        );

    \I__6770\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31351\
        );

    \I__6769\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31351\
        );

    \I__6768\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31351\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31347\
        );

    \I__6766\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31344\
        );

    \I__6765\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31339\
        );

    \I__6764\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31339\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__31364\,
            I => \N__31336\
        );

    \I__6762\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31333\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__31358\,
            I => \N__31327\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__31351\,
            I => \N__31327\
        );

    \I__6759\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31324\
        );

    \I__6758\ : Span4Mux_s1_v
    port map (
            O => \N__31347\,
            I => \N__31319\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__31344\,
            I => \N__31319\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31316\
        );

    \I__6755\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31313\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__31333\,
            I => \N__31306\
        );

    \I__6753\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31303\
        );

    \I__6752\ : Span4Mux_v
    port map (
            O => \N__31327\,
            I => \N__31298\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__31324\,
            I => \N__31298\
        );

    \I__6750\ : Span4Mux_v
    port map (
            O => \N__31319\,
            I => \N__31291\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__31316\,
            I => \N__31291\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__31313\,
            I => \N__31291\
        );

    \I__6747\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31288\
        );

    \I__6746\ : InMux
    port map (
            O => \N__31311\,
            I => \N__31283\
        );

    \I__6745\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31283\
        );

    \I__6744\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31280\
        );

    \I__6743\ : Span4Mux_h
    port map (
            O => \N__31306\,
            I => \N__31277\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__31303\,
            I => \N__31272\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__31298\,
            I => \N__31272\
        );

    \I__6740\ : Span4Mux_h
    port map (
            O => \N__31291\,
            I => \N__31267\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31267\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__31283\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__31280\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__31277\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6735\ : Odrv4
    port map (
            O => \N__31272\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6734\ : Odrv4
    port map (
            O => \N__31267\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6733\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31253\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__31253\,
            I => \b2v_inst11.dutycycle_eena_0\
        );

    \I__6731\ : IoInMux
    port map (
            O => \N__31250\,
            I => \N__31245\
        );

    \I__6730\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31241\
        );

    \I__6729\ : CascadeMux
    port map (
            O => \N__31248\,
            I => \N__31232\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__31245\,
            I => \N__31229\
        );

    \I__6727\ : CascadeMux
    port map (
            O => \N__31244\,
            I => \N__31222\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__31241\,
            I => \N__31218\
        );

    \I__6725\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31215\
        );

    \I__6724\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31212\
        );

    \I__6723\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31200\
        );

    \I__6722\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31200\
        );

    \I__6721\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31200\
        );

    \I__6720\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31200\
        );

    \I__6719\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31197\
        );

    \I__6718\ : IoSpan4Mux
    port map (
            O => \N__31229\,
            I => \N__31186\
        );

    \I__6717\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31177\
        );

    \I__6716\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31177\
        );

    \I__6715\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31177\
        );

    \I__6714\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31177\
        );

    \I__6713\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31172\
        );

    \I__6712\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31172\
        );

    \I__6711\ : Span4Mux_h
    port map (
            O => \N__31218\,
            I => \N__31165\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__31215\,
            I => \N__31165\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__31212\,
            I => \N__31165\
        );

    \I__6708\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31162\
        );

    \I__6707\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31157\
        );

    \I__6706\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31157\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31154\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31148\
        );

    \I__6703\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31145\
        );

    \I__6702\ : InMux
    port map (
            O => \N__31195\,
            I => \N__31140\
        );

    \I__6701\ : InMux
    port map (
            O => \N__31194\,
            I => \N__31140\
        );

    \I__6700\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31135\
        );

    \I__6699\ : InMux
    port map (
            O => \N__31192\,
            I => \N__31135\
        );

    \I__6698\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31128\
        );

    \I__6697\ : InMux
    port map (
            O => \N__31190\,
            I => \N__31128\
        );

    \I__6696\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31128\
        );

    \I__6695\ : Span4Mux_s0_v
    port map (
            O => \N__31186\,
            I => \N__31125\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__31177\,
            I => \N__31119\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__31172\,
            I => \N__31119\
        );

    \I__6692\ : Span4Mux_v
    port map (
            O => \N__31165\,
            I => \N__31114\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__31162\,
            I => \N__31114\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31111\
        );

    \I__6689\ : Span4Mux_v
    port map (
            O => \N__31154\,
            I => \N__31108\
        );

    \I__6688\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31101\
        );

    \I__6687\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31101\
        );

    \I__6686\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31101\
        );

    \I__6685\ : Span4Mux_h
    port map (
            O => \N__31148\,
            I => \N__31088\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__31145\,
            I => \N__31088\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__31140\,
            I => \N__31088\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__31135\,
            I => \N__31088\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31088\
        );

    \I__6680\ : Span4Mux_v
    port map (
            O => \N__31125\,
            I => \N__31088\
        );

    \I__6679\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31085\
        );

    \I__6678\ : Span4Mux_v
    port map (
            O => \N__31119\,
            I => \N__31082\
        );

    \I__6677\ : Span4Mux_v
    port map (
            O => \N__31114\,
            I => \N__31079\
        );

    \I__6676\ : Span4Mux_h
    port map (
            O => \N__31111\,
            I => \N__31070\
        );

    \I__6675\ : Span4Mux_h
    port map (
            O => \N__31108\,
            I => \N__31070\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__31101\,
            I => \N__31070\
        );

    \I__6673\ : Span4Mux_v
    port map (
            O => \N__31088\,
            I => \N__31070\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__31085\,
            I => \G_146\
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__31082\,
            I => \G_146\
        );

    \I__6670\ : Odrv4
    port map (
            O => \N__31079\,
            I => \G_146\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__31070\,
            I => \G_146\
        );

    \I__6668\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31058\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__31058\,
            I => \b2v_inst11.dutycycle_1_0_1\
        );

    \I__6666\ : CascadeMux
    port map (
            O => \N__31055\,
            I => \b2v_inst11.dutycycle_eena_0_cascade_\
        );

    \I__6665\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31046\
        );

    \I__6664\ : InMux
    port map (
            O => \N__31051\,
            I => \N__31046\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__31046\,
            I => \b2v_inst11.dutycycleZ1Z_1\
        );

    \I__6662\ : SRMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__31040\,
            I => \N__31033\
        );

    \I__6660\ : SRMux
    port map (
            O => \N__31039\,
            I => \N__31028\
        );

    \I__6659\ : SRMux
    port map (
            O => \N__31038\,
            I => \N__31025\
        );

    \I__6658\ : SRMux
    port map (
            O => \N__31037\,
            I => \N__31022\
        );

    \I__6657\ : SRMux
    port map (
            O => \N__31036\,
            I => \N__31017\
        );

    \I__6656\ : Span4Mux_h
    port map (
            O => \N__31033\,
            I => \N__31014\
        );

    \I__6655\ : SRMux
    port map (
            O => \N__31032\,
            I => \N__31011\
        );

    \I__6654\ : SRMux
    port map (
            O => \N__31031\,
            I => \N__31008\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__31028\,
            I => \N__31005\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__31025\,
            I => \N__31002\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__31022\,
            I => \N__30999\
        );

    \I__6650\ : SRMux
    port map (
            O => \N__31021\,
            I => \N__30996\
        );

    \I__6649\ : SRMux
    port map (
            O => \N__31020\,
            I => \N__30993\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__30990\
        );

    \I__6647\ : Span4Mux_s2_h
    port map (
            O => \N__31014\,
            I => \N__30985\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__31011\,
            I => \N__30985\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__30981\
        );

    \I__6644\ : Span4Mux_v
    port map (
            O => \N__31005\,
            I => \N__30978\
        );

    \I__6643\ : Span4Mux_v
    port map (
            O => \N__31002\,
            I => \N__30975\
        );

    \I__6642\ : Span4Mux_v
    port map (
            O => \N__30999\,
            I => \N__30970\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30970\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30967\
        );

    \I__6639\ : Span4Mux_v
    port map (
            O => \N__30990\,
            I => \N__30964\
        );

    \I__6638\ : Span4Mux_h
    port map (
            O => \N__30985\,
            I => \N__30961\
        );

    \I__6637\ : SRMux
    port map (
            O => \N__30984\,
            I => \N__30958\
        );

    \I__6636\ : Span4Mux_h
    port map (
            O => \N__30981\,
            I => \N__30955\
        );

    \I__6635\ : Span4Mux_h
    port map (
            O => \N__30978\,
            I => \N__30952\
        );

    \I__6634\ : Span4Mux_h
    port map (
            O => \N__30975\,
            I => \N__30947\
        );

    \I__6633\ : Span4Mux_v
    port map (
            O => \N__30970\,
            I => \N__30947\
        );

    \I__6632\ : Span4Mux_h
    port map (
            O => \N__30967\,
            I => \N__30944\
        );

    \I__6631\ : Span4Mux_s1_h
    port map (
            O => \N__30964\,
            I => \N__30939\
        );

    \I__6630\ : Span4Mux_h
    port map (
            O => \N__30961\,
            I => \N__30939\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__30958\,
            I => \N__30936\
        );

    \I__6628\ : Span4Mux_h
    port map (
            O => \N__30955\,
            I => \N__30931\
        );

    \I__6627\ : Span4Mux_s1_h
    port map (
            O => \N__30952\,
            I => \N__30931\
        );

    \I__6626\ : Span4Mux_h
    port map (
            O => \N__30947\,
            I => \N__30928\
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__30944\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__30939\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__6623\ : Odrv12
    port map (
            O => \N__30936\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__30931\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__30928\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__6620\ : CascadeMux
    port map (
            O => \N__30917\,
            I => \b2v_inst11.count_off_1_0_cascade_\
        );

    \I__6619\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30911\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__30911\,
            I => \N__30908\
        );

    \I__6617\ : Span4Mux_h
    port map (
            O => \N__30908\,
            I => \N__30905\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__30905\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_330_N\
        );

    \I__6615\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30899\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__30899\,
            I => \N__30890\
        );

    \I__6613\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30885\
        );

    \I__6612\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30885\
        );

    \I__6611\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30879\
        );

    \I__6610\ : InMux
    port map (
            O => \N__30895\,
            I => \N__30876\
        );

    \I__6609\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30871\
        );

    \I__6608\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30871\
        );

    \I__6607\ : Span4Mux_v
    port map (
            O => \N__30890\,
            I => \N__30866\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__30885\,
            I => \N__30866\
        );

    \I__6605\ : InMux
    port map (
            O => \N__30884\,
            I => \N__30859\
        );

    \I__6604\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30859\
        );

    \I__6603\ : InMux
    port map (
            O => \N__30882\,
            I => \N__30859\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__30879\,
            I => \b2v_inst11.func_state\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__30876\,
            I => \b2v_inst11.func_state\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__30871\,
            I => \b2v_inst11.func_state\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__30866\,
            I => \b2v_inst11.func_state\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__30859\,
            I => \b2v_inst11.func_state\
        );

    \I__6597\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30845\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__30845\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0\
        );

    \I__6595\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30838\
        );

    \I__6594\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30835\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30832\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__30835\,
            I => \b2v_inst11.N_382\
        );

    \I__6591\ : Odrv12
    port map (
            O => \N__30832\,
            I => \b2v_inst11.N_382\
        );

    \I__6590\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30821\
        );

    \I__6589\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30821\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__30821\,
            I => \N__30817\
        );

    \I__6587\ : InMux
    port map (
            O => \N__30820\,
            I => \N__30814\
        );

    \I__6586\ : Span4Mux_h
    port map (
            O => \N__30817\,
            I => \N__30811\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__30814\,
            I => \N__30808\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__30811\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_1\
        );

    \I__6583\ : Odrv4
    port map (
            O => \N__30808\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_1\
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__30803\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__30800\,
            I => \b2v_inst11.N_315_cascade_\
        );

    \I__6580\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__6578\ : Span4Mux_s3_h
    port map (
            O => \N__30791\,
            I => \N__30788\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__30788\,
            I => \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7\
        );

    \I__6576\ : CascadeMux
    port map (
            O => \N__30785\,
            I => \N__30782\
        );

    \I__6575\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30779\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30774\
        );

    \I__6573\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30769\
        );

    \I__6572\ : InMux
    port map (
            O => \N__30777\,
            I => \N__30769\
        );

    \I__6571\ : Odrv4
    port map (
            O => \N__30774\,
            I => \b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__30769\,
            I => \b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__30764\,
            I => \b2v_inst11.func_state_1_ss0_i_0_o3_0_cascade_\
        );

    \I__6568\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30758\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30754\
        );

    \I__6566\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30751\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__30754\,
            I => \N__30748\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__30751\,
            I => \N__30745\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__30748\,
            I => \N__30742\
        );

    \I__6562\ : Span4Mux_h
    port map (
            O => \N__30745\,
            I => \N__30739\
        );

    \I__6561\ : Odrv4
    port map (
            O => \N__30742\,
            I => \b2v_inst11.N_430\
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__30739\,
            I => \b2v_inst11.N_430\
        );

    \I__6559\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30719\
        );

    \I__6558\ : InMux
    port map (
            O => \N__30733\,
            I => \N__30719\
        );

    \I__6557\ : InMux
    port map (
            O => \N__30732\,
            I => \N__30714\
        );

    \I__6556\ : InMux
    port map (
            O => \N__30731\,
            I => \N__30714\
        );

    \I__6555\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30707\
        );

    \I__6554\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30707\
        );

    \I__6553\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30707\
        );

    \I__6552\ : CascadeMux
    port map (
            O => \N__30727\,
            I => \N__30702\
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__30726\,
            I => \N__30695\
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__30725\,
            I => \N__30685\
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__30724\,
            I => \N__30682\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__30719\,
            I => \N__30673\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__30714\,
            I => \N__30673\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__30707\,
            I => \N__30673\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__30706\,
            I => \N__30670\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__30705\,
            I => \N__30667\
        );

    \I__6543\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30664\
        );

    \I__6542\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30661\
        );

    \I__6541\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30658\
        );

    \I__6540\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30653\
        );

    \I__6539\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30653\
        );

    \I__6538\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30644\
        );

    \I__6537\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30644\
        );

    \I__6536\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30644\
        );

    \I__6535\ : InMux
    port map (
            O => \N__30692\,
            I => \N__30644\
        );

    \I__6534\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30639\
        );

    \I__6533\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30639\
        );

    \I__6532\ : CascadeMux
    port map (
            O => \N__30689\,
            I => \N__30628\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__30688\,
            I => \N__30624\
        );

    \I__6530\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30614\
        );

    \I__6529\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30614\
        );

    \I__6528\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30614\
        );

    \I__6527\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30614\
        );

    \I__6526\ : Span4Mux_v
    port map (
            O => \N__30673\,
            I => \N__30608\
        );

    \I__6525\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30605\
        );

    \I__6524\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30599\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30592\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__30661\,
            I => \N__30583\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__30658\,
            I => \N__30583\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__30653\,
            I => \N__30583\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__30644\,
            I => \N__30583\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30580\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__30638\,
            I => \N__30571\
        );

    \I__6516\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30568\
        );

    \I__6515\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30563\
        );

    \I__6514\ : InMux
    port map (
            O => \N__30635\,
            I => \N__30563\
        );

    \I__6513\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30560\
        );

    \I__6512\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30552\
        );

    \I__6511\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30552\
        );

    \I__6510\ : InMux
    port map (
            O => \N__30631\,
            I => \N__30549\
        );

    \I__6509\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30544\
        );

    \I__6508\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30544\
        );

    \I__6507\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30540\
        );

    \I__6506\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30537\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__30614\,
            I => \N__30534\
        );

    \I__6504\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30527\
        );

    \I__6503\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30527\
        );

    \I__6502\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30527\
        );

    \I__6501\ : Span4Mux_h
    port map (
            O => \N__30608\,
            I => \N__30522\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__30605\,
            I => \N__30522\
        );

    \I__6499\ : InMux
    port map (
            O => \N__30604\,
            I => \N__30519\
        );

    \I__6498\ : InMux
    port map (
            O => \N__30603\,
            I => \N__30516\
        );

    \I__6497\ : CascadeMux
    port map (
            O => \N__30602\,
            I => \N__30511\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__30599\,
            I => \N__30506\
        );

    \I__6495\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30503\
        );

    \I__6494\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30496\
        );

    \I__6493\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30496\
        );

    \I__6492\ : InMux
    port map (
            O => \N__30595\,
            I => \N__30496\
        );

    \I__6491\ : Span4Mux_s3_v
    port map (
            O => \N__30592\,
            I => \N__30489\
        );

    \I__6490\ : Span4Mux_s3_v
    port map (
            O => \N__30583\,
            I => \N__30489\
        );

    \I__6489\ : Span4Mux_s3_v
    port map (
            O => \N__30580\,
            I => \N__30489\
        );

    \I__6488\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30482\
        );

    \I__6487\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30482\
        );

    \I__6486\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30482\
        );

    \I__6485\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30477\
        );

    \I__6484\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30477\
        );

    \I__6483\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30474\
        );

    \I__6482\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30471\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__30568\,
            I => \N__30464\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__30563\,
            I => \N__30464\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__30560\,
            I => \N__30464\
        );

    \I__6478\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30457\
        );

    \I__6477\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30457\
        );

    \I__6476\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30457\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__30552\,
            I => \N__30454\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30451\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__30544\,
            I => \N__30448\
        );

    \I__6472\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30445\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30442\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__30537\,
            I => \N__30429\
        );

    \I__6469\ : Span4Mux_s1_v
    port map (
            O => \N__30534\,
            I => \N__30429\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__30527\,
            I => \N__30429\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__30522\,
            I => \N__30429\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30429\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30429\
        );

    \I__6464\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30424\
        );

    \I__6463\ : InMux
    port map (
            O => \N__30514\,
            I => \N__30424\
        );

    \I__6462\ : InMux
    port map (
            O => \N__30511\,
            I => \N__30421\
        );

    \I__6461\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30415\
        );

    \I__6460\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30415\
        );

    \I__6459\ : Span4Mux_v
    port map (
            O => \N__30506\,
            I => \N__30410\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__30503\,
            I => \N__30410\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30407\
        );

    \I__6456\ : Sp12to4
    port map (
            O => \N__30489\,
            I => \N__30402\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__30482\,
            I => \N__30402\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__30477\,
            I => \N__30399\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30392\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__30471\,
            I => \N__30392\
        );

    \I__6451\ : Sp12to4
    port map (
            O => \N__30464\,
            I => \N__30392\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__30457\,
            I => \N__30388\
        );

    \I__6449\ : Span4Mux_s2_v
    port map (
            O => \N__30454\,
            I => \N__30379\
        );

    \I__6448\ : Span4Mux_v
    port map (
            O => \N__30451\,
            I => \N__30379\
        );

    \I__6447\ : Span4Mux_h
    port map (
            O => \N__30448\,
            I => \N__30379\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__30445\,
            I => \N__30379\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__30442\,
            I => \N__30372\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__30429\,
            I => \N__30372\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30372\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__30421\,
            I => \N__30369\
        );

    \I__6441\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30366\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__30415\,
            I => \N__30361\
        );

    \I__6439\ : Span4Mux_v
    port map (
            O => \N__30410\,
            I => \N__30361\
        );

    \I__6438\ : Span4Mux_s3_h
    port map (
            O => \N__30407\,
            I => \N__30358\
        );

    \I__6437\ : Span12Mux_s7_h
    port map (
            O => \N__30402\,
            I => \N__30351\
        );

    \I__6436\ : Span12Mux_s7_h
    port map (
            O => \N__30399\,
            I => \N__30351\
        );

    \I__6435\ : Span12Mux_s3_v
    port map (
            O => \N__30392\,
            I => \N__30351\
        );

    \I__6434\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30348\
        );

    \I__6433\ : Span4Mux_s2_v
    port map (
            O => \N__30388\,
            I => \N__30337\
        );

    \I__6432\ : Span4Mux_h
    port map (
            O => \N__30379\,
            I => \N__30337\
        );

    \I__6431\ : Span4Mux_v
    port map (
            O => \N__30372\,
            I => \N__30337\
        );

    \I__6430\ : Span4Mux_s3_h
    port map (
            O => \N__30369\,
            I => \N__30337\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__30366\,
            I => \N__30337\
        );

    \I__6428\ : Odrv4
    port map (
            O => \N__30361\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__30358\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__6426\ : Odrv12
    port map (
            O => \N__30351\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__30348\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__6424\ : Odrv4
    port map (
            O => \N__30337\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__30326\,
            I => \N__30321\
        );

    \I__6422\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \N__30318\
        );

    \I__6421\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30315\
        );

    \I__6420\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30310\
        );

    \I__6419\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30310\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__30315\,
            I => \N__30303\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__30310\,
            I => \N__30300\
        );

    \I__6416\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30297\
        );

    \I__6415\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30294\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__30307\,
            I => \N__30291\
        );

    \I__6413\ : CascadeMux
    port map (
            O => \N__30306\,
            I => \N__30287\
        );

    \I__6412\ : Span4Mux_v
    port map (
            O => \N__30303\,
            I => \N__30283\
        );

    \I__6411\ : Span4Mux_s2_h
    port map (
            O => \N__30300\,
            I => \N__30278\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__30297\,
            I => \N__30278\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__30294\,
            I => \N__30272\
        );

    \I__6408\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30265\
        );

    \I__6407\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30265\
        );

    \I__6406\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30265\
        );

    \I__6405\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30262\
        );

    \I__6404\ : Sp12to4
    port map (
            O => \N__30283\,
            I => \N__30259\
        );

    \I__6403\ : Span4Mux_h
    port map (
            O => \N__30278\,
            I => \N__30256\
        );

    \I__6402\ : InMux
    port map (
            O => \N__30277\,
            I => \N__30251\
        );

    \I__6401\ : InMux
    port map (
            O => \N__30276\,
            I => \N__30251\
        );

    \I__6400\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30248\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__30272\,
            I => \N__30241\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__30265\,
            I => \N__30241\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__30262\,
            I => \N__30241\
        );

    \I__6396\ : Odrv12
    port map (
            O => \N__30259\,
            I => \b2v_inst11.N_161\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__30256\,
            I => \b2v_inst11.N_161\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__30251\,
            I => \b2v_inst11.N_161\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__30248\,
            I => \b2v_inst11.N_161\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__30241\,
            I => \b2v_inst11.N_161\
        );

    \I__6391\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30227\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__30227\,
            I => \b2v_inst11.N_339\
        );

    \I__6389\ : InMux
    port map (
            O => \N__30224\,
            I => \N__30221\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__30221\,
            I => \N__30218\
        );

    \I__6387\ : Span4Mux_s2_h
    port map (
            O => \N__30218\,
            I => \N__30215\
        );

    \I__6386\ : Span4Mux_v
    port map (
            O => \N__30215\,
            I => \N__30212\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__30212\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__30209\,
            I => \b2v_inst11.dutycycle_1_0_1_cascade_\
        );

    \I__6383\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30203\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__30203\,
            I => \b2v_inst11.dutycycle_eena\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__30200\,
            I => \N__30197\
        );

    \I__6380\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30191\
        );

    \I__6379\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30191\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__30191\,
            I => \b2v_inst11.dutycycleZ1Z_0\
        );

    \I__6377\ : CascadeMux
    port map (
            O => \N__30188\,
            I => \b2v_inst11.dutycycle_eena_cascade_\
        );

    \I__6376\ : CascadeMux
    port map (
            O => \N__30185\,
            I => \N__30180\
        );

    \I__6375\ : CascadeMux
    port map (
            O => \N__30184\,
            I => \N__30177\
        );

    \I__6374\ : InMux
    port map (
            O => \N__30183\,
            I => \N__30172\
        );

    \I__6373\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30169\
        );

    \I__6372\ : InMux
    port map (
            O => \N__30177\,
            I => \N__30161\
        );

    \I__6371\ : InMux
    port map (
            O => \N__30176\,
            I => \N__30161\
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__30175\,
            I => \N__30158\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30155\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30151\
        );

    \I__6367\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30148\
        );

    \I__6366\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30145\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__30166\,
            I => \N__30139\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__30161\,
            I => \N__30136\
        );

    \I__6363\ : InMux
    port map (
            O => \N__30158\,
            I => \N__30133\
        );

    \I__6362\ : Span4Mux_s1_v
    port map (
            O => \N__30155\,
            I => \N__30130\
        );

    \I__6361\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30127\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__30151\,
            I => \N__30119\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__30148\,
            I => \N__30119\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__30145\,
            I => \N__30119\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__30144\,
            I => \N__30116\
        );

    \I__6356\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30112\
        );

    \I__6355\ : InMux
    port map (
            O => \N__30142\,
            I => \N__30107\
        );

    \I__6354\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30107\
        );

    \I__6353\ : Span4Mux_v
    port map (
            O => \N__30136\,
            I => \N__30102\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__30133\,
            I => \N__30102\
        );

    \I__6351\ : Span4Mux_h
    port map (
            O => \N__30130\,
            I => \N__30097\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30097\
        );

    \I__6349\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30094\
        );

    \I__6348\ : Span4Mux_v
    port map (
            O => \N__30119\,
            I => \N__30091\
        );

    \I__6347\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30088\
        );

    \I__6346\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30085\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30078\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30078\
        );

    \I__6343\ : Span4Mux_h
    port map (
            O => \N__30102\,
            I => \N__30078\
        );

    \I__6342\ : Span4Mux_v
    port map (
            O => \N__30097\,
            I => \N__30073\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__30094\,
            I => \N__30073\
        );

    \I__6340\ : Span4Mux_h
    port map (
            O => \N__30091\,
            I => \N__30068\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__30088\,
            I => \N__30068\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__30085\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__30078\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__6336\ : Odrv4
    port map (
            O => \N__30073\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__6335\ : Odrv4
    port map (
            O => \N__30068\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__30059\,
            I => \b2v_inst11.dutycycleZ0Z_0_cascade_\
        );

    \I__6333\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30050\
        );

    \I__6332\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30050\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__30050\,
            I => \b2v_inst11.dutycycle_1_0_0\
        );

    \I__6330\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__30044\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__30041\,
            I => \b2v_inst11.dutycycleZ0Z_2_cascade_\
        );

    \I__6327\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__30035\,
            I => \N__30032\
        );

    \I__6325\ : Span4Mux_h
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__6324\ : Span4Mux_h
    port map (
            O => \N__30029\,
            I => \N__30026\
        );

    \I__6323\ : Span4Mux_v
    port map (
            O => \N__30026\,
            I => \N__30023\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__30023\,
            I => \b2v_inst11.mult1_un152_sum_i\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__30020\,
            I => \N__30016\
        );

    \I__6320\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30011\
        );

    \I__6319\ : InMux
    port map (
            O => \N__30016\,
            I => \N__30011\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__30011\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_0_2\
        );

    \I__6317\ : InMux
    port map (
            O => \N__30008\,
            I => \N__30002\
        );

    \I__6316\ : InMux
    port map (
            O => \N__30007\,
            I => \N__30002\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__6314\ : Odrv4
    port map (
            O => \N__29999\,
            I => \b2v_inst11.N_168\
        );

    \I__6313\ : InMux
    port map (
            O => \N__29996\,
            I => \N__29990\
        );

    \I__6312\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29990\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29987\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__29987\,
            I => \b2v_inst11.dutycycle_RNIAEUL3Z0Z_2\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__6308\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29975\
        );

    \I__6307\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29975\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__29975\,
            I => \b2v_inst11.dutycycleZ1Z_2\
        );

    \I__6305\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29958\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__29971\,
            I => \N__29954\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29948\
        );

    \I__6302\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29948\
        );

    \I__6301\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29943\
        );

    \I__6300\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29943\
        );

    \I__6299\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29938\
        );

    \I__6298\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29935\
        );

    \I__6297\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29932\
        );

    \I__6296\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29927\
        );

    \I__6295\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29927\
        );

    \I__6294\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29923\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29920\
        );

    \I__6292\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29917\
        );

    \I__6291\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29912\
        );

    \I__6290\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29912\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__29948\,
            I => \N__29907\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29907\
        );

    \I__6287\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29903\
        );

    \I__6286\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29900\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__29938\,
            I => \N__29897\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__29935\,
            I => \N__29892\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__29932\,
            I => \N__29892\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__29927\,
            I => \N__29887\
        );

    \I__6281\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29883\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__29923\,
            I => \N__29878\
        );

    \I__6279\ : Span4Mux_v
    port map (
            O => \N__29920\,
            I => \N__29878\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29917\,
            I => \N__29871\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__29912\,
            I => \N__29871\
        );

    \I__6276\ : Span4Mux_h
    port map (
            O => \N__29907\,
            I => \N__29871\
        );

    \I__6275\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29868\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__29903\,
            I => \N__29865\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__29900\,
            I => \N__29858\
        );

    \I__6272\ : Span4Mux_v
    port map (
            O => \N__29897\,
            I => \N__29858\
        );

    \I__6271\ : Span4Mux_h
    port map (
            O => \N__29892\,
            I => \N__29858\
        );

    \I__6270\ : InMux
    port map (
            O => \N__29891\,
            I => \N__29855\
        );

    \I__6269\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29852\
        );

    \I__6268\ : Span4Mux_v
    port map (
            O => \N__29887\,
            I => \N__29849\
        );

    \I__6267\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29846\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29841\
        );

    \I__6265\ : Span4Mux_h
    port map (
            O => \N__29878\,
            I => \N__29841\
        );

    \I__6264\ : Span4Mux_v
    port map (
            O => \N__29871\,
            I => \N__29838\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__29868\,
            I => \N__29835\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__29865\,
            I => \N__29826\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__29858\,
            I => \N__29826\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29826\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29826\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__29849\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__29846\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__29841\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__29838\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__6254\ : Odrv12
    port map (
            O => \N__29835\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__29826\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__6252\ : CascadeMux
    port map (
            O => \N__29813\,
            I => \N__29810\
        );

    \I__6251\ : InMux
    port map (
            O => \N__29810\,
            I => \N__29804\
        );

    \I__6250\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29804\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__29804\,
            I => \N__29801\
        );

    \I__6248\ : Span4Mux_v
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__6247\ : Sp12to4
    port map (
            O => \N__29798\,
            I => \N__29794\
        );

    \I__6246\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29791\
        );

    \I__6245\ : Odrv12
    port map (
            O => \N__29794\,
            I => \b2v_inst11.N_365\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__29791\,
            I => \b2v_inst11.N_365\
        );

    \I__6243\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29783\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__29783\,
            I => \N__29780\
        );

    \I__6241\ : Span4Mux_v
    port map (
            O => \N__29780\,
            I => \N__29777\
        );

    \I__6240\ : Span4Mux_h
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__6239\ : Odrv4
    port map (
            O => \N__29774\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1\
        );

    \I__6238\ : CascadeMux
    port map (
            O => \N__29771\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_\
        );

    \I__6237\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29765\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__29765\,
            I => \N__29762\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__29762\,
            I => \N__29759\
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__29759\,
            I => \b2v_inst11.N_186_i\
        );

    \I__6233\ : InMux
    port map (
            O => \N__29756\,
            I => \N__29750\
        );

    \I__6232\ : InMux
    port map (
            O => \N__29755\,
            I => \N__29743\
        );

    \I__6231\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29743\
        );

    \I__6230\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29743\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__29750\,
            I => \N__29738\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__29743\,
            I => \N__29738\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__29738\,
            I => \N__29735\
        );

    \I__6226\ : Span4Mux_h
    port map (
            O => \N__29735\,
            I => \N__29732\
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__29732\,
            I => \b2v_inst6.N_192\
        );

    \I__6224\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29726\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29722\
        );

    \I__6222\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29719\
        );

    \I__6221\ : Odrv12
    port map (
            O => \N__29722\,
            I => \N_241\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__29719\,
            I => \N_241\
        );

    \I__6219\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29708\
        );

    \I__6218\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29708\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__29708\,
            I => \b2v_inst6.N_276_0\
        );

    \I__6216\ : CascadeMux
    port map (
            O => \N__29705\,
            I => \N__29701\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__6214\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29694\
        );

    \I__6213\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29691\
        );

    \I__6212\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29688\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__29694\,
            I => \b2v_inst6.curr_state_RNIUP4B1Z0Z_0\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__29691\,
            I => \b2v_inst6.curr_state_RNIUP4B1Z0Z_0\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__29688\,
            I => \b2v_inst6.curr_state_RNIUP4B1Z0Z_0\
        );

    \I__6208\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29675\
        );

    \I__6207\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29675\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__29675\,
            I => \b2v_inst6.delayed_vccin_vccinaux_ok_0\
        );

    \I__6205\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29669\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__29669\,
            I => \N__29666\
        );

    \I__6203\ : Span4Mux_v
    port map (
            O => \N__29666\,
            I => \N__29663\
        );

    \I__6202\ : Span4Mux_h
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__6201\ : Odrv4
    port map (
            O => \N__29660\,
            I => \b2v_inst11.N_9\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__29657\,
            I => \b2v_inst11.N_172_cascade_\
        );

    \I__6199\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29651\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__29651\,
            I => \N__29648\
        );

    \I__6197\ : Span4Mux_v
    port map (
            O => \N__29648\,
            I => \N__29645\
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__29645\,
            I => \b2v_inst11.g0_i_a7_1_3\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__29642\,
            I => \b2v_inst11.g0_i_0_cascade_\
        );

    \I__6194\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29631\
        );

    \I__6193\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29631\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__29637\,
            I => \N__29628\
        );

    \I__6191\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29625\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__29631\,
            I => \N__29620\
        );

    \I__6189\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29617\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__29625\,
            I => \N__29614\
        );

    \I__6187\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29609\
        );

    \I__6186\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29609\
        );

    \I__6185\ : Sp12to4
    port map (
            O => \N__29620\,
            I => \N__29602\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__29617\,
            I => \N__29602\
        );

    \I__6183\ : Span4Mux_s3_h
    port map (
            O => \N__29614\,
            I => \N__29597\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__29609\,
            I => \N__29597\
        );

    \I__6181\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29592\
        );

    \I__6180\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29592\
        );

    \I__6179\ : Odrv12
    port map (
            O => \N__29602\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__29597\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__29592\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__6176\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__29579\,
            I => \N__29576\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__29576\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__29573\,
            I => \b2v_inst11.N_295_cascade_\
        );

    \I__6171\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__29567\,
            I => \N__29564\
        );

    \I__6169\ : Odrv12
    port map (
            O => \N__29564\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3_out\
        );

    \I__6168\ : InMux
    port map (
            O => \N__29561\,
            I => \N__29558\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__29558\,
            I => \N__29555\
        );

    \I__6166\ : Span4Mux_v
    port map (
            O => \N__29555\,
            I => \N__29552\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__6164\ : Odrv4
    port map (
            O => \N__29549\,
            I => \b2v_inst11.N_355\
        );

    \I__6163\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29543\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__29543\,
            I => \b2v_inst6.curr_state_1_1\
        );

    \I__6161\ : CascadeMux
    port map (
            O => \N__29540\,
            I => \b2v_inst6.N_42_cascade_\
        );

    \I__6160\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29530\
        );

    \I__6159\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29530\
        );

    \I__6158\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29527\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__29530\,
            I => \b2v_inst6.curr_stateZ0Z_1\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__29527\,
            I => \b2v_inst6.curr_stateZ0Z_1\
        );

    \I__6155\ : CascadeMux
    port map (
            O => \N__29522\,
            I => \b2v_inst6.curr_stateZ0Z_1_cascade_\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__29519\,
            I => \b2v_inst6.N_3053_i_cascade_\
        );

    \I__6153\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29511\
        );

    \I__6152\ : InMux
    port map (
            O => \N__29515\,
            I => \N__29506\
        );

    \I__6151\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29506\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__29511\,
            I => \b2v_inst6.N_3034_i\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__29506\,
            I => \b2v_inst6.N_3034_i\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__29501\,
            I => \b2v_inst6.N_3034_i_cascade_\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__29498\,
            I => \b2v_inst6.curr_state_RNIUP4B1Z0Z_0_cascade_\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__29495\,
            I => \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\
        );

    \I__6145\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29484\
        );

    \I__6144\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29477\
        );

    \I__6143\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29477\
        );

    \I__6142\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29477\
        );

    \I__6141\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29472\
        );

    \I__6140\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29472\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29465\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__29477\,
            I => \N__29465\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__29472\,
            I => \N__29465\
        );

    \I__6136\ : Span4Mux_s2_v
    port map (
            O => \N__29465\,
            I => \N__29462\
        );

    \I__6135\ : Span4Mux_v
    port map (
            O => \N__29462\,
            I => \N__29459\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__6133\ : Odrv4
    port map (
            O => \N__29456\,
            I => \N_222\
        );

    \I__6132\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29444\
        );

    \I__6131\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29444\
        );

    \I__6130\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29444\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__29444\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__29441\,
            I => \N__29437\
        );

    \I__6127\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29429\
        );

    \I__6126\ : InMux
    port map (
            O => \N__29437\,
            I => \N__29429\
        );

    \I__6125\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29429\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__29429\,
            I => \b2v_inst6.N_3053_i\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__29426\,
            I => \N__29422\
        );

    \I__6122\ : InMux
    port map (
            O => \N__29425\,
            I => \N__29419\
        );

    \I__6121\ : InMux
    port map (
            O => \N__29422\,
            I => \N__29416\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__29419\,
            I => \N__29413\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__29416\,
            I => \b2v_inst6.un2_count_1_axb_9\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__29413\,
            I => \b2v_inst6.un2_count_1_axb_9\
        );

    \I__6117\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29402\
        );

    \I__6116\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29402\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__29402\,
            I => \N__29399\
        );

    \I__6114\ : Odrv12
    port map (
            O => \N__29399\,
            I => \b2v_inst6.un2_count_1_cry_8_THRU_CO\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__29396\,
            I => \b2v_inst6.un2_count_1_axb_9_cascade_\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__29393\,
            I => \b2v_inst6.count_rst_6_cascade_\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__29390\,
            I => \N__29386\
        );

    \I__6110\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29381\
        );

    \I__6109\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29381\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__29381\,
            I => \N__29378\
        );

    \I__6107\ : Odrv12
    port map (
            O => \N__29378\,
            I => \b2v_inst6.un2_count_1_cry_7_THRU_CO\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__29375\,
            I => \b2v_inst6.countZ0Z_8_cascade_\
        );

    \I__6105\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29369\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__29369\,
            I => \N__29366\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__29366\,
            I => \b2v_inst6.count_0_8\
        );

    \I__6102\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29360\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__29360\,
            I => \b2v_inst6.curr_state_1_0\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__29357\,
            I => \b2v_inst6.curr_state_7_0_cascade_\
        );

    \I__6099\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29351\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__29351\,
            I => \b2v_inst6.N_42\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__29348\,
            I => \b2v_inst6.countZ0Z_6_cascade_\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__29345\,
            I => \b2v_inst6.count_1_i_a3_0_0_cascade_\
        );

    \I__6095\ : InMux
    port map (
            O => \N__29342\,
            I => \N__29338\
        );

    \I__6094\ : InMux
    port map (
            O => \N__29341\,
            I => \N__29335\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__29338\,
            I => \N__29330\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__29335\,
            I => \N__29327\
        );

    \I__6091\ : CascadeMux
    port map (
            O => \N__29334\,
            I => \N__29322\
        );

    \I__6090\ : CascadeMux
    port map (
            O => \N__29333\,
            I => \N__29319\
        );

    \I__6089\ : Sp12to4
    port map (
            O => \N__29330\,
            I => \N__29315\
        );

    \I__6088\ : Span4Mux_s2_h
    port map (
            O => \N__29327\,
            I => \N__29312\
        );

    \I__6087\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29301\
        );

    \I__6086\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29301\
        );

    \I__6085\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29301\
        );

    \I__6084\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29301\
        );

    \I__6083\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29301\
        );

    \I__6082\ : Odrv12
    port map (
            O => \N__29315\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__6081\ : Odrv4
    port map (
            O => \N__29312\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__29301\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__6079\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29289\
        );

    \I__6078\ : CascadeMux
    port map (
            O => \N__29293\,
            I => \N__29286\
        );

    \I__6077\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29279\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__29289\,
            I => \N__29276\
        );

    \I__6075\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29273\
        );

    \I__6074\ : InMux
    port map (
            O => \N__29285\,
            I => \N__29264\
        );

    \I__6073\ : InMux
    port map (
            O => \N__29284\,
            I => \N__29264\
        );

    \I__6072\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29264\
        );

    \I__6071\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29264\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29261\
        );

    \I__6069\ : Span4Mux_v
    port map (
            O => \N__29276\,
            I => \N__29252\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__29273\,
            I => \N__29252\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__29264\,
            I => \N__29252\
        );

    \I__6066\ : Span4Mux_v
    port map (
            O => \N__29261\,
            I => \N__29252\
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__29252\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__6064\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29239\
        );

    \I__6063\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29228\
        );

    \I__6062\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29228\
        );

    \I__6061\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29228\
        );

    \I__6060\ : InMux
    port map (
            O => \N__29245\,
            I => \N__29228\
        );

    \I__6059\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29228\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__29243\,
            I => \N__29225\
        );

    \I__6057\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29222\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__29239\,
            I => \N__29217\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__29228\,
            I => \N__29217\
        );

    \I__6054\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29214\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__29222\,
            I => \N__29211\
        );

    \I__6052\ : Span4Mux_h
    port map (
            O => \N__29217\,
            I => \N__29206\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29206\
        );

    \I__6050\ : Span4Mux_h
    port map (
            O => \N__29211\,
            I => \N__29203\
        );

    \I__6049\ : Sp12to4
    port map (
            O => \N__29206\,
            I => \N__29198\
        );

    \I__6048\ : Sp12to4
    port map (
            O => \N__29203\,
            I => \N__29198\
        );

    \I__6047\ : Span12Mux_v
    port map (
            O => \N__29198\,
            I => \N__29195\
        );

    \I__6046\ : Odrv12
    port map (
            O => \N__29195\,
            I => v33dsw_ok
        );

    \I__6045\ : CascadeMux
    port map (
            O => \N__29192\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_\
        );

    \I__6044\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29185\
        );

    \I__6043\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29182\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29179\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__29182\,
            I => \N__29176\
        );

    \I__6040\ : Span4Mux_h
    port map (
            O => \N__29179\,
            I => \N__29173\
        );

    \I__6039\ : Odrv12
    port map (
            O => \N__29176\,
            I => \b2v_inst36.countZ0Z_9\
        );

    \I__6038\ : Odrv4
    port map (
            O => \N__29173\,
            I => \b2v_inst36.countZ0Z_9\
        );

    \I__6037\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29162\
        );

    \I__6036\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29162\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__29162\,
            I => \N__29159\
        );

    \I__6034\ : Odrv4
    port map (
            O => \N__29159\,
            I => \b2v_inst36.count_rst_5\
        );

    \I__6033\ : InMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__29153\,
            I => \b2v_inst36.count_2_9\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__29150\,
            I => \N__29142\
        );

    \I__6030\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29136\
        );

    \I__6029\ : CEMux
    port map (
            O => \N__29148\,
            I => \N__29136\
        );

    \I__6028\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29127\
        );

    \I__6027\ : CEMux
    port map (
            O => \N__29146\,
            I => \N__29127\
        );

    \I__6026\ : CEMux
    port map (
            O => \N__29145\,
            I => \N__29123\
        );

    \I__6025\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29111\
        );

    \I__6024\ : CEMux
    port map (
            O => \N__29141\,
            I => \N__29111\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29103\
        );

    \I__6022\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29098\
        );

    \I__6021\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29098\
        );

    \I__6020\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29088\
        );

    \I__6019\ : CEMux
    port map (
            O => \N__29132\,
            I => \N__29088\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__29127\,
            I => \N__29085\
        );

    \I__6017\ : CEMux
    port map (
            O => \N__29126\,
            I => \N__29082\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__29123\,
            I => \N__29079\
        );

    \I__6015\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29070\
        );

    \I__6014\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29070\
        );

    \I__6013\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29070\
        );

    \I__6012\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29070\
        );

    \I__6011\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29063\
        );

    \I__6010\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29063\
        );

    \I__6009\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29063\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__29111\,
            I => \N__29060\
        );

    \I__6007\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29053\
        );

    \I__6006\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29053\
        );

    \I__6005\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29053\
        );

    \I__6004\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29048\
        );

    \I__6003\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29048\
        );

    \I__6002\ : Span4Mux_h
    port map (
            O => \N__29103\,
            I => \N__29043\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29043\
        );

    \I__6000\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29032\
        );

    \I__5999\ : CEMux
    port map (
            O => \N__29096\,
            I => \N__29032\
        );

    \I__5998\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29032\
        );

    \I__5997\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29032\
        );

    \I__5996\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29032\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__29088\,
            I => \N__29029\
        );

    \I__5994\ : Span4Mux_h
    port map (
            O => \N__29085\,
            I => \N__29024\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__29082\,
            I => \N__29024\
        );

    \I__5992\ : Span4Mux_s3_v
    port map (
            O => \N__29079\,
            I => \N__29021\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__29070\,
            I => \N__29016\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29016\
        );

    \I__5989\ : Span4Mux_s1_v
    port map (
            O => \N__29060\,
            I => \N__29005\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__29053\,
            I => \N__29005\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__29048\,
            I => \N__29005\
        );

    \I__5986\ : Span4Mux_s1_v
    port map (
            O => \N__29043\,
            I => \N__29005\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__29032\,
            I => \N__29005\
        );

    \I__5984\ : Span4Mux_h
    port map (
            O => \N__29029\,
            I => \N__29002\
        );

    \I__5983\ : Sp12to4
    port map (
            O => \N__29024\,
            I => \N__28999\
        );

    \I__5982\ : Span4Mux_v
    port map (
            O => \N__29021\,
            I => \N__28994\
        );

    \I__5981\ : Span4Mux_s3_v
    port map (
            O => \N__29016\,
            I => \N__28994\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__29005\,
            I => \N__28991\
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__29002\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__5978\ : Odrv12
    port map (
            O => \N__28999\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__28994\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__28991\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__5975\ : SRMux
    port map (
            O => \N__28982\,
            I => \N__28977\
        );

    \I__5974\ : SRMux
    port map (
            O => \N__28981\,
            I => \N__28969\
        );

    \I__5973\ : SRMux
    port map (
            O => \N__28980\,
            I => \N__28966\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__28977\,
            I => \N__28956\
        );

    \I__5971\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28951\
        );

    \I__5970\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28951\
        );

    \I__5969\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28946\
        );

    \I__5968\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28946\
        );

    \I__5967\ : SRMux
    port map (
            O => \N__28972\,
            I => \N__28942\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__28969\,
            I => \N__28931\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__28966\,
            I => \N__28928\
        );

    \I__5964\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28921\
        );

    \I__5963\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28921\
        );

    \I__5962\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28921\
        );

    \I__5961\ : SRMux
    port map (
            O => \N__28962\,
            I => \N__28911\
        );

    \I__5960\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28904\
        );

    \I__5959\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28904\
        );

    \I__5958\ : SRMux
    port map (
            O => \N__28959\,
            I => \N__28904\
        );

    \I__5957\ : Span4Mux_s2_v
    port map (
            O => \N__28956\,
            I => \N__28899\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28899\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__28946\,
            I => \N__28896\
        );

    \I__5954\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28893\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28890\
        );

    \I__5952\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28883\
        );

    \I__5951\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28883\
        );

    \I__5950\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28883\
        );

    \I__5949\ : SRMux
    port map (
            O => \N__28938\,
            I => \N__28878\
        );

    \I__5948\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28878\
        );

    \I__5947\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28871\
        );

    \I__5946\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28871\
        );

    \I__5945\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28871\
        );

    \I__5944\ : Span4Mux_h
    port map (
            O => \N__28931\,
            I => \N__28866\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__28928\,
            I => \N__28866\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__28921\,
            I => \N__28863\
        );

    \I__5941\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28856\
        );

    \I__5940\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28856\
        );

    \I__5939\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28856\
        );

    \I__5938\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28853\
        );

    \I__5937\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28850\
        );

    \I__5936\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28845\
        );

    \I__5935\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28845\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28834\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__28904\,
            I => \N__28834\
        );

    \I__5932\ : Span4Mux_v
    port map (
            O => \N__28899\,
            I => \N__28834\
        );

    \I__5931\ : Span4Mux_h
    port map (
            O => \N__28896\,
            I => \N__28834\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__28893\,
            I => \N__28834\
        );

    \I__5929\ : Span4Mux_v
    port map (
            O => \N__28890\,
            I => \N__28827\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__28883\,
            I => \N__28827\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__28878\,
            I => \N__28827\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__28871\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__28866\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5924\ : Odrv4
    port map (
            O => \N__28863\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__28856\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__28853\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__28850\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__28845\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5919\ : Odrv4
    port map (
            O => \N__28834\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__28827\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__5917\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28802\
        );

    \I__5916\ : InMux
    port map (
            O => \N__28807\,
            I => \N__28802\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__28799\,
            I => \b2v_inst6.count_0_10\
        );

    \I__5913\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28791\
        );

    \I__5912\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28788\
        );

    \I__5911\ : InMux
    port map (
            O => \N__28794\,
            I => \N__28785\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__28791\,
            I => \N__28780\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__28788\,
            I => \N__28780\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__28785\,
            I => \b2v_inst6.count_rst_4\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__28780\,
            I => \b2v_inst6.count_rst_4\
        );

    \I__5906\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28772\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__28772\,
            I => \N__28769\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__28769\,
            I => \b2v_inst6.un2_count_1_axb_10\
        );

    \I__5903\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28763\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__28763\,
            I => \N__28760\
        );

    \I__5901\ : Sp12to4
    port map (
            O => \N__28760\,
            I => \N__28757\
        );

    \I__5900\ : Span12Mux_v
    port map (
            O => \N__28757\,
            I => \N__28754\
        );

    \I__5899\ : Odrv12
    port map (
            O => \N__28754\,
            I => v33a_ok
        );

    \I__5898\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__28748\,
            I => \N__28745\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__28745\,
            I => \N__28742\
        );

    \I__5895\ : Odrv4
    port map (
            O => \N__28742\,
            I => vccst_cpu_ok
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__28739\,
            I => \N__28736\
        );

    \I__5893\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28733\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__28733\,
            I => \N__28730\
        );

    \I__5891\ : Span4Mux_v
    port map (
            O => \N__28730\,
            I => \N__28727\
        );

    \I__5890\ : Span4Mux_v
    port map (
            O => \N__28727\,
            I => \N__28724\
        );

    \I__5889\ : Sp12to4
    port map (
            O => \N__28724\,
            I => \N__28721\
        );

    \I__5888\ : Odrv12
    port map (
            O => \N__28721\,
            I => v1p8a_ok
        );

    \I__5887\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28715\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__28715\,
            I => \N__28712\
        );

    \I__5885\ : Odrv12
    port map (
            O => \N__28712\,
            I => v5a_ok
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__28709\,
            I => \b2v_inst6.count_rst_5_cascade_\
        );

    \I__5883\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28703\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__28703\,
            I => \b2v_inst6.count_0_15\
        );

    \I__5881\ : InMux
    port map (
            O => \N__28700\,
            I => \N__28694\
        );

    \I__5880\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28694\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__28694\,
            I => \b2v_inst6.count_rst\
        );

    \I__5878\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28688\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__28688\,
            I => \b2v_inst6.countZ0Z_15\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__28685\,
            I => \b2v_inst6.countZ0Z_15_cascade_\
        );

    \I__5875\ : InMux
    port map (
            O => \N__28682\,
            I => \N__28678\
        );

    \I__5874\ : InMux
    port map (
            O => \N__28681\,
            I => \N__28675\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__28678\,
            I => \N__28672\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__28675\,
            I => \b2v_inst6.un2_count_1_axb_7\
        );

    \I__5871\ : Odrv4
    port map (
            O => \N__28672\,
            I => \b2v_inst6.un2_count_1_axb_7\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__28667\,
            I => \N__28664\
        );

    \I__5869\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28658\
        );

    \I__5868\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28658\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28655\
        );

    \I__5866\ : Odrv12
    port map (
            O => \N__28655\,
            I => \b2v_inst6.un2_count_1_cry_6_THRU_CO\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__28652\,
            I => \b2v_inst6.un2_count_1_axb_7_cascade_\
        );

    \I__5864\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28646\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__28646\,
            I => \b2v_inst6.count_rst_7\
        );

    \I__5862\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28637\
        );

    \I__5861\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28637\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__28637\,
            I => \b2v_inst6.count_0_7\
        );

    \I__5859\ : CascadeMux
    port map (
            O => \N__28634\,
            I => \b2v_inst6.count_rst_7_cascade_\
        );

    \I__5858\ : CascadeMux
    port map (
            O => \N__28631\,
            I => \b2v_inst6.count_en_cascade_\
        );

    \I__5857\ : InMux
    port map (
            O => \N__28628\,
            I => \N__28625\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__28625\,
            I => \N__28622\
        );

    \I__5855\ : Odrv4
    port map (
            O => \N__28622\,
            I => \b2v_inst6.countZ0Z_6\
        );

    \I__5854\ : InMux
    port map (
            O => \N__28619\,
            I => \bfn_11_2_0_\
        );

    \I__5853\ : InMux
    port map (
            O => \N__28616\,
            I => \b2v_inst6.un2_count_1_cry_9\
        );

    \I__5852\ : InMux
    port map (
            O => \N__28613\,
            I => \b2v_inst6.un2_count_1_cry_10\
        );

    \I__5851\ : InMux
    port map (
            O => \N__28610\,
            I => \b2v_inst6.un2_count_1_cry_11\
        );

    \I__5850\ : InMux
    port map (
            O => \N__28607\,
            I => \b2v_inst6.un2_count_1_cry_12\
        );

    \I__5849\ : InMux
    port map (
            O => \N__28604\,
            I => \b2v_inst6.un2_count_1_cry_13\
        );

    \I__5848\ : InMux
    port map (
            O => \N__28601\,
            I => \b2v_inst6.un2_count_1_cry_14\
        );

    \I__5847\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28592\
        );

    \I__5846\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28592\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__28592\,
            I => \b2v_inst11.count_clk_1_13\
        );

    \I__5844\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__28586\,
            I => \b2v_inst11.count_clk_0_13\
        );

    \I__5842\ : CEMux
    port map (
            O => \N__28583\,
            I => \N__28579\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__28582\,
            I => \N__28576\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__28579\,
            I => \N__28573\
        );

    \I__5839\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28565\
        );

    \I__5838\ : Span4Mux_s3_v
    port map (
            O => \N__28573\,
            I => \N__28562\
        );

    \I__5837\ : CEMux
    port map (
            O => \N__28572\,
            I => \N__28559\
        );

    \I__5836\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28551\
        );

    \I__5835\ : CEMux
    port map (
            O => \N__28570\,
            I => \N__28548\
        );

    \I__5834\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28543\
        );

    \I__5833\ : CEMux
    port map (
            O => \N__28568\,
            I => \N__28543\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__28565\,
            I => \N__28531\
        );

    \I__5831\ : Span4Mux_h
    port map (
            O => \N__28562\,
            I => \N__28531\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__28559\,
            I => \N__28531\
        );

    \I__5829\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28522\
        );

    \I__5828\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28522\
        );

    \I__5827\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28522\
        );

    \I__5826\ : CEMux
    port map (
            O => \N__28555\,
            I => \N__28522\
        );

    \I__5825\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28519\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28516\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__28548\,
            I => \N__28513\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__28543\,
            I => \N__28510\
        );

    \I__5821\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28501\
        );

    \I__5820\ : CEMux
    port map (
            O => \N__28541\,
            I => \N__28501\
        );

    \I__5819\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28501\
        );

    \I__5818\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28501\
        );

    \I__5817\ : CEMux
    port map (
            O => \N__28538\,
            I => \N__28498\
        );

    \I__5816\ : IoSpan4Mux
    port map (
            O => \N__28531\,
            I => \N__28493\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28493\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__28519\,
            I => \N__28490\
        );

    \I__5813\ : Span4Mux_s2_v
    port map (
            O => \N__28516\,
            I => \N__28480\
        );

    \I__5812\ : Span4Mux_h
    port map (
            O => \N__28513\,
            I => \N__28480\
        );

    \I__5811\ : Span4Mux_s1_v
    port map (
            O => \N__28510\,
            I => \N__28475\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__28501\,
            I => \N__28475\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__28498\,
            I => \N__28468\
        );

    \I__5808\ : Span4Mux_s1_v
    port map (
            O => \N__28493\,
            I => \N__28468\
        );

    \I__5807\ : Span4Mux_s1_v
    port map (
            O => \N__28490\,
            I => \N__28468\
        );

    \I__5806\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28465\
        );

    \I__5805\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28456\
        );

    \I__5804\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28456\
        );

    \I__5803\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28456\
        );

    \I__5802\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28456\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__28480\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__28475\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__28468\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__28465\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__28456\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__5796\ : InMux
    port map (
            O => \N__28445\,
            I => \b2v_inst6.un2_count_1_cry_1\
        );

    \I__5795\ : InMux
    port map (
            O => \N__28442\,
            I => \b2v_inst6.un2_count_1_cry_2\
        );

    \I__5794\ : InMux
    port map (
            O => \N__28439\,
            I => \b2v_inst6.un2_count_1_cry_3\
        );

    \I__5793\ : InMux
    port map (
            O => \N__28436\,
            I => \b2v_inst6.un2_count_1_cry_4\
        );

    \I__5792\ : InMux
    port map (
            O => \N__28433\,
            I => \b2v_inst6.un2_count_1_cry_5\
        );

    \I__5791\ : InMux
    port map (
            O => \N__28430\,
            I => \b2v_inst6.un2_count_1_cry_6\
        );

    \I__5790\ : InMux
    port map (
            O => \N__28427\,
            I => \b2v_inst6.un2_count_1_cry_7\
        );

    \I__5789\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28419\
        );

    \I__5788\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28414\
        );

    \I__5787\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28414\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__28419\,
            I => \N__28408\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__28414\,
            I => \N__28408\
        );

    \I__5784\ : InMux
    port map (
            O => \N__28413\,
            I => \N__28405\
        );

    \I__5783\ : Span4Mux_h
    port map (
            O => \N__28408\,
            I => \N__28402\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__28405\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__28402\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__5780\ : CascadeMux
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__5779\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28388\
        );

    \I__5778\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28388\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__28388\,
            I => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\
        );

    \I__5776\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28382\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__28382\,
            I => \b2v_inst11.count_clk_0_7\
        );

    \I__5774\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28376\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__28376\,
            I => \b2v_inst11.count_clk_0_10\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__28373\,
            I => \N__28370\
        );

    \I__5771\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28366\
        );

    \I__5770\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28363\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__28366\,
            I => \b2v_inst11.count_clk_1_10\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__28363\,
            I => \b2v_inst11.count_clk_1_10\
        );

    \I__5767\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__28355\,
            I => \b2v_inst11.count_clkZ0Z_13\
        );

    \I__5765\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28348\
        );

    \I__5764\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__28348\,
            I => \b2v_inst11.count_clkZ0Z_11\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__28345\,
            I => \b2v_inst11.count_clkZ0Z_11\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__28340\,
            I => \b2v_inst11.count_clkZ0Z_13_cascade_\
        );

    \I__5760\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28333\
        );

    \I__5759\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28330\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__28333\,
            I => \b2v_inst11.count_clkZ0Z_10\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__28330\,
            I => \b2v_inst11.count_clkZ0Z_10\
        );

    \I__5756\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__28322\,
            I => \N__28319\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__28319\,
            I => \b2v_inst11.un2_count_clk_17_0_o2_4\
        );

    \I__5753\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28312\
        );

    \I__5752\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28309\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__28312\,
            I => \b2v_inst11.count_clk_1_12\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__28309\,
            I => \b2v_inst11.count_clk_1_12\
        );

    \I__5749\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28301\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__28301\,
            I => \b2v_inst11.count_clk_0_12\
        );

    \I__5747\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28294\
        );

    \I__5746\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28291\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__28294\,
            I => \b2v_inst11.count_clkZ0Z_12\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__28291\,
            I => \b2v_inst11.count_clkZ0Z_12\
        );

    \I__5743\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28279\
        );

    \I__5742\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28279\
        );

    \I__5741\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28276\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__28279\,
            I => \N__28273\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__28276\,
            I => \b2v_inst11.func_state_enZ0\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__28273\,
            I => \b2v_inst11.func_state_enZ0\
        );

    \I__5737\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__28265\,
            I => \b2v_inst11.func_state_1_m2_1\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__5734\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28255\
        );

    \I__5733\ : InMux
    port map (
            O => \N__28258\,
            I => \N__28252\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__28255\,
            I => \b2v_inst11.func_stateZ0Z_1\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__28252\,
            I => \b2v_inst11.func_stateZ0Z_1\
        );

    \I__5730\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28243\
        );

    \I__5729\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28240\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__28243\,
            I => \N__28237\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28234\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__28237\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_5\
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__28234\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_5\
        );

    \I__5724\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28226\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__28226\,
            I => \b2v_inst11.func_state_1_m2s2_i_0\
        );

    \I__5722\ : InMux
    port map (
            O => \N__28223\,
            I => \N__28220\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28216\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__28219\,
            I => \N__28211\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__28216\,
            I => \N__28208\
        );

    \I__5718\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28205\
        );

    \I__5717\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28202\
        );

    \I__5716\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28199\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__28208\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__28205\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__28202\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__28199\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__5711\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28187\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__5709\ : Span4Mux_s2_v
    port map (
            O => \N__28184\,
            I => \N__28181\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__28181\,
            I => \b2v_inst11.count_clk_RNIZ0Z_0\
        );

    \I__5707\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28174\
        );

    \I__5706\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28170\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__28174\,
            I => \N__28166\
        );

    \I__5704\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28163\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28160\
        );

    \I__5702\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28157\
        );

    \I__5701\ : Span12Mux_s7_h
    port map (
            O => \N__28166\,
            I => \N__28152\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__28163\,
            I => \N__28149\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__28160\,
            I => \N__28144\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__28157\,
            I => \N__28144\
        );

    \I__5697\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28139\
        );

    \I__5696\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28139\
        );

    \I__5695\ : Odrv12
    port map (
            O => \N__28152\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__28149\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__28144\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__28139\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__5691\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28123\
        );

    \I__5690\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28114\
        );

    \I__5689\ : InMux
    port map (
            O => \N__28128\,
            I => \N__28114\
        );

    \I__5688\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28114\
        );

    \I__5687\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28114\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__28123\,
            I => \N__28111\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__28114\,
            I => \N__28100\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__28111\,
            I => \N__28094\
        );

    \I__5683\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28091\
        );

    \I__5682\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28080\
        );

    \I__5681\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28080\
        );

    \I__5680\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28080\
        );

    \I__5679\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28080\
        );

    \I__5678\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28073\
        );

    \I__5677\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28073\
        );

    \I__5676\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28073\
        );

    \I__5675\ : Span4Mux_s2_v
    port map (
            O => \N__28100\,
            I => \N__28070\
        );

    \I__5674\ : InMux
    port map (
            O => \N__28099\,
            I => \N__28063\
        );

    \I__5673\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28063\
        );

    \I__5672\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28063\
        );

    \I__5671\ : Span4Mux_v
    port map (
            O => \N__28094\,
            I => \N__28060\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__28091\,
            I => \N__28057\
        );

    \I__5669\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28052\
        );

    \I__5668\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28052\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__28080\,
            I => \N__28043\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__28073\,
            I => \N__28043\
        );

    \I__5665\ : Span4Mux_s3_h
    port map (
            O => \N__28070\,
            I => \N__28043\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__28063\,
            I => \N__28043\
        );

    \I__5663\ : Span4Mux_h
    port map (
            O => \N__28060\,
            I => \N__28040\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__28057\,
            I => \N__28037\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__28052\,
            I => \N__28032\
        );

    \I__5660\ : Span4Mux_s2_v
    port map (
            O => \N__28043\,
            I => \N__28032\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__28040\,
            I => \b2v_inst11.func_state_RNINIV94_0_0\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__28037\,
            I => \b2v_inst11.func_state_RNINIV94_0_0\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__28032\,
            I => \b2v_inst11.func_state_RNINIV94_0_0\
        );

    \I__5656\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28022\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__28022\,
            I => \b2v_inst11.count_clk_0_0\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__28019\,
            I => \b2v_inst11.func_state_1_m2_ns_1_0_cascade_\
        );

    \I__5653\ : InMux
    port map (
            O => \N__28016\,
            I => \N__28010\
        );

    \I__5652\ : InMux
    port map (
            O => \N__28015\,
            I => \N__28010\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__28010\,
            I => \b2v_inst11.func_state_1_m2_0\
        );

    \I__5650\ : InMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__28004\,
            I => \b2v_inst11.N_327\
        );

    \I__5648\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27998\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__27998\,
            I => \N__27995\
        );

    \I__5646\ : Odrv4
    port map (
            O => \N__27995\,
            I => \b2v_inst11.func_state_1_m2_ns_1_1_1\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__27992\,
            I => \b2v_inst11.N_382_cascade_\
        );

    \I__5644\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27986\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__27986\,
            I => \b2v_inst11.un1_func_state25_6_0_2\
        );

    \I__5642\ : CascadeMux
    port map (
            O => \N__27983\,
            I => \N__27979\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__27982\,
            I => \N__27976\
        );

    \I__5640\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27971\
        );

    \I__5639\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27968\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__27975\,
            I => \N__27965\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__27974\,
            I => \N__27962\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__27971\,
            I => \N__27959\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27956\
        );

    \I__5634\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27951\
        );

    \I__5633\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27951\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__27959\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_0\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__27956\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_0\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__27951\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_0\
        );

    \I__5629\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27941\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__27941\,
            I => \N__27938\
        );

    \I__5627\ : Span4Mux_v
    port map (
            O => \N__27938\,
            I => \N__27935\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__27935\,
            I => \b2v_inst11.un1_func_state25_6_0_a3_1\
        );

    \I__5625\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27929\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27924\
        );

    \I__5623\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27919\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27927\,
            I => \N__27919\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__27924\,
            I => \b2v_inst11.N_406\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__27919\,
            I => \b2v_inst11.N_406\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__27914\,
            I => \N__27911\
        );

    \I__5618\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27908\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__27908\,
            I => \b2v_inst11.func_state_1_m2_ns_1_1\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__27905\,
            I => \b2v_inst11.func_state_1_m2_1_cascade_\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__27902\,
            I => \b2v_inst11.func_stateZ0Z_0_cascade_\
        );

    \I__5614\ : InMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__5612\ : Span4Mux_v
    port map (
            O => \N__27893\,
            I => \N__27890\
        );

    \I__5611\ : Odrv4
    port map (
            O => \N__27890\,
            I => \b2v_inst11.N_337\
        );

    \I__5610\ : CascadeMux
    port map (
            O => \N__27887\,
            I => \b2v_inst11.N_338_cascade_\
        );

    \I__5609\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27880\
        );

    \I__5608\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27877\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__27880\,
            I => \b2v_inst11.N_76\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__27877\,
            I => \b2v_inst11.N_76\
        );

    \I__5605\ : CascadeMux
    port map (
            O => \N__27872\,
            I => \b2v_inst11.N_406_cascade_\
        );

    \I__5604\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27863\
        );

    \I__5603\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27863\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__27863\,
            I => \b2v_inst11.func_stateZ1Z_0\
        );

    \I__5601\ : CascadeMux
    port map (
            O => \N__27860\,
            I => \b2v_inst11.func_state_enZ0_cascade_\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__27857\,
            I => \b2v_inst11.func_state_cascade_\
        );

    \I__5599\ : CascadeMux
    port map (
            O => \N__27854\,
            I => \N__27851\
        );

    \I__5598\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27848\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__27848\,
            I => \N__27845\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__27845\,
            I => \N__27841\
        );

    \I__5595\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27838\
        );

    \I__5594\ : Odrv4
    port map (
            O => \N__27841\,
            I => \b2v_inst11.N_428\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__27838\,
            I => \b2v_inst11.N_428\
        );

    \I__5592\ : CascadeMux
    port map (
            O => \N__27833\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0_cascade_\
        );

    \I__5591\ : InMux
    port map (
            O => \N__27830\,
            I => \N__27827\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__27827\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0\
        );

    \I__5589\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27818\
        );

    \I__5588\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27818\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__27815\,
            I => \N__27812\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__27812\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__27809\,
            I => \N__27804\
        );

    \I__5583\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27798\
        );

    \I__5582\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27798\
        );

    \I__5581\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27793\
        );

    \I__5580\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27793\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__27798\,
            I => \b2v_inst11.N_369\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__27793\,
            I => \b2v_inst11.N_369\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__27788\,
            I => \b2v_inst11.func_state_1_m2_ns_1_1_0_cascade_\
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__27785\,
            I => \N__27782\
        );

    \I__5575\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27779\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27776\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__27776\,
            I => \N__27773\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__27773\,
            I => \b2v_inst11.g0_i_a7_1_2\
        );

    \I__5571\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27766\
        );

    \I__5570\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27763\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__27766\,
            I => \N__27760\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__27763\,
            I => \N__27756\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__27760\,
            I => \N__27753\
        );

    \I__5566\ : InMux
    port map (
            O => \N__27759\,
            I => \N__27750\
        );

    \I__5565\ : Span12Mux_s7_h
    port map (
            O => \N__27756\,
            I => \N__27747\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__27753\,
            I => \b2v_inst16.curr_state_RNIUCAD1Z0Z_0\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__27750\,
            I => \b2v_inst16.curr_state_RNIUCAD1Z0Z_0\
        );

    \I__5562\ : Odrv12
    port map (
            O => \N__27747\,
            I => \b2v_inst16.curr_state_RNIUCAD1Z0Z_0\
        );

    \I__5561\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27737\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__27737\,
            I => \N__27731\
        );

    \I__5559\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27726\
        );

    \I__5558\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27726\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__27734\,
            I => \N__27723\
        );

    \I__5556\ : Span4Mux_v
    port map (
            O => \N__27731\,
            I => \N__27717\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27714\
        );

    \I__5554\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27709\
        );

    \I__5553\ : InMux
    port map (
            O => \N__27722\,
            I => \N__27709\
        );

    \I__5552\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27704\
        );

    \I__5551\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27704\
        );

    \I__5550\ : Span4Mux_h
    port map (
            O => \N__27717\,
            I => \N__27699\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__27714\,
            I => \N__27699\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__27709\,
            I => \N__27694\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27694\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__27699\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__5545\ : Odrv12
    port map (
            O => \N__27694\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__5544\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27683\
        );

    \I__5543\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27683\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__27683\,
            I => \N__27680\
        );

    \I__5541\ : Span4Mux_v
    port map (
            O => \N__27680\,
            I => \N__27677\
        );

    \I__5540\ : Span4Mux_v
    port map (
            O => \N__27677\,
            I => \N__27674\
        );

    \I__5539\ : Span4Mux_h
    port map (
            O => \N__27674\,
            I => \N__27671\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__27671\,
            I => \b2v_inst16.N_268\
        );

    \I__5537\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27665\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__27665\,
            I => \b2v_inst11.N_395\
        );

    \I__5535\ : InMux
    port map (
            O => \N__27662\,
            I => \N__27656\
        );

    \I__5534\ : InMux
    port map (
            O => \N__27661\,
            I => \N__27656\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__27656\,
            I => \b2v_inst11.N_159\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__27653\,
            I => \b2v_inst11.N_159_cascade_\
        );

    \I__5531\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27647\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__27647\,
            I => \N__27640\
        );

    \I__5529\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27637\
        );

    \I__5528\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27633\
        );

    \I__5527\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27628\
        );

    \I__5526\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27628\
        );

    \I__5525\ : Span4Mux_v
    port map (
            O => \N__27640\,
            I => \N__27623\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__27637\,
            I => \N__27623\
        );

    \I__5523\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27618\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__27633\,
            I => \N__27615\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__27628\,
            I => \N__27612\
        );

    \I__5520\ : Span4Mux_h
    port map (
            O => \N__27623\,
            I => \N__27609\
        );

    \I__5519\ : InMux
    port map (
            O => \N__27622\,
            I => \N__27606\
        );

    \I__5518\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27603\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__27618\,
            I => \b2v_inst11.N_425\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__27615\,
            I => \b2v_inst11.N_425\
        );

    \I__5515\ : Odrv4
    port map (
            O => \N__27612\,
            I => \b2v_inst11.N_425\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__27609\,
            I => \b2v_inst11.N_425\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__27606\,
            I => \b2v_inst11.N_425\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__27603\,
            I => \b2v_inst11.N_425\
        );

    \I__5511\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27587\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__27587\,
            I => \b2v_inst11.g2\
        );

    \I__5509\ : InMux
    port map (
            O => \N__27584\,
            I => \N__27581\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__27581\,
            I => \N__27576\
        );

    \I__5507\ : InMux
    port map (
            O => \N__27580\,
            I => \N__27570\
        );

    \I__5506\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27567\
        );

    \I__5505\ : Span4Mux_s3_h
    port map (
            O => \N__27576\,
            I => \N__27564\
        );

    \I__5504\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27561\
        );

    \I__5503\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27558\
        );

    \I__5502\ : InMux
    port map (
            O => \N__27573\,
            I => \N__27555\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__27570\,
            I => \N__27552\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__27567\,
            I => \b2v_inst11.N_366\
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__27564\,
            I => \b2v_inst11.N_366\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__27561\,
            I => \b2v_inst11.N_366\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__27558\,
            I => \b2v_inst11.N_366\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__27555\,
            I => \b2v_inst11.N_366\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__27552\,
            I => \b2v_inst11.N_366\
        );

    \I__5494\ : CascadeMux
    port map (
            O => \N__27539\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_0_cascade_\
        );

    \I__5493\ : CascadeMux
    port map (
            O => \N__27536\,
            I => \b2v_inst11.N_168_cascade_\
        );

    \I__5492\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27529\
        );

    \I__5491\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27524\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__27529\,
            I => \N__27521\
        );

    \I__5489\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27518\
        );

    \I__5488\ : CascadeMux
    port map (
            O => \N__27527\,
            I => \N__27515\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__27524\,
            I => \N__27509\
        );

    \I__5486\ : Span4Mux_v
    port map (
            O => \N__27521\,
            I => \N__27506\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__27518\,
            I => \N__27503\
        );

    \I__5484\ : InMux
    port map (
            O => \N__27515\,
            I => \N__27500\
        );

    \I__5483\ : CascadeMux
    port map (
            O => \N__27514\,
            I => \N__27496\
        );

    \I__5482\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27490\
        );

    \I__5481\ : InMux
    port map (
            O => \N__27512\,
            I => \N__27490\
        );

    \I__5480\ : Span4Mux_h
    port map (
            O => \N__27509\,
            I => \N__27487\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__27506\,
            I => \N__27480\
        );

    \I__5478\ : Span4Mux_v
    port map (
            O => \N__27503\,
            I => \N__27480\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__27500\,
            I => \N__27480\
        );

    \I__5476\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27473\
        );

    \I__5475\ : InMux
    port map (
            O => \N__27496\,
            I => \N__27473\
        );

    \I__5474\ : InMux
    port map (
            O => \N__27495\,
            I => \N__27473\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__27490\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__27487\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__27480\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__27473\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5469\ : InMux
    port map (
            O => \N__27464\,
            I => \N__27460\
        );

    \I__5468\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27455\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__27460\,
            I => \N__27452\
        );

    \I__5466\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27449\
        );

    \I__5465\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27446\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__27455\,
            I => \N__27442\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__27452\,
            I => \N__27437\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__27449\,
            I => \N__27437\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27434\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__27445\,
            I => \N__27429\
        );

    \I__5459\ : Span4Mux_v
    port map (
            O => \N__27442\,
            I => \N__27424\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__27437\,
            I => \N__27424\
        );

    \I__5457\ : Span12Mux_s3_h
    port map (
            O => \N__27434\,
            I => \N__27421\
        );

    \I__5456\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27414\
        );

    \I__5455\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27414\
        );

    \I__5454\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27414\
        );

    \I__5453\ : Odrv4
    port map (
            O => \N__27424\,
            I => \RSMRSTn_0\
        );

    \I__5452\ : Odrv12
    port map (
            O => \N__27421\,
            I => \RSMRSTn_0\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__27414\,
            I => \RSMRSTn_0\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__27407\,
            I => \b2v_inst11.count_clk_RNIDQ4A1Z0Z_6_cascade_\
        );

    \I__5449\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__27401\,
            I => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__27398\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_\
        );

    \I__5446\ : CascadeMux
    port map (
            O => \N__27395\,
            I => \b2v_inst11.N_186_i_cascade_\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__27392\,
            I => \b2v_inst11.N_115_f0_cascade_\
        );

    \I__5444\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27386\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__27386\,
            I => \b2v_inst11.N_381\
        );

    \I__5442\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27374\
        );

    \I__5441\ : InMux
    port map (
            O => \N__27382\,
            I => \N__27374\
        );

    \I__5440\ : InMux
    port map (
            O => \N__27381\,
            I => \N__27374\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__27374\,
            I => \N__27370\
        );

    \I__5438\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27367\
        );

    \I__5437\ : Odrv4
    port map (
            O => \N__27370\,
            I => \b2v_inst5.curr_state_RNIZ0Z_1\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__27367\,
            I => \b2v_inst5.curr_state_RNIZ0Z_1\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__5434\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27352\
        );

    \I__5433\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27352\
        );

    \I__5432\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27349\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__27352\,
            I => \b2v_inst5.N_2898_i\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__27349\,
            I => \b2v_inst5.N_2898_i\
        );

    \I__5429\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27336\
        );

    \I__5428\ : SRMux
    port map (
            O => \N__27343\,
            I => \N__27336\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__27342\,
            I => \N__27332\
        );

    \I__5426\ : SRMux
    port map (
            O => \N__27341\,
            I => \N__27326\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__27336\,
            I => \N__27320\
        );

    \I__5424\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27315\
        );

    \I__5423\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27315\
        );

    \I__5422\ : SRMux
    port map (
            O => \N__27331\,
            I => \N__27310\
        );

    \I__5421\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27297\
        );

    \I__5420\ : SRMux
    port map (
            O => \N__27329\,
            I => \N__27297\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27294\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__27325\,
            I => \N__27290\
        );

    \I__5417\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27284\
        );

    \I__5416\ : SRMux
    port map (
            O => \N__27323\,
            I => \N__27284\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__27320\,
            I => \N__27279\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__27315\,
            I => \N__27279\
        );

    \I__5413\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27274\
        );

    \I__5412\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27274\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__27310\,
            I => \N__27271\
        );

    \I__5410\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27262\
        );

    \I__5409\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27262\
        );

    \I__5408\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27262\
        );

    \I__5407\ : InMux
    port map (
            O => \N__27306\,
            I => \N__27262\
        );

    \I__5406\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27257\
        );

    \I__5405\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27257\
        );

    \I__5404\ : SRMux
    port map (
            O => \N__27303\,
            I => \N__27254\
        );

    \I__5403\ : SRMux
    port map (
            O => \N__27302\,
            I => \N__27251\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__27297\,
            I => \N__27248\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__27294\,
            I => \N__27245\
        );

    \I__5400\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27240\
        );

    \I__5399\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27240\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__27289\,
            I => \N__27237\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__27284\,
            I => \N__27232\
        );

    \I__5396\ : Span4Mux_s2_v
    port map (
            O => \N__27279\,
            I => \N__27232\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__27274\,
            I => \N__27229\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__27271\,
            I => \N__27226\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__27262\,
            I => \N__27221\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__27257\,
            I => \N__27221\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__27254\,
            I => \N__27210\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__27251\,
            I => \N__27207\
        );

    \I__5389\ : Span4Mux_v
    port map (
            O => \N__27248\,
            I => \N__27204\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__27245\,
            I => \N__27199\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__27240\,
            I => \N__27199\
        );

    \I__5386\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27196\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__27232\,
            I => \N__27193\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__27229\,
            I => \N__27190\
        );

    \I__5383\ : Span4Mux_v
    port map (
            O => \N__27226\,
            I => \N__27185\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__27221\,
            I => \N__27185\
        );

    \I__5381\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27174\
        );

    \I__5380\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27174\
        );

    \I__5379\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27174\
        );

    \I__5378\ : InMux
    port map (
            O => \N__27217\,
            I => \N__27174\
        );

    \I__5377\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27174\
        );

    \I__5376\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27169\
        );

    \I__5375\ : InMux
    port map (
            O => \N__27214\,
            I => \N__27169\
        );

    \I__5374\ : InMux
    port map (
            O => \N__27213\,
            I => \N__27166\
        );

    \I__5373\ : Odrv12
    port map (
            O => \N__27210\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5372\ : Odrv12
    port map (
            O => \N__27207\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5371\ : Odrv4
    port map (
            O => \N__27204\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__27199\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__27196\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__27193\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__27190\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5366\ : Odrv4
    port map (
            O => \N__27185\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__27174\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__27169\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__27166\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__27143\,
            I => \N__27136\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__27142\,
            I => \N__27132\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__27141\,
            I => \N__27127\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__27140\,
            I => \N__27123\
        );

    \I__5358\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27111\
        );

    \I__5357\ : InMux
    port map (
            O => \N__27136\,
            I => \N__27111\
        );

    \I__5356\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27111\
        );

    \I__5355\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27102\
        );

    \I__5354\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27102\
        );

    \I__5353\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27102\
        );

    \I__5352\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27102\
        );

    \I__5351\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27093\
        );

    \I__5350\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27093\
        );

    \I__5349\ : InMux
    port map (
            O => \N__27122\,
            I => \N__27093\
        );

    \I__5348\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27093\
        );

    \I__5347\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27086\
        );

    \I__5346\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27086\
        );

    \I__5345\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27086\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__27111\,
            I => \N__27081\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__27102\,
            I => \N__27081\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__27093\,
            I => \N__27074\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__27086\,
            I => \N__27074\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__27081\,
            I => \N__27074\
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__27074\,
            I => \b2v_inst11.N_172_i\
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__27071\,
            I => \N__27068\
        );

    \I__5337\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27065\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__27065\,
            I => \N__27062\
        );

    \I__5335\ : Span4Mux_h
    port map (
            O => \N__27062\,
            I => \N__27059\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__27059\,
            I => \b2v_inst11.un1_clk_100khz_2_i_o3_out\
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__27056\,
            I => \b2v_inst11.N_19_cascade_\
        );

    \I__5332\ : CascadeMux
    port map (
            O => \N__27053\,
            I => \rsmrstn_cascade_\
        );

    \I__5331\ : CascadeMux
    port map (
            O => \N__27050\,
            I => \N__27047\
        );

    \I__5330\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27039\
        );

    \I__5329\ : InMux
    port map (
            O => \N__27046\,
            I => \N__27039\
        );

    \I__5328\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27036\
        );

    \I__5327\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27033\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__27030\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__27036\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__27033\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__27030\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__5322\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27020\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__27020\,
            I => \N__27016\
        );

    \I__5320\ : InMux
    port map (
            O => \N__27019\,
            I => \N__27012\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__27016\,
            I => \N__27009\
        );

    \I__5318\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27006\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__27012\,
            I => \b2v_inst5.countZ0Z_9\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__27009\,
            I => \b2v_inst5.countZ0Z_9\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__27006\,
            I => \b2v_inst5.countZ0Z_9\
        );

    \I__5314\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26995\
        );

    \I__5313\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26992\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__26995\,
            I => \N__26989\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__26992\,
            I => \N__26984\
        );

    \I__5310\ : Span4Mux_v
    port map (
            O => \N__26989\,
            I => \N__26984\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__26984\,
            I => \b2v_inst5.un2_count_1_cry_8_THRU_CO\
        );

    \I__5308\ : CascadeMux
    port map (
            O => \N__26981\,
            I => \N__26976\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__26980\,
            I => \N__26970\
        );

    \I__5306\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26965\
        );

    \I__5305\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26965\
        );

    \I__5304\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26955\
        );

    \I__5303\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26955\
        );

    \I__5302\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26955\
        );

    \I__5301\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26952\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__26965\,
            I => \N__26949\
        );

    \I__5299\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26942\
        );

    \I__5298\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26942\
        );

    \I__5297\ : InMux
    port map (
            O => \N__26962\,
            I => \N__26942\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__26955\,
            I => \N__26935\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__26952\,
            I => \N__26928\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__26949\,
            I => \N__26928\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__26942\,
            I => \N__26928\
        );

    \I__5292\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26921\
        );

    \I__5291\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26921\
        );

    \I__5290\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26921\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26918\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__26935\,
            I => \b2v_inst5.N_1_i\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__26928\,
            I => \b2v_inst5.N_1_i\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__26921\,
            I => \b2v_inst5.N_1_i\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__26918\,
            I => \b2v_inst5.N_1_i\
        );

    \I__5284\ : InMux
    port map (
            O => \N__26909\,
            I => \N__26906\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__26906\,
            I => \b2v_inst5.count_rst_5\
        );

    \I__5282\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26899\
        );

    \I__5281\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26896\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__26899\,
            I => \N__26893\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__26896\,
            I => \N__26890\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__26893\,
            I => \N__26885\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__26890\,
            I => \N__26885\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__26885\,
            I => \b2v_inst5.count_rst_9\
        );

    \I__5275\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26879\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__26876\,
            I => \b2v_inst5.count_1_5\
        );

    \I__5272\ : InMux
    port map (
            O => \N__26873\,
            I => \N__26869\
        );

    \I__5271\ : CEMux
    port map (
            O => \N__26872\,
            I => \N__26866\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__26869\,
            I => \N__26858\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__26866\,
            I => \N__26858\
        );

    \I__5268\ : CEMux
    port map (
            O => \N__26865\,
            I => \N__26852\
        );

    \I__5267\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26849\
        );

    \I__5266\ : CEMux
    port map (
            O => \N__26863\,
            I => \N__26845\
        );

    \I__5265\ : Span4Mux_h
    port map (
            O => \N__26858\,
            I => \N__26842\
        );

    \I__5264\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26835\
        );

    \I__5263\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26835\
        );

    \I__5262\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26835\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__26852\,
            I => \N__26832\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__26849\,
            I => \N__26829\
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__26848\,
            I => \N__26822\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__26845\,
            I => \N__26816\
        );

    \I__5257\ : Span4Mux_s2_h
    port map (
            O => \N__26842\,
            I => \N__26808\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__26835\,
            I => \N__26808\
        );

    \I__5255\ : Span4Mux_v
    port map (
            O => \N__26832\,
            I => \N__26803\
        );

    \I__5254\ : Span4Mux_v
    port map (
            O => \N__26829\,
            I => \N__26803\
        );

    \I__5253\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26787\
        );

    \I__5252\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26787\
        );

    \I__5251\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26787\
        );

    \I__5250\ : InMux
    port map (
            O => \N__26825\,
            I => \N__26787\
        );

    \I__5249\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26782\
        );

    \I__5248\ : CEMux
    port map (
            O => \N__26821\,
            I => \N__26782\
        );

    \I__5247\ : CEMux
    port map (
            O => \N__26820\,
            I => \N__26779\
        );

    \I__5246\ : CEMux
    port map (
            O => \N__26819\,
            I => \N__26776\
        );

    \I__5245\ : Sp12to4
    port map (
            O => \N__26816\,
            I => \N__26773\
        );

    \I__5244\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26766\
        );

    \I__5243\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26766\
        );

    \I__5242\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26766\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__26808\,
            I => \N__26763\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__26803\,
            I => \N__26760\
        );

    \I__5239\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26755\
        );

    \I__5238\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26755\
        );

    \I__5237\ : CEMux
    port map (
            O => \N__26800\,
            I => \N__26744\
        );

    \I__5236\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26744\
        );

    \I__5235\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26744\
        );

    \I__5234\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26744\
        );

    \I__5233\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26744\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__26787\,
            I => \N__26741\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__26782\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__26779\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__26776\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5228\ : Odrv12
    port map (
            O => \N__26773\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__26766\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__26763\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__26760\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__26755\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__26744\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__26741\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__26720\,
            I => \b2v_inst5.curr_stateZ0Z_0_cascade_\
        );

    \I__5220\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26714\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__26714\,
            I => \b2v_inst5.m4_0\
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__26711\,
            I => \b2v_inst5.N_2898_i_cascade_\
        );

    \I__5217\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26699\
        );

    \I__5216\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26699\
        );

    \I__5215\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26699\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N_413\
        );

    \I__5213\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26693\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__26693\,
            I => \b2v_inst5.curr_state_0_0\
        );

    \I__5211\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26681\
        );

    \I__5210\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26681\
        );

    \I__5209\ : InMux
    port map (
            O => \N__26688\,
            I => \N__26681\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__26681\,
            I => \b2v_inst5.curr_stateZ0Z_0\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__26678\,
            I => \b2v_inst5.countZ0Z_9_cascade_\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__26675\,
            I => \N__26672\
        );

    \I__5205\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26669\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__26669\,
            I => \b2v_inst5.count_1_9\
        );

    \I__5203\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26660\
        );

    \I__5202\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26660\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__26654\,
            I => \b2v_inst5.un2_count_1_cry_9_THRU_CO\
        );

    \I__5198\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__26648\,
            I => \N__26644\
        );

    \I__5196\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26641\
        );

    \I__5195\ : Span4Mux_h
    port map (
            O => \N__26644\,
            I => \N__26638\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__26641\,
            I => \b2v_inst5.un2_count_1_axb_10\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__26638\,
            I => \b2v_inst5.un2_count_1_axb_10\
        );

    \I__5192\ : InMux
    port map (
            O => \N__26633\,
            I => \N__26627\
        );

    \I__5191\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26627\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__26627\,
            I => \b2v_inst5.count_rst_4\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__26624\,
            I => \b2v_inst5.curr_stateZ0Z_1_cascade_\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__26621\,
            I => \b2v_inst5.curr_state_RNIZ0Z_1_cascade_\
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__26618\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_\
        );

    \I__5186\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26611\
        );

    \I__5185\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26608\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__26611\,
            I => \N__26605\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__26608\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__5182\ : Odrv12
    port map (
            O => \N__26605\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__5181\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26594\
        );

    \I__5180\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26594\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__26594\,
            I => \N__26591\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__26591\,
            I => \b2v_inst5.count_rst\
        );

    \I__5177\ : InMux
    port map (
            O => \N__26588\,
            I => \N__26585\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__26585\,
            I => \b2v_inst5.count_1_15\
        );

    \I__5175\ : InMux
    port map (
            O => \N__26582\,
            I => \N__26579\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__26579\,
            I => \b2v_inst5.curr_stateZ0Z_1\
        );

    \I__5173\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26570\
        );

    \I__5172\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26570\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__26570\,
            I => \N__26567\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__26567\,
            I => \N__26564\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__26564\,
            I => \b2v_inst5.count_rst_11\
        );

    \I__5168\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__26558\,
            I => \b2v_inst5.count_1_3\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__26555\,
            I => \N__26552\
        );

    \I__5165\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26549\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__5163\ : Span4Mux_v
    port map (
            O => \N__26546\,
            I => \N__26543\
        );

    \I__5162\ : Odrv4
    port map (
            O => \N__26543\,
            I => \b2v_inst5.countZ0Z_3\
        );

    \I__5161\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26532\
        );

    \I__5159\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26529\
        );

    \I__5158\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26526\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__26532\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__26529\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__26526\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__5154\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26516\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__26516\,
            I => \N__26512\
        );

    \I__5152\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26509\
        );

    \I__5151\ : Span4Mux_h
    port map (
            O => \N__26512\,
            I => \N__26506\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__26509\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__5149\ : Odrv4
    port map (
            O => \N__26506\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__26501\,
            I => \b2v_inst5.countZ0Z_3_cascade_\
        );

    \I__5147\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__26495\,
            I => \N__26491\
        );

    \I__5145\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26488\
        );

    \I__5144\ : Span4Mux_h
    port map (
            O => \N__26491\,
            I => \N__26485\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__26488\,
            I => \b2v_inst5.countZ0Z_2\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__26485\,
            I => \b2v_inst5.countZ0Z_2\
        );

    \I__5141\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__26474\,
            I => \b2v_inst5.un12_clk_100khz_11\
        );

    \I__5138\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26468\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__5136\ : Odrv4
    port map (
            O => \N__26465\,
            I => \b2v_inst5.un12_clk_100khz_4\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__26462\,
            I => \b2v_inst5.un12_clk_100khz_5_cascade_\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__26459\,
            I => \b2v_inst5.un2_count_1_axb_10_cascade_\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__26456\,
            I => \N__26452\
        );

    \I__5132\ : CascadeMux
    port map (
            O => \N__26455\,
            I => \N__26449\
        );

    \I__5131\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26444\
        );

    \I__5130\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26444\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__26444\,
            I => \b2v_inst5.count_1_10\
        );

    \I__5128\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26438\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26435\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__26435\,
            I => \N__26432\
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__26432\,
            I => \b2v_inst5.un12_clk_100khz_1\
        );

    \I__5124\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__26426\,
            I => \N__26422\
        );

    \I__5122\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26419\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__26422\,
            I => \N__26416\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__26419\,
            I => \b2v_inst5.countZ0Z_5\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__26416\,
            I => \b2v_inst5.countZ0Z_5\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__26411\,
            I => \N__26408\
        );

    \I__5117\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26405\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__26405\,
            I => \b2v_inst5.un12_clk_100khz_9\
        );

    \I__5115\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__26399\,
            I => \N__26395\
        );

    \I__5113\ : InMux
    port map (
            O => \N__26398\,
            I => \N__26392\
        );

    \I__5112\ : Span4Mux_v
    port map (
            O => \N__26395\,
            I => \N__26389\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__26392\,
            I => \N__26386\
        );

    \I__5110\ : Span4Mux_v
    port map (
            O => \N__26389\,
            I => \N__26383\
        );

    \I__5109\ : Span4Mux_v
    port map (
            O => \N__26386\,
            I => \N__26380\
        );

    \I__5108\ : Odrv4
    port map (
            O => \N__26383\,
            I => \b2v_inst5.countZ0Z_6\
        );

    \I__5107\ : Odrv4
    port map (
            O => \N__26380\,
            I => \b2v_inst5.countZ0Z_6\
        );

    \I__5106\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__26372\,
            I => \b2v_inst5.un12_clk_100khz_12\
        );

    \I__5104\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26364\
        );

    \I__5103\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26359\
        );

    \I__5102\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26359\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__26364\,
            I => \b2v_inst36.count_rst_8\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__26359\,
            I => \b2v_inst36.count_rst_8\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__26354\,
            I => \b2v_inst36.countZ0Z_4_cascade_\
        );

    \I__5098\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26345\
        );

    \I__5097\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26345\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__26345\,
            I => \b2v_inst36.count_2_6\
        );

    \I__5095\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__26339\,
            I => \b2v_inst36.un12_clk_100khz_0\
        );

    \I__5093\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__26333\,
            I => \b2v_inst36.un2_count_1_axb_12\
        );

    \I__5091\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26324\
        );

    \I__5090\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26324\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__26324\,
            I => \b2v_inst36.count_2_12\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__5087\ : InMux
    port map (
            O => \N__26318\,
            I => \N__26313\
        );

    \I__5086\ : InMux
    port map (
            O => \N__26317\,
            I => \N__26308\
        );

    \I__5085\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26308\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__26313\,
            I => \b2v_inst36.count_rst_2\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__26308\,
            I => \b2v_inst36.count_rst_2\
        );

    \I__5082\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26300\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__26300\,
            I => \b2v_inst36.un12_clk_100khz_1\
        );

    \I__5080\ : InMux
    port map (
            O => \N__26297\,
            I => \N__26291\
        );

    \I__5079\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26291\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__5077\ : Span4Mux_v
    port map (
            O => \N__26288\,
            I => \N__26285\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__26285\,
            I => \b2v_inst5.count_rst_13\
        );

    \I__5075\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26279\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__26279\,
            I => \b2v_inst5.count_1_1\
        );

    \I__5073\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26270\
        );

    \I__5072\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26270\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__5070\ : Span4Mux_h
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__5069\ : Odrv4
    port map (
            O => \N__26264\,
            I => \b2v_inst5.count_rst_12\
        );

    \I__5068\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__26258\,
            I => \b2v_inst5.count_1_2\
        );

    \I__5066\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__26252\,
            I => \b2v_inst36.un12_clk_100khz_5\
        );

    \I__5064\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26246\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__26246\,
            I => \b2v_inst36.un12_clk_100khz_4\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__26243\,
            I => \b2v_inst36.un12_clk_100khz_6_cascade_\
        );

    \I__5061\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26237\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26234\
        );

    \I__5059\ : Span4Mux_v
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__26231\,
            I => \b2v_inst36.un12_clk_100khz_7\
        );

    \I__5057\ : InMux
    port map (
            O => \N__26228\,
            I => \N__26225\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__5055\ : Odrv12
    port map (
            O => \N__26222\,
            I => \b2v_inst36.un12_clk_100khz_9\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__26219\,
            I => \b2v_inst36.un12_clk_100khz_13_cascade_\
        );

    \I__5053\ : CascadeMux
    port map (
            O => \N__26216\,
            I => \b2v_inst36.N_1_i_cascade_\
        );

    \I__5052\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26210\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__26210\,
            I => \b2v_inst36.count_rst_4\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__26207\,
            I => \b2v_inst36.count_rst_4_cascade_\
        );

    \I__5049\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26201\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__26201\,
            I => \N__26197\
        );

    \I__5047\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26194\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__26197\,
            I => \b2v_inst36.un2_count_1_axb_10\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__26194\,
            I => \b2v_inst36.un2_count_1_axb_10\
        );

    \I__5044\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26183\
        );

    \I__5043\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26183\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26180\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__26180\,
            I => \b2v_inst36.un2_count_1_cry_9_THRU_CO\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__26177\,
            I => \b2v_inst36.un2_count_1_axb_10_cascade_\
        );

    \I__5039\ : CascadeMux
    port map (
            O => \N__26174\,
            I => \N__26166\
        );

    \I__5038\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26163\
        );

    \I__5037\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26156\
        );

    \I__5036\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26156\
        );

    \I__5035\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26156\
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__26169\,
            I => \N__26149\
        );

    \I__5033\ : InMux
    port map (
            O => \N__26166\,
            I => \N__26139\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__26163\,
            I => \N__26134\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__26156\,
            I => \N__26134\
        );

    \I__5030\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26127\
        );

    \I__5029\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26127\
        );

    \I__5028\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26124\
        );

    \I__5027\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26119\
        );

    \I__5026\ : InMux
    port map (
            O => \N__26149\,
            I => \N__26119\
        );

    \I__5025\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26112\
        );

    \I__5024\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26112\
        );

    \I__5023\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26112\
        );

    \I__5022\ : InMux
    port map (
            O => \N__26145\,
            I => \N__26103\
        );

    \I__5021\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26103\
        );

    \I__5020\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26103\
        );

    \I__5019\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26103\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__26139\,
            I => \N__26100\
        );

    \I__5017\ : Span4Mux_s1_v
    port map (
            O => \N__26134\,
            I => \N__26097\
        );

    \I__5016\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26092\
        );

    \I__5015\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26092\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__26127\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__26124\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__26119\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__26112\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__26103\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__26100\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__26097\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__26092\,
            I => \b2v_inst36.N_1_i\
        );

    \I__5006\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26069\
        );

    \I__5005\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26069\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__26069\,
            I => \b2v_inst36.count_2_10\
        );

    \I__5003\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26063\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__26063\,
            I => \b2v_inst36.un2_count_1_axb_6\
        );

    \I__5001\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26054\
        );

    \I__5000\ : InMux
    port map (
            O => \N__26059\,
            I => \N__26054\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__26054\,
            I => \b2v_inst36.count_rst_10\
        );

    \I__4998\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__26048\,
            I => \b2v_inst36.count_2_4\
        );

    \I__4996\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__26042\,
            I => \b2v_inst36.countZ0Z_4\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__26039\,
            I => \b2v_inst36.curr_stateZ0Z_0_cascade_\
        );

    \I__4993\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26033\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__26033\,
            I => \b2v_inst36.curr_state_0_0\
        );

    \I__4991\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26027\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__26027\,
            I => \b2v_inst36.curr_state_0_1\
        );

    \I__4989\ : InMux
    port map (
            O => \N__26024\,
            I => \N__26021\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__26021\,
            I => \b2v_inst36.curr_state_7_1\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__26018\,
            I => \b2v_inst36.curr_stateZ0Z_1_cascade_\
        );

    \I__4986\ : InMux
    port map (
            O => \N__26015\,
            I => \N__26012\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__4984\ : Span4Mux_v
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__26006\,
            I => \b2v_inst36.DSW_PWROK_0\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__4981\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25996\
        );

    \I__4980\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25993\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__25996\,
            I => \N__25990\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__25993\,
            I => \N__25987\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__25990\,
            I => \b2v_inst36.un2_count_1_cry_7_THRU_CO\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__25987\,
            I => \b2v_inst36.un2_count_1_cry_7_THRU_CO\
        );

    \I__4975\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__25979\,
            I => \b2v_inst36.count_2_8\
        );

    \I__4973\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25973\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__25973\,
            I => \b2v_inst36.count_rst_6\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__25970\,
            I => \N__25966\
        );

    \I__4970\ : CascadeMux
    port map (
            O => \N__25969\,
            I => \N__25963\
        );

    \I__4969\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25959\
        );

    \I__4968\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25956\
        );

    \I__4967\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25953\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__25959\,
            I => \N__25948\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__25956\,
            I => \N__25948\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__25953\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__25948\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__25943\,
            I => \b2v_inst36.countZ0Z_8_cascade_\
        );

    \I__4961\ : InMux
    port map (
            O => \N__25940\,
            I => \b2v_inst11.un1_count_clk_2_cry_10\
        );

    \I__4960\ : InMux
    port map (
            O => \N__25937\,
            I => \b2v_inst11.un1_count_clk_2_cry_11\
        );

    \I__4959\ : InMux
    port map (
            O => \N__25934\,
            I => \b2v_inst11.un1_count_clk_2_cry_12\
        );

    \I__4958\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25927\
        );

    \I__4957\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25924\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__25927\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__25924\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__4954\ : InMux
    port map (
            O => \N__25919\,
            I => \N__25913\
        );

    \I__4953\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25913\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__25913\,
            I => \b2v_inst11.count_clk_1_14\
        );

    \I__4951\ : InMux
    port map (
            O => \N__25910\,
            I => \b2v_inst11.un1_count_clk_2_cry_13\
        );

    \I__4950\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__25904\,
            I => \b2v_inst11.count_clkZ0Z_15\
        );

    \I__4948\ : InMux
    port map (
            O => \N__25901\,
            I => \b2v_inst11.un1_count_clk_2_cry_14\
        );

    \I__4947\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25892\
        );

    \I__4946\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25892\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__25892\,
            I => \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\
        );

    \I__4944\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25886\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__25886\,
            I => \b2v_inst11.count_clk_0_11\
        );

    \I__4942\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25879\
        );

    \I__4941\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25876\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__25879\,
            I => \b2v_inst11.count_clk_1_11\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__25876\,
            I => \b2v_inst11.count_clk_1_11\
        );

    \I__4938\ : CascadeMux
    port map (
            O => \N__25871\,
            I => \b2v_inst36.curr_state_7_0_cascade_\
        );

    \I__4937\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25865\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__25865\,
            I => \N__25860\
        );

    \I__4935\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25857\
        );

    \I__4934\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25854\
        );

    \I__4933\ : Odrv12
    port map (
            O => \N__25860\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__25857\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__25854\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__4930\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25841\
        );

    \I__4929\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25841\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__25841\,
            I => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\
        );

    \I__4927\ : InMux
    port map (
            O => \N__25838\,
            I => \b2v_inst11.un1_count_clk_2_cry_2\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__4925\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25827\
        );

    \I__4924\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25822\
        );

    \I__4923\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25822\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__25827\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__25822\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__25817\,
            I => \N__25814\
        );

    \I__4919\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25808\
        );

    \I__4918\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25808\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__25808\,
            I => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\
        );

    \I__4916\ : InMux
    port map (
            O => \N__25805\,
            I => \b2v_inst11.un1_count_clk_2_cry_3\
        );

    \I__4915\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25798\
        );

    \I__4914\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25795\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__25798\,
            I => \N__25792\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__25795\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__25792\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__4910\ : CascadeMux
    port map (
            O => \N__25787\,
            I => \N__25784\
        );

    \I__4909\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25778\
        );

    \I__4908\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25778\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__4906\ : Odrv4
    port map (
            O => \N__25775\,
            I => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\
        );

    \I__4905\ : InMux
    port map (
            O => \N__25772\,
            I => \b2v_inst11.un1_count_clk_2_cry_4\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__4903\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25761\
        );

    \I__4902\ : InMux
    port map (
            O => \N__25765\,
            I => \N__25756\
        );

    \I__4901\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25756\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__25761\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__25756\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__4897\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25742\
        );

    \I__4896\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25742\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__25742\,
            I => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\
        );

    \I__4894\ : InMux
    port map (
            O => \N__25739\,
            I => \b2v_inst11.un1_count_clk_2_cry_5\
        );

    \I__4893\ : InMux
    port map (
            O => \N__25736\,
            I => \b2v_inst11.un1_count_clk_2_cry_6\
        );

    \I__4892\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25729\
        );

    \I__4891\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25726\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__25729\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__25726\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__4888\ : CascadeMux
    port map (
            O => \N__25721\,
            I => \N__25718\
        );

    \I__4887\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25712\
        );

    \I__4886\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25712\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__25712\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\
        );

    \I__4884\ : InMux
    port map (
            O => \N__25709\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\
        );

    \I__4883\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25702\
        );

    \I__4882\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25699\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__25702\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__25699\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__4879\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25688\
        );

    \I__4878\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25688\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__25688\,
            I => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\
        );

    \I__4876\ : InMux
    port map (
            O => \N__25685\,
            I => \bfn_8_16_0_\
        );

    \I__4875\ : InMux
    port map (
            O => \N__25682\,
            I => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\
        );

    \I__4874\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__25676\,
            I => \b2v_inst11.count_clk_0_2\
        );

    \I__4872\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25670\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__25670\,
            I => \b2v_inst11.count_clk_0_3\
        );

    \I__4870\ : InMux
    port map (
            O => \N__25667\,
            I => \N__25664\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__25664\,
            I => \b2v_inst11.count_clk_0_4\
        );

    \I__4868\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25658\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__25658\,
            I => \b2v_inst11.count_clk_0_6\
        );

    \I__4866\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25650\
        );

    \I__4865\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25647\
        );

    \I__4864\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25644\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__25650\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__25647\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__25644\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__25637\,
            I => \N__25634\
        );

    \I__4859\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25628\
        );

    \I__4858\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25628\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__25628\,
            I => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\
        );

    \I__4856\ : InMux
    port map (
            O => \N__25625\,
            I => \b2v_inst11.un1_count_clk_2_cry_1\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__25622\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\
        );

    \I__4854\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25616\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__25616\,
            I => \N__25613\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__25613\,
            I => \b2v_inst11.count_clk_en_0\
        );

    \I__4851\ : CascadeMux
    port map (
            O => \N__25610\,
            I => \b2v_inst11.N_328_cascade_\
        );

    \I__4850\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25604\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__25604\,
            I => \N__25601\
        );

    \I__4848\ : Span12Mux_v
    port map (
            O => \N__25601\,
            I => \N__25598\
        );

    \I__4847\ : Odrv12
    port map (
            O => \N__25598\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_0\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__25595\,
            I => \b2v_inst11.count_clk_en_cascade_\
        );

    \I__4845\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__25589\,
            I => \N__25586\
        );

    \I__4843\ : Span4Mux_v
    port map (
            O => \N__25586\,
            I => \N__25583\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__25583\,
            I => \b2v_inst11.N_218\
        );

    \I__4841\ : CascadeMux
    port map (
            O => \N__25580\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_329_N_cascade_\
        );

    \I__4840\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25574\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__25574\,
            I => \b2v_inst11.un1_func_state25_6_0_0\
        );

    \I__4838\ : CascadeMux
    port map (
            O => \N__25571\,
            I => \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7_cascade_\
        );

    \I__4837\ : CascadeMux
    port map (
            O => \N__25568\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_\
        );

    \I__4836\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__25562\,
            I => \b2v_inst11.g0_4_2\
        );

    \I__4834\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25556\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__25556\,
            I => \b2v_inst11.g0_0_0\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__4831\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25544\
        );

    \I__4830\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25544\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__25544\,
            I => \N__25541\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__25541\,
            I => \b2v_inst11.un1_clk_100khz_36_and_i_o3_0_c_0\
        );

    \I__4827\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__25535\,
            I => \b2v_inst11.g0_0_0_1\
        );

    \I__4825\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25526\
        );

    \I__4824\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25526\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__25526\,
            I => \N__25523\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__25523\,
            I => \N__25518\
        );

    \I__4821\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25513\
        );

    \I__4820\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25513\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__25518\,
            I => \N__25509\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__25513\,
            I => \N__25506\
        );

    \I__4817\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25503\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__25509\,
            I => \b2v_inst11.func_state_RNI8H551Z0Z_0\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__25506\,
            I => \b2v_inst11.func_state_RNI8H551Z0Z_0\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__25503\,
            I => \b2v_inst11.func_state_RNI8H551Z0Z_0\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__25496\,
            I => \N__25493\
        );

    \I__4812\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25487\
        );

    \I__4811\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25487\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25484\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__25484\,
            I => \N__25480\
        );

    \I__4808\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25476\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__25480\,
            I => \N__25473\
        );

    \I__4806\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25470\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__25476\,
            I => \N__25467\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__25473\,
            I => \b2v_inst11.func_state_RNIDUQ02Z0Z_1\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__25470\,
            I => \b2v_inst11.func_state_RNIDUQ02Z0Z_1\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__25467\,
            I => \b2v_inst11.func_state_RNIDUQ02Z0Z_1\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__25460\,
            I => \N__25456\
        );

    \I__4800\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25444\
        );

    \I__4799\ : InMux
    port map (
            O => \N__25456\,
            I => \N__25444\
        );

    \I__4798\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25439\
        );

    \I__4797\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25439\
        );

    \I__4796\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25430\
        );

    \I__4795\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25430\
        );

    \I__4794\ : InMux
    port map (
            O => \N__25451\,
            I => \N__25430\
        );

    \I__4793\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25430\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__25449\,
            I => \N__25427\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__25444\,
            I => \N__25419\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__25439\,
            I => \N__25416\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__25430\,
            I => \N__25411\
        );

    \I__4788\ : InMux
    port map (
            O => \N__25427\,
            I => \N__25408\
        );

    \I__4787\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25403\
        );

    \I__4786\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25403\
        );

    \I__4785\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25398\
        );

    \I__4784\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25398\
        );

    \I__4783\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25395\
        );

    \I__4782\ : Span4Mux_v
    port map (
            O => \N__25419\,
            I => \N__25392\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__25416\,
            I => \N__25389\
        );

    \I__4780\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25384\
        );

    \I__4779\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25384\
        );

    \I__4778\ : Span4Mux_h
    port map (
            O => \N__25411\,
            I => \N__25381\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__25408\,
            I => \N__25368\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__25403\,
            I => \N__25368\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__25398\,
            I => \N__25368\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__25395\,
            I => \N__25368\
        );

    \I__4773\ : Span4Mux_h
    port map (
            O => \N__25392\,
            I => \N__25368\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__25389\,
            I => \N__25368\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__25384\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__25381\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__25368\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7\
        );

    \I__4768\ : CascadeMux
    port map (
            O => \N__25361\,
            I => \b2v_inst11.dutycycle_eena_5_d_1_1_cascade_\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__25358\,
            I => \b2v_inst11.dutycycle_eena_5_0_1_cascade_\
        );

    \I__4766\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25352\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__25352\,
            I => \N__25349\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__25349\,
            I => \b2v_inst11.un1_clk_100khz_36_and_i_0\
        );

    \I__4763\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25342\
        );

    \I__4762\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25339\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25334\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__25339\,
            I => \N__25334\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__25328\,
            I => \b2v_inst11.dutycycle_RNI2IQ6CZ0Z_7\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__25325\,
            I => \b2v_inst11.func_state_RNIDUQ02Z0Z_1_cascade_\
        );

    \I__4755\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25317\
        );

    \I__4754\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25313\
        );

    \I__4753\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25309\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25306\
        );

    \I__4751\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25303\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__25313\,
            I => \N__25298\
        );

    \I__4749\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25295\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__25309\,
            I => \N__25290\
        );

    \I__4747\ : Span4Mux_v
    port map (
            O => \N__25306\,
            I => \N__25290\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__25303\,
            I => \N__25287\
        );

    \I__4745\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25282\
        );

    \I__4744\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25282\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__25298\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__25295\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__25290\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__25287\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__25282\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__25271\,
            I => \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf0_cascade_\
        );

    \I__4737\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25265\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__25265\,
            I => \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf1\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__25262\,
            I => \b2v_inst11.N_14_0_cascade_\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__25259\,
            I => \N__25256\
        );

    \I__4733\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__25253\,
            I => \b2v_inst11.g2_i_2\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__25250\,
            I => \N__25247\
        );

    \I__4730\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25241\
        );

    \I__4729\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25241\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__25241\,
            I => \N__25235\
        );

    \I__4727\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25228\
        );

    \I__4726\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25228\
        );

    \I__4725\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25228\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__25235\,
            I => \b2v_inst11.func_state_RNI_6Z0Z_0\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__25228\,
            I => \b2v_inst11.func_state_RNI_6Z0Z_0\
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__25223\,
            I => \b2v_inst11.N_395_cascade_\
        );

    \I__4721\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25212\
        );

    \I__4720\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25207\
        );

    \I__4719\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25207\
        );

    \I__4718\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25204\
        );

    \I__4717\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25201\
        );

    \I__4716\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25198\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__25212\,
            I => \N__25193\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__25207\,
            I => \N__25190\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__25204\,
            I => \N__25187\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25182\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__25198\,
            I => \N__25182\
        );

    \I__4710\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25179\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__25196\,
            I => \N__25174\
        );

    \I__4708\ : Span4Mux_h
    port map (
            O => \N__25193\,
            I => \N__25171\
        );

    \I__4707\ : Span4Mux_h
    port map (
            O => \N__25190\,
            I => \N__25168\
        );

    \I__4706\ : Span4Mux_h
    port map (
            O => \N__25187\,
            I => \N__25161\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__25182\,
            I => \N__25161\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__25179\,
            I => \N__25161\
        );

    \I__4703\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25156\
        );

    \I__4702\ : InMux
    port map (
            O => \N__25177\,
            I => \N__25156\
        );

    \I__4701\ : InMux
    port map (
            O => \N__25174\,
            I => \N__25153\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__25171\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__25168\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__25161\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__25156\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__25153\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__25142\,
            I => \N__25135\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__25141\,
            I => \N__25131\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__25140\,
            I => \N__25128\
        );

    \I__4692\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25125\
        );

    \I__4691\ : InMux
    port map (
            O => \N__25138\,
            I => \N__25116\
        );

    \I__4690\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25116\
        );

    \I__4689\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25116\
        );

    \I__4688\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25116\
        );

    \I__4687\ : InMux
    port map (
            O => \N__25128\,
            I => \N__25113\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__25125\,
            I => \N__25104\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__25116\,
            I => \N__25104\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__25113\,
            I => \N__25104\
        );

    \I__4683\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25099\
        );

    \I__4682\ : InMux
    port map (
            O => \N__25111\,
            I => \N__25099\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__25104\,
            I => \N__25096\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__25099\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__25096\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__4678\ : CascadeMux
    port map (
            O => \N__25091\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__25088\,
            I => \N__25082\
        );

    \I__4676\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25076\
        );

    \I__4675\ : InMux
    port map (
            O => \N__25086\,
            I => \N__25071\
        );

    \I__4674\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25071\
        );

    \I__4673\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25068\
        );

    \I__4672\ : InMux
    port map (
            O => \N__25081\,
            I => \N__25065\
        );

    \I__4671\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25062\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__25079\,
            I => \N__25057\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__25076\,
            I => \N__25053\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__25071\,
            I => \N__25050\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__25068\,
            I => \N__25043\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__25065\,
            I => \N__25043\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__25062\,
            I => \N__25043\
        );

    \I__4664\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25038\
        );

    \I__4663\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25038\
        );

    \I__4662\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25030\
        );

    \I__4661\ : InMux
    port map (
            O => \N__25056\,
            I => \N__25030\
        );

    \I__4660\ : Span4Mux_h
    port map (
            O => \N__25053\,
            I => \N__25027\
        );

    \I__4659\ : Span4Mux_h
    port map (
            O => \N__25050\,
            I => \N__25020\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__25043\,
            I => \N__25020\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25020\
        );

    \I__4656\ : InMux
    port map (
            O => \N__25037\,
            I => \N__25017\
        );

    \I__4655\ : InMux
    port map (
            O => \N__25036\,
            I => \N__25012\
        );

    \I__4654\ : InMux
    port map (
            O => \N__25035\,
            I => \N__25012\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__25030\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__25027\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__25020\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__25017\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__25012\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__4648\ : CascadeMux
    port map (
            O => \N__25001\,
            I => \b2v_inst11.N_365_cascade_\
        );

    \I__4647\ : CascadeMux
    port map (
            O => \N__24998\,
            I => \b2v_inst11.N_366_cascade_\
        );

    \I__4646\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24988\
        );

    \I__4645\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24988\
        );

    \I__4644\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24983\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__24988\,
            I => \N__24980\
        );

    \I__4642\ : InMux
    port map (
            O => \N__24987\,
            I => \N__24977\
        );

    \I__4641\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24974\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__24983\,
            I => \N__24969\
        );

    \I__4639\ : Span4Mux_v
    port map (
            O => \N__24980\,
            I => \N__24969\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__24977\,
            I => \N__24964\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__24974\,
            I => \N__24964\
        );

    \I__4636\ : Span4Mux_v
    port map (
            O => \N__24969\,
            I => \N__24961\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__24964\,
            I => \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__24961\,
            I => \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1\
        );

    \I__4633\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24952\
        );

    \I__4632\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24947\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__24952\,
            I => \N__24944\
        );

    \I__4630\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24940\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__24950\,
            I => \N__24936\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__24947\,
            I => \N__24932\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__24944\,
            I => \N__24929\
        );

    \I__4626\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24926\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__24940\,
            I => \N__24923\
        );

    \I__4624\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24918\
        );

    \I__4623\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24918\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__24935\,
            I => \N__24913\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__24932\,
            I => \N__24908\
        );

    \I__4620\ : Span4Mux_h
    port map (
            O => \N__24929\,
            I => \N__24908\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__24926\,
            I => \N__24905\
        );

    \I__4618\ : Span4Mux_h
    port map (
            O => \N__24923\,
            I => \N__24902\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__24918\,
            I => \N__24899\
        );

    \I__4616\ : InMux
    port map (
            O => \N__24917\,
            I => \N__24896\
        );

    \I__4615\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24893\
        );

    \I__4614\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24890\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__24908\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__24905\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__24902\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__24899\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__24896\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__24893\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__24890\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__4606\ : CascadeMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__4605\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__24869\,
            I => \b2v_inst11.N_153_N\
        );

    \I__4603\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24860\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__24860\,
            I => \N__24857\
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__24857\,
            I => \b2v_inst11.g2_i_a6_0\
        );

    \I__4599\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24850\
        );

    \I__4598\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24847\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__24850\,
            I => \N__24844\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__24847\,
            I => \N__24841\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__24844\,
            I => \N__24838\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__24841\,
            I => \N__24835\
        );

    \I__4593\ : Span4Mux_h
    port map (
            O => \N__24838\,
            I => \N__24830\
        );

    \I__4592\ : Span4Mux_h
    port map (
            O => \N__24835\,
            I => \N__24830\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__24830\,
            I => \b2v_inst11.N_363\
        );

    \I__4590\ : InMux
    port map (
            O => \N__24827\,
            I => \N__24824\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__24824\,
            I => \N__24821\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__24821\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__24818\,
            I => \b2v_inst11.N_396_N_cascade_\
        );

    \I__4586\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \b2v_inst11.N_234_N_cascade_\
        );

    \I__4585\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__24806\,
            I => \b2v_inst11.dutycycle_eena_9\
        );

    \I__4582\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__24800\,
            I => \N__24796\
        );

    \I__4580\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24793\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__24796\,
            I => \b2v_inst11.dutycycle_rst_8\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__24793\,
            I => \b2v_inst11.dutycycle_rst_8\
        );

    \I__4577\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24782\
        );

    \I__4576\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24782\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__24782\,
            I => \b2v_inst11.dutycycleZ1Z_12\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__24779\,
            I => \b2v_inst11.dutycycle_eena_9_cascade_\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__4572\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__24770\,
            I => \b2v_inst11.N_234_N\
        );

    \I__4570\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24764\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__24764\,
            I => \b2v_inst11.dutycycle_eena_7\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__24761\,
            I => \N__24758\
        );

    \I__4567\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24755\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__24755\,
            I => \N__24751\
        );

    \I__4565\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24748\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__24751\,
            I => \b2v_inst11.dutycycleZ1Z_11\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__24748\,
            I => \b2v_inst11.dutycycleZ1Z_11\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__24743\,
            I => \b2v_inst11.dutycycle_eena_7_cascade_\
        );

    \I__4561\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24734\
        );

    \I__4560\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24734\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__24734\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUFZ0Z1\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__4557\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24722\
        );

    \I__4556\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24722\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__24722\,
            I => \N__24719\
        );

    \I__4554\ : Span4Mux_h
    port map (
            O => \N__24719\,
            I => \N__24716\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__24716\,
            I => \b2v_inst11.dutycycle_RNIT35D7Z0Z_13\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__24713\,
            I => \N__24708\
        );

    \I__4551\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24705\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__24711\,
            I => \N__24700\
        );

    \I__4549\ : InMux
    port map (
            O => \N__24708\,
            I => \N__24696\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__24705\,
            I => \N__24693\
        );

    \I__4547\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24690\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__24703\,
            I => \N__24685\
        );

    \I__4545\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24680\
        );

    \I__4544\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24680\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__24696\,
            I => \N__24677\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__24693\,
            I => \N__24671\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__24690\,
            I => \N__24671\
        );

    \I__4540\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24666\
        );

    \I__4539\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24666\
        );

    \I__4538\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24663\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24658\
        );

    \I__4536\ : Span4Mux_v
    port map (
            O => \N__24677\,
            I => \N__24658\
        );

    \I__4535\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24655\
        );

    \I__4534\ : Odrv4
    port map (
            O => \N__24671\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__24666\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__24663\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__24658\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__24655\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__4529\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__24635\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_11\
        );

    \I__4525\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24624\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__24631\,
            I => \N__24617\
        );

    \I__4523\ : InMux
    port map (
            O => \N__24630\,
            I => \N__24614\
        );

    \I__4522\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24609\
        );

    \I__4521\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24609\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__24627\,
            I => \N__24605\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__24624\,
            I => \N__24602\
        );

    \I__4518\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24599\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__24622\,
            I => \N__24592\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__24621\,
            I => \N__24589\
        );

    \I__4515\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24583\
        );

    \I__4514\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24583\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__24614\,
            I => \N__24580\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24577\
        );

    \I__4511\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24572\
        );

    \I__4510\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24572\
        );

    \I__4509\ : Span4Mux_v
    port map (
            O => \N__24602\,
            I => \N__24569\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__24599\,
            I => \N__24564\
        );

    \I__4507\ : InMux
    port map (
            O => \N__24598\,
            I => \N__24561\
        );

    \I__4506\ : InMux
    port map (
            O => \N__24597\,
            I => \N__24558\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__24596\,
            I => \N__24552\
        );

    \I__4504\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24543\
        );

    \I__4503\ : InMux
    port map (
            O => \N__24592\,
            I => \N__24543\
        );

    \I__4502\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24543\
        );

    \I__4501\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24543\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__24583\,
            I => \N__24540\
        );

    \I__4499\ : Span4Mux_h
    port map (
            O => \N__24580\,
            I => \N__24537\
        );

    \I__4498\ : Span4Mux_v
    port map (
            O => \N__24577\,
            I => \N__24530\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__24572\,
            I => \N__24530\
        );

    \I__4496\ : Span4Mux_s3_h
    port map (
            O => \N__24569\,
            I => \N__24530\
        );

    \I__4495\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24525\
        );

    \I__4494\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24525\
        );

    \I__4493\ : Span4Mux_v
    port map (
            O => \N__24564\,
            I => \N__24518\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__24561\,
            I => \N__24518\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__24558\,
            I => \N__24518\
        );

    \I__4490\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24511\
        );

    \I__4489\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24511\
        );

    \I__4488\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24511\
        );

    \I__4487\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24508\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__24543\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__24540\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__24537\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__24530\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__24525\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4481\ : Odrv4
    port map (
            O => \N__24518\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__24511\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__24508\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__4477\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24485\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__24482\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_5\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__24479\,
            I => \b2v_inst5.count_rst_6_cascade_\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__4472\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24469\
        );

    \I__4471\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24466\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__24469\,
            I => \b2v_inst5.un2_count_1_axb_8\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__24466\,
            I => \b2v_inst5.un2_count_1_axb_8\
        );

    \I__4468\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24455\
        );

    \I__4467\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24455\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__24455\,
            I => \b2v_inst5.un2_count_1_cry_7_THRU_CO\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__24452\,
            I => \b2v_inst5.un2_count_1_axb_8_cascade_\
        );

    \I__4464\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24443\
        );

    \I__4463\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24443\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__24443\,
            I => \b2v_inst5.count_1_8\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__24440\,
            I => \b2v_inst5.count_rst_10_cascade_\
        );

    \I__4460\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24434\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__24434\,
            I => \N__24429\
        );

    \I__4458\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24424\
        );

    \I__4457\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24424\
        );

    \I__4456\ : Span4Mux_h
    port map (
            O => \N__24429\,
            I => \N__24421\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__24424\,
            I => \b2v_inst5.countZ0Z_4\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__24421\,
            I => \b2v_inst5.countZ0Z_4\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__24416\,
            I => \N__24412\
        );

    \I__4452\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24407\
        );

    \I__4451\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24407\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__4448\ : Odrv4
    port map (
            O => \N__24401\,
            I => \b2v_inst5.un2_count_1_cry_3_THRU_CO\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__24398\,
            I => \b2v_inst5.countZ0Z_4_cascade_\
        );

    \I__4446\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__24392\,
            I => \b2v_inst5.count_1_4\
        );

    \I__4444\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24385\
        );

    \I__4443\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24382\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__24385\,
            I => \b2v_inst5.un2_count_1_cry_12_THRU_CO\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__24382\,
            I => \b2v_inst5.un2_count_1_cry_12_THRU_CO\
        );

    \I__4440\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24374\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__24374\,
            I => \b2v_inst5.count_rst_1\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__24371\,
            I => \b2v_inst5.countZ0Z_13_cascade_\
        );

    \I__4437\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__24365\,
            I => \b2v_inst5.count_1_13\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__24362\,
            I => \b2v_inst5.count_i_0_cascade_\
        );

    \I__4434\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24356\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__24356\,
            I => \b2v_inst5.count_rst_14\
        );

    \I__4432\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24347\
        );

    \I__4431\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24347\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__24347\,
            I => \b2v_inst5.count_1_0\
        );

    \I__4429\ : CascadeMux
    port map (
            O => \N__24344\,
            I => \b2v_inst5.count_rst_14_cascade_\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__4427\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24335\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__24335\,
            I => \b2v_inst5.un2_count_1_axb_0\
        );

    \I__4425\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24325\
        );

    \I__4423\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24322\
        );

    \I__4422\ : Odrv12
    port map (
            O => \N__24325\,
            I => \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__24322\,
            I => \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2\
        );

    \I__4420\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24314\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__24311\,
            I => \b2v_inst5.count_1_14\
        );

    \I__4417\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__24305\,
            I => \b2v_inst5.countZ0Z_14\
        );

    \I__4415\ : InMux
    port map (
            O => \N__24302\,
            I => \N__24296\
        );

    \I__4414\ : InMux
    port map (
            O => \N__24301\,
            I => \N__24296\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__24296\,
            I => \b2v_inst5.count_i_0\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__24293\,
            I => \b2v_inst5.countZ0Z_14_cascade_\
        );

    \I__4411\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24286\
        );

    \I__4410\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24283\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24280\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__24283\,
            I => \N__24277\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__24280\,
            I => \b2v_inst5.countZ0Z_12\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__24277\,
            I => \b2v_inst5.countZ0Z_12\
        );

    \I__4405\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__24269\,
            I => \N__24266\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__24266\,
            I => \b2v_inst5.count_rst_6\
        );

    \I__4402\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24257\
        );

    \I__4401\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24257\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__24257\,
            I => \N__24254\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__24254\,
            I => \b2v_inst36.count_rst\
        );

    \I__4398\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__24245\,
            I => \N__24242\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__24242\,
            I => \b2v_inst20.counter_1_cry_1_THRU_CO\
        );

    \I__4394\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24235\
        );

    \I__4393\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24232\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__24235\,
            I => \N__24229\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24223\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__24229\,
            I => \N__24223\
        );

    \I__4389\ : InMux
    port map (
            O => \N__24228\,
            I => \N__24220\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__24223\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__24220\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__24215\,
            I => \b2v_inst36.curr_state_RNI3E27Z0Z_0_cascade_\
        );

    \I__4385\ : IoInMux
    port map (
            O => \N__24212\,
            I => \N__24209\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__4383\ : Span4Mux_s3_h
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__24203\,
            I => \N__24200\
        );

    \I__4381\ : Span4Mux_v
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__24197\,
            I => dsw_pwrok
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__24194\,
            I => \N__24187\
        );

    \I__4378\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24176\
        );

    \I__4377\ : InMux
    port map (
            O => \N__24192\,
            I => \N__24176\
        );

    \I__4376\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24176\
        );

    \I__4375\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24176\
        );

    \I__4374\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24176\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24167\
        );

    \I__4372\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24164\
        );

    \I__4371\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24153\
        );

    \I__4370\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24153\
        );

    \I__4369\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24153\
        );

    \I__4368\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24153\
        );

    \I__4367\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24153\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__24167\,
            I => \N__24150\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__24164\,
            I => \N__24145\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__24153\,
            I => \N__24145\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__24150\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__24145\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4361\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__24137\,
            I => \N__24134\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__24134\,
            I => \N__24131\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__24131\,
            I => \b2v_inst20.counter_1_cry_2_THRU_CO\
        );

    \I__4357\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24125\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__24125\,
            I => \N__24121\
        );

    \I__4355\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24117\
        );

    \I__4354\ : Span4Mux_h
    port map (
            O => \N__24121\,
            I => \N__24114\
        );

    \I__4353\ : InMux
    port map (
            O => \N__24120\,
            I => \N__24111\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__24117\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__24114\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__24111\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__24104\,
            I => \N__24100\
        );

    \I__4348\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24094\
        );

    \I__4347\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24094\
        );

    \I__4346\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24091\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__24094\,
            I => \b2v_inst36.un2_count_1_axb_7\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__24091\,
            I => \b2v_inst36.un2_count_1_axb_7\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__24086\,
            I => \N__24083\
        );

    \I__4342\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24079\
        );

    \I__4341\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24076\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__24079\,
            I => \N__24073\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__24076\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__24073\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__4337\ : InMux
    port map (
            O => \N__24068\,
            I => \b2v_inst36.un2_count_1_cry_6\
        );

    \I__4336\ : InMux
    port map (
            O => \N__24065\,
            I => \bfn_8_4_0_\
        );

    \I__4335\ : InMux
    port map (
            O => \N__24062\,
            I => \b2v_inst36.un2_count_1_cry_8\
        );

    \I__4334\ : InMux
    port map (
            O => \N__24059\,
            I => \b2v_inst36.un2_count_1_cry_9\
        );

    \I__4333\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24051\
        );

    \I__4332\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24046\
        );

    \I__4331\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24046\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__24051\,
            I => \N__24043\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__24046\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__24043\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__24038\,
            I => \N__24034\
        );

    \I__4326\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24029\
        );

    \I__4325\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24029\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24026\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__24026\,
            I => \b2v_inst36.un2_count_1_cry_10_THRU_CO\
        );

    \I__4322\ : InMux
    port map (
            O => \N__24023\,
            I => \b2v_inst36.un2_count_1_cry_10\
        );

    \I__4321\ : InMux
    port map (
            O => \N__24020\,
            I => \b2v_inst36.un2_count_1_cry_11\
        );

    \I__4320\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24013\
        );

    \I__4319\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24010\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__24013\,
            I => \N__24007\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__24010\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__24007\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__4315\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23996\
        );

    \I__4314\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23996\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__23996\,
            I => \N__23993\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__23993\,
            I => \b2v_inst36.count_rst_1\
        );

    \I__4311\ : InMux
    port map (
            O => \N__23990\,
            I => \b2v_inst36.un2_count_1_cry_12\
        );

    \I__4310\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23983\
        );

    \I__4309\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23980\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23977\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__23980\,
            I => \b2v_inst36.countZ0Z_14\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__23977\,
            I => \b2v_inst36.countZ0Z_14\
        );

    \I__4305\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23966\
        );

    \I__4304\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23966\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__23966\,
            I => \N__23963\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__23963\,
            I => \N__23960\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__23960\,
            I => \b2v_inst36.count_rst_0\
        );

    \I__4300\ : InMux
    port map (
            O => \N__23957\,
            I => \b2v_inst36.un2_count_1_cry_13\
        );

    \I__4299\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23947\
        );

    \I__4297\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23944\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__23947\,
            I => \b2v_inst36.countZ0Z_15\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__23944\,
            I => \b2v_inst36.countZ0Z_15\
        );

    \I__4294\ : InMux
    port map (
            O => \N__23939\,
            I => \b2v_inst36.un2_count_1_cry_14\
        );

    \I__4293\ : InMux
    port map (
            O => \N__23936\,
            I => \N__23932\
        );

    \I__4292\ : InMux
    port map (
            O => \N__23935\,
            I => \N__23929\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__23932\,
            I => \b2v_inst36.count_2_0\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__23929\,
            I => \b2v_inst36.count_2_0\
        );

    \I__4289\ : InMux
    port map (
            O => \N__23924\,
            I => \N__23920\
        );

    \I__4288\ : InMux
    port map (
            O => \N__23923\,
            I => \N__23917\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__23920\,
            I => \b2v_inst36.count_rst_14\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__23917\,
            I => \b2v_inst36.count_rst_14\
        );

    \I__4285\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__23909\,
            I => \b2v_inst36.un2_count_1_axb_0\
        );

    \I__4283\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23903\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__23903\,
            I => \N__23900\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__23900\,
            I => \b2v_inst36.un2_count_1_axb_1\
        );

    \I__4280\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23888\
        );

    \I__4279\ : InMux
    port map (
            O => \N__23896\,
            I => \N__23888\
        );

    \I__4278\ : InMux
    port map (
            O => \N__23895\,
            I => \N__23888\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__23885\,
            I => \b2v_inst36.count_rst_13\
        );

    \I__4275\ : InMux
    port map (
            O => \N__23882\,
            I => \b2v_inst36.un2_count_1_cry_0\
        );

    \I__4274\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23874\
        );

    \I__4273\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23869\
        );

    \I__4272\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23869\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23866\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__23869\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__4269\ : Odrv4
    port map (
            O => \N__23866\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__4268\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23855\
        );

    \I__4267\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23855\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__23855\,
            I => \N__23852\
        );

    \I__4265\ : Odrv4
    port map (
            O => \N__23852\,
            I => \b2v_inst36.un2_count_1_cry_1_THRU_CO\
        );

    \I__4264\ : InMux
    port map (
            O => \N__23849\,
            I => \b2v_inst36.un2_count_1_cry_1\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__23846\,
            I => \N__23842\
        );

    \I__4262\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__4261\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23836\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23833\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__23836\,
            I => \b2v_inst36.un2_count_1_axb_3\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__23833\,
            I => \b2v_inst36.un2_count_1_axb_3\
        );

    \I__4257\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23822\
        );

    \I__4256\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23822\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__23822\,
            I => \N__23819\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__23819\,
            I => \b2v_inst36.un2_count_1_cry_2_THRU_CO\
        );

    \I__4253\ : InMux
    port map (
            O => \N__23816\,
            I => \b2v_inst36.un2_count_1_cry_2\
        );

    \I__4252\ : InMux
    port map (
            O => \N__23813\,
            I => \b2v_inst36.un2_count_1_cry_3\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__23810\,
            I => \N__23806\
        );

    \I__4250\ : CascadeMux
    port map (
            O => \N__23809\,
            I => \N__23803\
        );

    \I__4249\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23799\
        );

    \I__4248\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23796\
        );

    \I__4247\ : InMux
    port map (
            O => \N__23802\,
            I => \N__23793\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__23799\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__23796\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__23793\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__4243\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23783\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23779\
        );

    \I__4241\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23776\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__23779\,
            I => \b2v_inst36.un2_count_1_cry_4_THRU_CO\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__23776\,
            I => \b2v_inst36.un2_count_1_cry_4_THRU_CO\
        );

    \I__4238\ : InMux
    port map (
            O => \N__23771\,
            I => \b2v_inst36.un2_count_1_cry_4\
        );

    \I__4237\ : InMux
    port map (
            O => \N__23768\,
            I => \b2v_inst36.un2_count_1_cry_5\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__23765\,
            I => \b2v_inst36.countZ0Z_2_cascade_\
        );

    \I__4235\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23759\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__23759\,
            I => \b2v_inst36.count_2_2\
        );

    \I__4233\ : CascadeMux
    port map (
            O => \N__23756\,
            I => \b2v_inst36.count_rst_7_cascade_\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__23753\,
            I => \b2v_inst36.count_rst_9_cascade_\
        );

    \I__4231\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23747\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__23747\,
            I => \b2v_inst36.count_2_5\
        );

    \I__4229\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23738\
        );

    \I__4228\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23738\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__23738\,
            I => \b2v_inst36.count_2_7\
        );

    \I__4226\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23732\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__23732\,
            I => \b2v_inst36.count_rst_7\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__23729\,
            I => \b2v_inst36.countZ0Z_5_cascade_\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__23726\,
            I => \b2v_inst11.count_clkZ0Z_15_cascade_\
        );

    \I__4222\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23717\
        );

    \I__4221\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23717\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__23717\,
            I => \b2v_inst11.N_175\
        );

    \I__4219\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__23711\,
            I => \b2v_inst11.count_clk_0_14\
        );

    \I__4217\ : CascadeMux
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__4216\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23702\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__23702\,
            I => \b2v_inst11.count_clk_0_15\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__23699\,
            I => \b2v_inst36.un2_count_1_axb_3_cascade_\
        );

    \I__4213\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23693\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__23693\,
            I => \b2v_inst36.count_rst_11\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__23690\,
            I => \b2v_inst36.count_rst_11_cascade_\
        );

    \I__4210\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23681\
        );

    \I__4209\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23681\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__23681\,
            I => \b2v_inst36.count_2_3\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__23678\,
            I => \b2v_inst36.count_rst_12_cascade_\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__23675\,
            I => \N__23672\
        );

    \I__4205\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__23669\,
            I => \b2v_inst11.count_clk_0_9\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__23666\,
            I => \b2v_inst11.count_clkZ0Z_9_cascade_\
        );

    \I__4202\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23657\
        );

    \I__4201\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23657\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__23657\,
            I => \b2v_inst11.N_190\
        );

    \I__4199\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__23651\,
            I => \b2v_inst11.count_clk_0_5\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__23648\,
            I => \b2v_inst11.count_clkZ0Z_5_cascade_\
        );

    \I__4196\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__23642\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__23639\,
            I => \b2v_inst11.count_clkZ0Z_1_cascade_\
        );

    \I__4193\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__23633\,
            I => \b2v_inst11.count_clk_0_1\
        );

    \I__4191\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__23627\,
            I => \b2v_inst11.count_clk_0_8\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__23624\,
            I => \b2v_inst11.count_clkZ0Z_8_cascade_\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__23621\,
            I => \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__23618\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\
        );

    \I__4186\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__23612\,
            I => \b2v_inst11.N_379\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__23609\,
            I => \b2v_inst11.N_379_cascade_\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__23606\,
            I => \N__23602\
        );

    \I__4182\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23597\
        );

    \I__4181\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23597\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__23597\,
            I => \b2v_inst11.dutycycle_eena_13_0\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__23594\,
            I => \b2v_inst11.N_200_i_cascade_\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__23591\,
            I => \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1_cascade_\
        );

    \I__4177\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23582\
        );

    \I__4176\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23582\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__4174\ : Span4Mux_v
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__23576\,
            I => \b2v_inst11.dutycycle_eena_3\
        );

    \I__4172\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23565\
        );

    \I__4171\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23558\
        );

    \I__4170\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23558\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__23570\,
            I => \N__23555\
        );

    \I__4168\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23550\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__23568\,
            I => \N__23547\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__23565\,
            I => \N__23538\
        );

    \I__4165\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23533\
        );

    \I__4164\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23533\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23528\
        );

    \I__4162\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23525\
        );

    \I__4161\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23520\
        );

    \I__4160\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23520\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23517\
        );

    \I__4158\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23514\
        );

    \I__4157\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23511\
        );

    \I__4156\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23506\
        );

    \I__4155\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23506\
        );

    \I__4154\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23503\
        );

    \I__4153\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23498\
        );

    \I__4152\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23498\
        );

    \I__4151\ : Span4Mux_v
    port map (
            O => \N__23538\,
            I => \N__23493\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__23533\,
            I => \N__23493\
        );

    \I__4149\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23488\
        );

    \I__4148\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23488\
        );

    \I__4147\ : Span4Mux_h
    port map (
            O => \N__23528\,
            I => \N__23485\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__23525\,
            I => \N__23480\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__23520\,
            I => \N__23480\
        );

    \I__4144\ : Span4Mux_v
    port map (
            O => \N__23517\,
            I => \N__23475\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23475\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__23511\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__23506\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__23503\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__23498\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4138\ : Odrv4
    port map (
            O => \N__23493\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__23488\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__23485\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__23480\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__23475\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__4133\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23453\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__23453\,
            I => \b2v_inst11.un1_clk_100khz_32_and_i_0_c\
        );

    \I__4131\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23444\
        );

    \I__4130\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23444\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__23441\,
            I => \b2v_inst11.un1_clk_100khz_40_and_i_0_c\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__23438\,
            I => \N__23431\
        );

    \I__4126\ : InMux
    port map (
            O => \N__23437\,
            I => \N__23426\
        );

    \I__4125\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23426\
        );

    \I__4124\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23419\
        );

    \I__4123\ : InMux
    port map (
            O => \N__23434\,
            I => \N__23414\
        );

    \I__4122\ : InMux
    port map (
            O => \N__23431\,
            I => \N__23414\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__23426\,
            I => \N__23411\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__23425\,
            I => \N__23408\
        );

    \I__4119\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23405\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__23423\,
            I => \N__23402\
        );

    \I__4117\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23394\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23389\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23389\
        );

    \I__4114\ : Span4Mux_h
    port map (
            O => \N__23411\,
            I => \N__23386\
        );

    \I__4113\ : InMux
    port map (
            O => \N__23408\,
            I => \N__23383\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__23405\,
            I => \N__23380\
        );

    \I__4111\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23377\
        );

    \I__4110\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23366\
        );

    \I__4109\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23366\
        );

    \I__4108\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23366\
        );

    \I__4107\ : InMux
    port map (
            O => \N__23398\,
            I => \N__23366\
        );

    \I__4106\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23366\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23363\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__23389\,
            I => \N__23360\
        );

    \I__4103\ : Span4Mux_h
    port map (
            O => \N__23386\,
            I => \N__23355\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23355\
        );

    \I__4101\ : Odrv12
    port map (
            O => \N__23380\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__23377\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__23366\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__23363\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__23360\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__23355\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__4095\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__23339\,
            I => \b2v_inst11.mult1_un145_sum\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__23336\,
            I => \b2v_inst11.mult1_un145_sum_cascade_\
        );

    \I__4092\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__4090\ : Span4Mux_s3_v
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__23324\,
            I => \b2v_inst11.mult1_un145_sum_i\
        );

    \I__4088\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23318\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__23315\,
            I => \b2v_inst11.N_10\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__23312\,
            I => \b2v_inst11.dutycycleZ0Z_12_cascade_\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__4083\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23302\
        );

    \I__4082\ : InMux
    port map (
            O => \N__23305\,
            I => \N__23299\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__23302\,
            I => \N__23296\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__23299\,
            I => \N__23293\
        );

    \I__4079\ : Span4Mux_v
    port map (
            O => \N__23296\,
            I => \N__23290\
        );

    \I__4078\ : Span4Mux_h
    port map (
            O => \N__23293\,
            I => \N__23287\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__23290\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_13\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__23287\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_13\
        );

    \I__4075\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23276\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__23276\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_14\
        );

    \I__4072\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23270\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23267\
        );

    \I__4070\ : Odrv12
    port map (
            O => \N__23267\,
            I => \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__23264\,
            I => \b2v_inst11.dutycycle_set_1_cascade_\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__4067\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__23255\,
            I => \b2v_inst11.N_300\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__23252\,
            I => \b2v_inst11.N_300_0_cascade_\
        );

    \I__4064\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23246\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__23240\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29\
        );

    \I__4060\ : InMux
    port map (
            O => \N__23237\,
            I => \N__23234\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__23234\,
            I => \b2v_inst11.dutycycle_set_0_0\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__23231\,
            I => \b2v_inst11.dutycycle_set_0_0_cascade_\
        );

    \I__4057\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__4056\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23222\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__23222\,
            I => \b2v_inst11.dutycycle_0_6\
        );

    \I__4054\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23213\
        );

    \I__4053\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23213\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__23213\,
            I => \b2v_inst11.dutycycle_0_5\
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__4050\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__23204\,
            I => \b2v_inst11.dutycycle_set_1\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__23201\,
            I => \b2v_inst11.un1_clk_100khz_40_and_i_0_0_0_cascade_\
        );

    \I__4047\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23192\
        );

    \I__4046\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23192\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__23192\,
            I => \N__23189\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__23189\,
            I => \b2v_inst11.dutycycle_RNIT35D7Z0Z_4\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__23186\,
            I => \N__23183\
        );

    \I__4042\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23180\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__23180\,
            I => \N__23177\
        );

    \I__4040\ : Span4Mux_h
    port map (
            O => \N__23177\,
            I => \N__23174\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__23174\,
            I => \b2v_inst11.N_155_N\
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__23171\,
            I => \b2v_inst11.dutycycle_en_11_cascade_\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__23168\,
            I => \b2v_inst11.N_158_N_cascade_\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__23165\,
            I => \N__23162\
        );

    \I__4035\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__23159\,
            I => \b2v_inst11.dutycycle_RNIT35D7Z0Z_15\
        );

    \I__4033\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23150\
        );

    \I__4032\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23150\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__23147\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__23144\,
            I => \b2v_inst11.dutycycle_RNIT35D7Z0Z_15_cascade_\
        );

    \I__4028\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23135\
        );

    \I__4027\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23135\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__23132\,
            I => \b2v_inst11.dutycycleZ0Z_15\
        );

    \I__4024\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23123\
        );

    \I__4023\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23123\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__23123\,
            I => \b2v_inst11.dutycycleZ0Z_14\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__4020\ : InMux
    port map (
            O => \N__23117\,
            I => \N__23114\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__23114\,
            I => \b2v_inst11.dutycycle_en_11\
        );

    \I__4018\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23105\
        );

    \I__4017\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23105\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__23105\,
            I => \N__23102\
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__23102\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__4013\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23092\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \N__23088\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__23083\
        );

    \I__4010\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23080\
        );

    \I__4009\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23077\
        );

    \I__4008\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23073\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__23086\,
            I => \N__23070\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__23083\,
            I => \N__23065\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__23065\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23062\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__23076\,
            I => \N__23058\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__23073\,
            I => \N__23054\
        );

    \I__4001\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23051\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__23065\,
            I => \N__23048\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__23062\,
            I => \N__23045\
        );

    \I__3998\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23040\
        );

    \I__3997\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23040\
        );

    \I__3996\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23037\
        );

    \I__3995\ : Span4Mux_h
    port map (
            O => \N__23054\,
            I => \N__23032\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__23051\,
            I => \N__23032\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__23048\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__23045\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__23040\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__23037\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__23032\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3988\ : InMux
    port map (
            O => \N__23021\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11_cZ0\
        );

    \I__3987\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23012\
        );

    \I__3986\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23012\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__23012\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\
        );

    \I__3984\ : InMux
    port map (
            O => \N__23009\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_cZ0\
        );

    \I__3983\ : InMux
    port map (
            O => \N__23006\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_cZ0\
        );

    \I__3982\ : InMux
    port map (
            O => \N__23003\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14\
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__23000\,
            I => \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0_cascade_\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__22997\,
            I => \b2v_inst11.dutycycleZ0Z_3_cascade_\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \N__22991\
        );

    \I__3978\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22988\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__22988\,
            I => \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0\
        );

    \I__3976\ : InMux
    port map (
            O => \N__22985\,
            I => \N__22982\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__22979\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\
        );

    \I__3973\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__22973\,
            I => \b2v_inst11.dutycycle_e_1_3\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__22967\,
            I => \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__22964\,
            I => \b2v_inst11.dutycycle_e_1_3_cascade_\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__3967\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22953\
        );

    \I__3966\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22948\
        );

    \I__3965\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22948\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__22953\,
            I => \b2v_inst11.dutycycle_0_3\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__22948\,
            I => \b2v_inst11.dutycycle_0_3\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__22943\,
            I => \N__22940\
        );

    \I__3961\ : InMux
    port map (
            O => \N__22940\,
            I => \N__22934\
        );

    \I__3960\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22934\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__22931\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\
        );

    \I__3957\ : InMux
    port map (
            O => \N__22928\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3\
        );

    \I__3956\ : InMux
    port map (
            O => \N__22925\,
            I => \b2v_inst11.un1_dutycycle_94_cry_4\
        );

    \I__3955\ : InMux
    port map (
            O => \N__22922\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__22919\,
            I => \N__22909\
        );

    \I__3953\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22905\
        );

    \I__3952\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22900\
        );

    \I__3951\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22900\
        );

    \I__3950\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22895\
        );

    \I__3949\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22895\
        );

    \I__3948\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22892\
        );

    \I__3947\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22889\
        );

    \I__3946\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22886\
        );

    \I__3945\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22883\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__22905\,
            I => \N__22878\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__22900\,
            I => \N__22878\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__22895\,
            I => \N__22874\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__22892\,
            I => \N__22871\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__22889\,
            I => \N__22866\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__22886\,
            I => \N__22866\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__22883\,
            I => \N__22861\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__22878\,
            I => \N__22861\
        );

    \I__3936\ : InMux
    port map (
            O => \N__22877\,
            I => \N__22858\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__22874\,
            I => \N__22853\
        );

    \I__3934\ : Span4Mux_v
    port map (
            O => \N__22871\,
            I => \N__22853\
        );

    \I__3933\ : Span4Mux_h
    port map (
            O => \N__22866\,
            I => \N__22850\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__22861\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__22858\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__22853\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__22850\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__22841\,
            I => \N__22837\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__22840\,
            I => \N__22834\
        );

    \I__3926\ : InMux
    port map (
            O => \N__22837\,
            I => \N__22831\
        );

    \I__3925\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22828\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__22831\,
            I => \N__22823\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__22828\,
            I => \N__22823\
        );

    \I__3922\ : Span4Mux_h
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__22820\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\
        );

    \I__3920\ : InMux
    port map (
            O => \N__22817\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__22814\,
            I => \N__22810\
        );

    \I__3918\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22805\
        );

    \I__3917\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22805\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__22802\,
            I => \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9JZ0Z1\
        );

    \I__3914\ : InMux
    port map (
            O => \N__22799\,
            I => \bfn_7_8_0_\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__22796\,
            I => \N__22792\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__22795\,
            I => \N__22785\
        );

    \I__3911\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22782\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__22791\,
            I => \N__22765\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__22790\,
            I => \N__22762\
        );

    \I__3908\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22753\
        );

    \I__3907\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22753\
        );

    \I__3906\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22753\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22750\
        );

    \I__3904\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22747\
        );

    \I__3903\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22742\
        );

    \I__3902\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22742\
        );

    \I__3901\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22735\
        );

    \I__3900\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22735\
        );

    \I__3899\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22735\
        );

    \I__3898\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22732\
        );

    \I__3897\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22723\
        );

    \I__3896\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22723\
        );

    \I__3895\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22723\
        );

    \I__3894\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22723\
        );

    \I__3893\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22716\
        );

    \I__3892\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22716\
        );

    \I__3891\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22716\
        );

    \I__3890\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22707\
        );

    \I__3889\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22707\
        );

    \I__3888\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22707\
        );

    \I__3887\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22707\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__22753\,
            I => \N__22702\
        );

    \I__3885\ : Span4Mux_h
    port map (
            O => \N__22750\,
            I => \N__22702\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__22747\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__22742\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__22735\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__22732\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__22723\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__22716\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__22707\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__22702\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3876\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22679\
        );

    \I__3875\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22679\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__22673\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJZ0Z1\
        );

    \I__3871\ : InMux
    port map (
            O => \N__22670\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__22667\,
            I => \N__22662\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__22666\,
            I => \N__22654\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__22665\,
            I => \N__22651\
        );

    \I__3867\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22647\
        );

    \I__3866\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22643\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__22660\,
            I => \N__22638\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__22659\,
            I => \N__22632\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__22658\,
            I => \N__22628\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__22657\,
            I => \N__22625\
        );

    \I__3861\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22620\
        );

    \I__3860\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22620\
        );

    \I__3859\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22617\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__22647\,
            I => \N__22614\
        );

    \I__3857\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22611\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__22643\,
            I => \N__22608\
        );

    \I__3855\ : InMux
    port map (
            O => \N__22642\,
            I => \N__22603\
        );

    \I__3854\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22603\
        );

    \I__3853\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22596\
        );

    \I__3852\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22596\
        );

    \I__3851\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22596\
        );

    \I__3850\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22591\
        );

    \I__3849\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22591\
        );

    \I__3848\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22588\
        );

    \I__3847\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22583\
        );

    \I__3846\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22583\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__22620\,
            I => \N__22578\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22578\
        );

    \I__3843\ : Span4Mux_v
    port map (
            O => \N__22614\,
            I => \N__22575\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__22611\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__22608\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__22603\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__22596\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__22591\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__22588\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__22583\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__22578\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__22575\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__3833\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22550\
        );

    \I__3832\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22550\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__3830\ : Span4Mux_v
    port map (
            O => \N__22547\,
            I => \N__22544\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__22544\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJZ0Z1\
        );

    \I__3828\ : InMux
    port map (
            O => \N__22541\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9\
        );

    \I__3827\ : InMux
    port map (
            O => \N__22538\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10\
        );

    \I__3826\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__3824\ : Span4Mux_v
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__22526\,
            I => \b2v_inst5.un2_count_1_axb_11\
        );

    \I__3822\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22514\
        );

    \I__3821\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22514\
        );

    \I__3820\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22514\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__22511\,
            I => \b2v_inst5.count_rst_3\
        );

    \I__3817\ : InMux
    port map (
            O => \N__22508\,
            I => \b2v_inst5.un2_count_1_cry_10\
        );

    \I__3816\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22499\
        );

    \I__3815\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22499\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__22496\,
            I => \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2\
        );

    \I__3812\ : InMux
    port map (
            O => \N__22493\,
            I => \b2v_inst5.un2_count_1_cry_11\
        );

    \I__3811\ : InMux
    port map (
            O => \N__22490\,
            I => \b2v_inst5.un2_count_1_cry_12\
        );

    \I__3810\ : InMux
    port map (
            O => \N__22487\,
            I => \b2v_inst5.un2_count_1_cry_13\
        );

    \I__3809\ : InMux
    port map (
            O => \N__22484\,
            I => \b2v_inst5.un2_count_1_cry_14\
        );

    \I__3808\ : InMux
    port map (
            O => \N__22481\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__3807\ : InMux
    port map (
            O => \N__22478\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__3806\ : InMux
    port map (
            O => \N__22475\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2\
        );

    \I__3805\ : InMux
    port map (
            O => \N__22472\,
            I => \b2v_inst5.un2_count_1_cry_1\
        );

    \I__3804\ : InMux
    port map (
            O => \N__22469\,
            I => \b2v_inst5.un2_count_1_cry_2\
        );

    \I__3803\ : InMux
    port map (
            O => \N__22466\,
            I => \b2v_inst5.un2_count_1_cry_3\
        );

    \I__3802\ : InMux
    port map (
            O => \N__22463\,
            I => \b2v_inst5.un2_count_1_cry_4\
        );

    \I__3801\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22454\
        );

    \I__3800\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22454\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__3798\ : Span4Mux_v
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__22448\,
            I => \b2v_inst5.count_rst_8\
        );

    \I__3796\ : InMux
    port map (
            O => \N__22445\,
            I => \b2v_inst5.un2_count_1_cry_5\
        );

    \I__3795\ : InMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__3793\ : Odrv12
    port map (
            O => \N__22436\,
            I => \b2v_inst5.countZ0Z_7\
        );

    \I__3792\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22427\
        );

    \I__3791\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22427\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__22424\,
            I => \b2v_inst5.count_rst_7\
        );

    \I__3788\ : InMux
    port map (
            O => \N__22421\,
            I => \b2v_inst5.un2_count_1_cry_6\
        );

    \I__3787\ : InMux
    port map (
            O => \N__22418\,
            I => \bfn_7_6_0_\
        );

    \I__3786\ : InMux
    port map (
            O => \N__22415\,
            I => \b2v_inst5.un2_count_1_cry_8\
        );

    \I__3785\ : InMux
    port map (
            O => \N__22412\,
            I => \b2v_inst5.un2_count_1_cry_9\
        );

    \I__3784\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__22403\,
            I => \b2v_inst20.counter_1_cry_5_THRU_CO\
        );

    \I__3781\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22396\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__22399\,
            I => \N__22392\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22389\
        );

    \I__3778\ : InMux
    port map (
            O => \N__22395\,
            I => \N__22384\
        );

    \I__3777\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22384\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__22389\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__22384\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__3774\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22375\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__22378\,
            I => \N__22372\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__22375\,
            I => \N__22368\
        );

    \I__3771\ : InMux
    port map (
            O => \N__22372\,
            I => \N__22363\
        );

    \I__3770\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22363\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__22368\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__22363\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__3766\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22346\
        );

    \I__3764\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22339\
        );

    \I__3763\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22339\
        );

    \I__3762\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22339\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__22346\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__22339\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__3758\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__22325\,
            I => \b2v_inst20.un4_counter_0_and\
        );

    \I__3755\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__3753\ : Span4Mux_h
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__22313\,
            I => \b2v_inst20.counter_1_cry_4_THRU_CO\
        );

    \I__3751\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22302\
        );

    \I__3749\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22297\
        );

    \I__3748\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22297\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__22302\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__22297\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__3745\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__22289\,
            I => \N__22286\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__22286\,
            I => \b2v_inst20.counter_1_cry_3_THRU_CO\
        );

    \I__3742\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22279\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22275\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22272\
        );

    \I__3739\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22267\
        );

    \I__3738\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22267\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__22272\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__22267\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__3735\ : InMux
    port map (
            O => \N__22262\,
            I => \b2v_inst5.un2_count_1_cry_0\
        );

    \I__3734\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__22256\,
            I => \b2v_inst5.count_1_7\
        );

    \I__3732\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22247\
        );

    \I__3731\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22247\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__22247\,
            I => \b2v_inst5.count_1_11\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__22244\,
            I => \b2v_inst5.countZ0Z_7_cascade_\
        );

    \I__3728\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__22238\,
            I => \b2v_inst5.count_1_12\
        );

    \I__3726\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22231\
        );

    \I__3725\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22228\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22225\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__22228\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__22225\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__3720\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__3718\ : Odrv12
    port map (
            O => \N__22211\,
            I => \b2v_inst20.un4_counter_1_and\
        );

    \I__3717\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__22205\,
            I => \b2v_inst36.count_2_15\
        );

    \I__3715\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__22199\,
            I => \b2v_inst36.count_2_13\
        );

    \I__3713\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__22193\,
            I => \b2v_inst36.count_2_14\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__3710\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22182\
        );

    \I__3709\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22177\
        );

    \I__3708\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22177\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__22182\,
            I => \b2v_inst36.count_i_0\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__22177\,
            I => \b2v_inst36.count_i_0\
        );

    \I__3705\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__22169\,
            I => \b2v_inst11.mult1_un145_sum_cry_6_s\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__22166\,
            I => \N__22162\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__22165\,
            I => \N__22158\
        );

    \I__3701\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22151\
        );

    \I__3700\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22151\
        );

    \I__3699\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22151\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__22151\,
            I => \b2v_inst11.mult1_un145_sum_i_0_8\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__3696\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__22142\,
            I => \b2v_inst11.mult1_un159_sum_axb_7\
        );

    \I__3694\ : InMux
    port map (
            O => \N__22139\,
            I => \b2v_inst11.mult1_un152_sum_cry_6\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__3692\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22130\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__22130\,
            I => \b2v_inst11.mult1_un152_sum_axb_8\
        );

    \I__3690\ : InMux
    port map (
            O => \N__22127\,
            I => \b2v_inst11.mult1_un152_sum_cry_7\
        );

    \I__3689\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22117\
        );

    \I__3687\ : CascadeMux
    port map (
            O => \N__22120\,
            I => \N__22113\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__22117\,
            I => \N__22109\
        );

    \I__3685\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22104\
        );

    \I__3684\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22104\
        );

    \I__3683\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22101\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__22109\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__22104\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__22101\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__22094\,
            I => \b2v_inst11.mult1_un152_sum_s_8_cascade_\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__22091\,
            I => \N__22087\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__22090\,
            I => \N__22083\
        );

    \I__3676\ : InMux
    port map (
            O => \N__22087\,
            I => \N__22076\
        );

    \I__3675\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22076\
        );

    \I__3674\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22076\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__22076\,
            I => \b2v_inst11.mult1_un152_sum_i_0_8\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__22073\,
            I => \b2v_inst36.count_rst_3_cascade_\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__22070\,
            I => \b2v_inst36.countZ0Z_11_cascade_\
        );

    \I__3670\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__22064\,
            I => \b2v_inst36.count_2_11\
        );

    \I__3668\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22055\
        );

    \I__3667\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22055\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__22055\,
            I => \b2v_inst36.count_2_1\
        );

    \I__3665\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__22049\,
            I => \b2v_inst11.mult1_un138_sum_cry_6_s\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__22046\,
            I => \N__22042\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__22045\,
            I => \N__22038\
        );

    \I__3661\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22031\
        );

    \I__3660\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22031\
        );

    \I__3659\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22031\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__22031\,
            I => \b2v_inst11.mult1_un138_sum_i_0_8\
        );

    \I__3657\ : InMux
    port map (
            O => \N__22028\,
            I => \b2v_inst11.mult1_un145_sum_cry_6\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__3655\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22019\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__22019\,
            I => \b2v_inst11.mult1_un145_sum_axb_8\
        );

    \I__3653\ : InMux
    port map (
            O => \N__22016\,
            I => \b2v_inst11.mult1_un145_sum_cry_7\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__22013\,
            I => \b2v_inst11.mult1_un145_sum_s_8_cascade_\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__3650\ : InMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__22004\,
            I => \b2v_inst11.mult1_un152_sum_cry_3_s\
        );

    \I__3648\ : InMux
    port map (
            O => \N__22001\,
            I => \b2v_inst11.mult1_un152_sum_cry_2\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__3646\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__21992\,
            I => \b2v_inst11.mult1_un145_sum_cry_3_s\
        );

    \I__3644\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__21986\,
            I => \b2v_inst11.mult1_un152_sum_cry_4_s\
        );

    \I__3642\ : InMux
    port map (
            O => \N__21983\,
            I => \b2v_inst11.mult1_un152_sum_cry_3\
        );

    \I__3641\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__21977\,
            I => \b2v_inst11.mult1_un145_sum_cry_4_s\
        );

    \I__3639\ : CascadeMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__3638\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__21968\,
            I => \b2v_inst11.mult1_un152_sum_cry_5_s\
        );

    \I__3636\ : InMux
    port map (
            O => \N__21965\,
            I => \b2v_inst11.mult1_un152_sum_cry_4\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__3634\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21955\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__21958\,
            I => \N__21951\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__21955\,
            I => \N__21947\
        );

    \I__3631\ : InMux
    port map (
            O => \N__21954\,
            I => \N__21942\
        );

    \I__3630\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21942\
        );

    \I__3629\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21939\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__21947\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__21942\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__21939\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__3624\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__21926\,
            I => \b2v_inst11.mult1_un145_sum_cry_5_s\
        );

    \I__3622\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__21920\,
            I => \b2v_inst11.mult1_un152_sum_cry_6_s\
        );

    \I__3620\ : InMux
    port map (
            O => \N__21917\,
            I => \b2v_inst11.mult1_un152_sum_cry_5\
        );

    \I__3619\ : InMux
    port map (
            O => \N__21914\,
            I => \b2v_inst11.mult1_un138_sum_cry_5_c\
        );

    \I__3618\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21908\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__21908\,
            I => \b2v_inst11.mult1_un131_sum_cry_6_s\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__21905\,
            I => \N__21901\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__21904\,
            I => \N__21897\
        );

    \I__3614\ : InMux
    port map (
            O => \N__21901\,
            I => \N__21890\
        );

    \I__3613\ : InMux
    port map (
            O => \N__21900\,
            I => \N__21890\
        );

    \I__3612\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21890\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__21890\,
            I => \b2v_inst11.mult1_un131_sum_i_0_8\
        );

    \I__3610\ : InMux
    port map (
            O => \N__21887\,
            I => \b2v_inst11.mult1_un138_sum_cry_6_c\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__3608\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21878\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__21878\,
            I => \b2v_inst11.mult1_un138_sum_axb_8\
        );

    \I__3606\ : InMux
    port map (
            O => \N__21875\,
            I => \b2v_inst11.mult1_un138_sum_cry_7\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__21872\,
            I => \b2v_inst11.mult1_un138_sum_s_8_cascade_\
        );

    \I__3604\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__3602\ : Odrv12
    port map (
            O => \N__21863\,
            I => \b2v_inst11.mult1_un138_sum_i\
        );

    \I__3601\ : InMux
    port map (
            O => \N__21860\,
            I => \b2v_inst11.mult1_un145_sum_cry_2\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__3599\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__21851\,
            I => \b2v_inst11.mult1_un138_sum_cry_3_s\
        );

    \I__3597\ : InMux
    port map (
            O => \N__21848\,
            I => \b2v_inst11.mult1_un145_sum_cry_3\
        );

    \I__3596\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__21842\,
            I => \b2v_inst11.mult1_un138_sum_cry_4_s\
        );

    \I__3594\ : InMux
    port map (
            O => \N__21839\,
            I => \b2v_inst11.mult1_un145_sum_cry_4\
        );

    \I__3593\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21832\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__21835\,
            I => \N__21828\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__21832\,
            I => \N__21824\
        );

    \I__3590\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21819\
        );

    \I__3589\ : InMux
    port map (
            O => \N__21828\,
            I => \N__21819\
        );

    \I__3588\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21816\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__21824\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__21819\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__21816\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__3584\ : CascadeMux
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__3583\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__21803\,
            I => \b2v_inst11.mult1_un138_sum_cry_5_s\
        );

    \I__3581\ : InMux
    port map (
            O => \N__21800\,
            I => \b2v_inst11.mult1_un145_sum_cry_5\
        );

    \I__3580\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__21794\,
            I => \b2v_inst5.count_1_6\
        );

    \I__3578\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__21776\,
            I => vr_ready_vccinaux
        );

    \I__3572\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__3570\ : Span12Mux_s7_v
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__3569\ : Odrv12
    port map (
            O => \N__21764\,
            I => vr_ready_vccin
        );

    \I__3568\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21754\
        );

    \I__3566\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21751\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__21754\,
            I => \b2v_inst11.mult1_un124_sum_cry_3_s\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__21751\,
            I => \b2v_inst11.mult1_un124_sum_cry_3_s\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__21746\,
            I => \N__21741\
        );

    \I__3562\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21737\
        );

    \I__3561\ : InMux
    port map (
            O => \N__21744\,
            I => \N__21731\
        );

    \I__3560\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21731\
        );

    \I__3559\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21728\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__21737\,
            I => \N__21724\
        );

    \I__3557\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21721\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__21731\,
            I => \N__21716\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__21728\,
            I => \N__21716\
        );

    \I__3554\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21713\
        );

    \I__3553\ : Odrv12
    port map (
            O => \N__21724\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__21721\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__21716\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__21713\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__3548\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__21698\,
            I => \b2v_inst11.mult1_un131_sum_axb_4_l_fx\
        );

    \I__3546\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21691\
        );

    \I__3545\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21688\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__21691\,
            I => \N__21683\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__21688\,
            I => \N__21683\
        );

    \I__3542\ : Odrv12
    port map (
            O => \N__21683\,
            I => \b2v_inst11.mult1_un138_sum\
        );

    \I__3541\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__3539\ : Odrv12
    port map (
            O => \N__21674\,
            I => \b2v_inst11.mult1_un131_sum_i\
        );

    \I__3538\ : InMux
    port map (
            O => \N__21671\,
            I => \b2v_inst11.mult1_un138_sum_cry_2_c\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__3536\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__21662\,
            I => \b2v_inst11.mult1_un131_sum_cry_3_s\
        );

    \I__3534\ : InMux
    port map (
            O => \N__21659\,
            I => \b2v_inst11.mult1_un138_sum_cry_3_c\
        );

    \I__3533\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__21653\,
            I => \b2v_inst11.mult1_un131_sum_cry_4_s\
        );

    \I__3531\ : InMux
    port map (
            O => \N__21650\,
            I => \b2v_inst11.mult1_un138_sum_cry_4_c\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__21647\,
            I => \N__21642\
        );

    \I__3529\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21638\
        );

    \I__3528\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21633\
        );

    \I__3527\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21633\
        );

    \I__3526\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21630\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__21638\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__21633\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__21630\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__3521\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21617\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__21617\,
            I => \b2v_inst11.mult1_un131_sum_cry_5_s\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__3518\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__21608\,
            I => \N__21605\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__21605\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_13\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__21602\,
            I => \N__21598\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__21601\,
            I => \N__21595\
        );

    \I__3513\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21590\
        );

    \I__3512\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21590\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__21590\,
            I => \b2v_inst11.mult1_un47_sum\
        );

    \I__3510\ : InMux
    port map (
            O => \N__21587\,
            I => \b2v_inst11.un1_dutycycle_53_cry_13\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__21584\,
            I => \N__21579\
        );

    \I__3508\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21569\
        );

    \I__3507\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21569\
        );

    \I__3506\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21569\
        );

    \I__3505\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21569\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__21569\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\
        );

    \I__3503\ : InMux
    port map (
            O => \N__21566\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__21563\,
            I => \N__21559\
        );

    \I__3501\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21551\
        );

    \I__3500\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21551\
        );

    \I__3499\ : InMux
    port map (
            O => \N__21558\,
            I => \N__21551\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__21551\,
            I => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\
        );

    \I__3497\ : InMux
    port map (
            O => \N__21548\,
            I => \bfn_6_11_0_\
        );

    \I__3496\ : InMux
    port map (
            O => \N__21545\,
            I => \b2v_inst11.CO2\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__21542\,
            I => \N__21539\
        );

    \I__3494\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21533\
        );

    \I__3493\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21533\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__21533\,
            I => \b2v_inst11.CO2_THRU_CO\
        );

    \I__3491\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21526\
        );

    \I__3490\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21523\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__21526\,
            I => \N__21518\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__21523\,
            I => \N__21518\
        );

    \I__3487\ : Span4Mux_v
    port map (
            O => \N__21518\,
            I => \N__21515\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__21515\,
            I => \b2v_inst11.mult1_un131_sum\
        );

    \I__3485\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21509\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__21509\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_14\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__21506\,
            I => \N__21503\
        );

    \I__3482\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21500\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__21500\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_5\
        );

    \I__3480\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21493\
        );

    \I__3479\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21490\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__21493\,
            I => \N__21487\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21484\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__21487\,
            I => \N__21481\
        );

    \I__3475\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21478\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__21481\,
            I => \b2v_inst11.mult1_un103_sum\
        );

    \I__3473\ : Odrv4
    port map (
            O => \N__21478\,
            I => \b2v_inst11.mult1_un103_sum\
        );

    \I__3472\ : InMux
    port map (
            O => \N__21473\,
            I => \b2v_inst11.un1_dutycycle_53_cry_5\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__3470\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__21464\,
            I => \N__21461\
        );

    \I__3468\ : Span4Mux_v
    port map (
            O => \N__21461\,
            I => \N__21458\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__21458\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_10\
        );

    \I__3466\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21451\
        );

    \I__3465\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21448\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__21451\,
            I => \N__21445\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__21448\,
            I => \N__21440\
        );

    \I__3462\ : Span4Mux_s1_h
    port map (
            O => \N__21445\,
            I => \N__21440\
        );

    \I__3461\ : Span4Mux_h
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__21437\,
            I => \b2v_inst11.mult1_un96_sum\
        );

    \I__3459\ : InMux
    port map (
            O => \N__21434\,
            I => \b2v_inst11.un1_dutycycle_53_cry_6\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__21431\,
            I => \N__21428\
        );

    \I__3457\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__21422\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_11\
        );

    \I__3454\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21415\
        );

    \I__3453\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21412\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__21415\,
            I => \N__21409\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__21412\,
            I => \N__21404\
        );

    \I__3450\ : Span4Mux_s1_h
    port map (
            O => \N__21409\,
            I => \N__21404\
        );

    \I__3449\ : Span4Mux_h
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__3448\ : Odrv4
    port map (
            O => \N__21401\,
            I => \b2v_inst11.mult1_un89_sum\
        );

    \I__3447\ : InMux
    port map (
            O => \N__21398\,
            I => \bfn_6_10_0_\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__3445\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__21389\,
            I => \N__21386\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__21386\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_12\
        );

    \I__3442\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21376\
        );

    \I__3440\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21373\
        );

    \I__3439\ : Span4Mux_h
    port map (
            O => \N__21376\,
            I => \N__21370\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__21373\,
            I => \N__21367\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__21370\,
            I => \b2v_inst11.mult1_un82_sum\
        );

    \I__3436\ : Odrv12
    port map (
            O => \N__21367\,
            I => \b2v_inst11.mult1_un82_sum\
        );

    \I__3435\ : InMux
    port map (
            O => \N__21362\,
            I => \b2v_inst11.un1_dutycycle_53_cry_8\
        );

    \I__3434\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__3432\ : Span4Mux_v
    port map (
            O => \N__21353\,
            I => \N__21350\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__21350\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_13\
        );

    \I__3430\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21343\
        );

    \I__3429\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21340\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__21343\,
            I => \N__21337\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__21340\,
            I => \N__21334\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__21337\,
            I => \b2v_inst11.mult1_un75_sum\
        );

    \I__3425\ : Odrv12
    port map (
            O => \N__21334\,
            I => \b2v_inst11.mult1_un75_sum\
        );

    \I__3424\ : InMux
    port map (
            O => \N__21329\,
            I => \b2v_inst11.un1_dutycycle_53_cry_9\
        );

    \I__3423\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21323\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21320\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__21320\,
            I => \N__21317\
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__21317\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_14\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__21314\,
            I => \N__21310\
        );

    \I__3418\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21307\
        );

    \I__3417\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21304\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21301\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21298\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__21301\,
            I => \N__21295\
        );

    \I__3413\ : Span12Mux_s5_h
    port map (
            O => \N__21298\,
            I => \N__21292\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__21295\,
            I => \b2v_inst11.mult1_un68_sum\
        );

    \I__3411\ : Odrv12
    port map (
            O => \N__21292\,
            I => \b2v_inst11.mult1_un68_sum\
        );

    \I__3410\ : InMux
    port map (
            O => \N__21287\,
            I => \b2v_inst11.un1_dutycycle_53_cry_10\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__21284\,
            I => \N__21281\
        );

    \I__3408\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21278\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__21278\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_15\
        );

    \I__3406\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21271\
        );

    \I__3405\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21268\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__21271\,
            I => \N__21265\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21262\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__21265\,
            I => \N__21259\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__21262\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__21259\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__3399\ : InMux
    port map (
            O => \N__21254\,
            I => \b2v_inst11.un1_dutycycle_53_cry_11\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__3397\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__21245\,
            I => \N__21242\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__21239\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_13\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__3392\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21229\
        );

    \I__3391\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21223\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21220\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__21223\,
            I => \N__21217\
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__21220\,
            I => \b2v_inst11.mult1_un54_sum\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__21217\,
            I => \b2v_inst11.mult1_un54_sum\
        );

    \I__3385\ : InMux
    port map (
            O => \N__21212\,
            I => \b2v_inst11.un1_dutycycle_53_cry_12\
        );

    \I__3384\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21206\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__21206\,
            I => \b2v_inst11.d_i3_mux\
        );

    \I__3382\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__21200\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_0\
        );

    \I__3380\ : InMux
    port map (
            O => \N__21197\,
            I => \b2v_inst11.un1_dutycycle_53_cry_0\
        );

    \I__3379\ : InMux
    port map (
            O => \N__21194\,
            I => \b2v_inst11.un1_dutycycle_53_cry_1\
        );

    \I__3378\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__21188\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_2\
        );

    \I__3376\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21181\
        );

    \I__3375\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21178\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__21181\,
            I => \N__21175\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__21178\,
            I => \N__21172\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__21175\,
            I => \N__21167\
        );

    \I__3371\ : Span4Mux_v
    port map (
            O => \N__21172\,
            I => \N__21167\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__21167\,
            I => \b2v_inst11.mult1_un124_sum\
        );

    \I__3369\ : InMux
    port map (
            O => \N__21164\,
            I => \b2v_inst11.un1_dutycycle_53_cry_2\
        );

    \I__3368\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21157\
        );

    \I__3367\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21154\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__21157\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_7\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__21154\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_7\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__3363\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__21143\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_5\
        );

    \I__3361\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21136\
        );

    \I__3360\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21133\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__21136\,
            I => \N__21130\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__21133\,
            I => \N__21125\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__21130\,
            I => \N__21125\
        );

    \I__3356\ : Span4Mux_v
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__21122\,
            I => \b2v_inst11.mult1_un117_sum\
        );

    \I__3354\ : InMux
    port map (
            O => \N__21119\,
            I => \b2v_inst11.un1_dutycycle_53_cry_3\
        );

    \I__3353\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__21113\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_7\
        );

    \I__3351\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21106\
        );

    \I__3350\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21103\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__21106\,
            I => \N__21100\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__21103\,
            I => \N__21097\
        );

    \I__3347\ : Span12Mux_s5_h
    port map (
            O => \N__21100\,
            I => \N__21094\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__21097\,
            I => \b2v_inst11.mult1_un110_sum\
        );

    \I__3345\ : Odrv12
    port map (
            O => \N__21094\,
            I => \b2v_inst11.mult1_un110_sum\
        );

    \I__3344\ : InMux
    port map (
            O => \N__21089\,
            I => \b2v_inst11.un1_dutycycle_53_cry_4\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__21086\,
            I => \b2v_inst11.dutycycleZ0Z_7_cascade_\
        );

    \I__3342\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__21080\,
            I => \b2v_inst11.dutycycle_RNI_8Z0Z_7\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__21077\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_4_cascade_\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__21074\,
            I => \b2v_inst11.un1_dutycycle_53_axb_8_cascade_\
        );

    \I__3338\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21068\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__21068\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_11\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__21065\,
            I => \b2v_inst11.un1_dutycycle_53_axb_3_1_0_cascade_\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__21062\,
            I => \b2v_inst11.un1_dutycycle_53_axb_3_cascade_\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__21059\,
            I => \b2v_inst11.un1_i3_mux_cascade_\
        );

    \I__3333\ : InMux
    port map (
            O => \N__21056\,
            I => \N__21050\
        );

    \I__3332\ : InMux
    port map (
            O => \N__21055\,
            I => \N__21050\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__21050\,
            I => \b2v_inst11.dutycycleZ1Z_8\
        );

    \I__3330\ : InMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__21044\,
            I => \b2v_inst11.un1_dutycycle_53_3_0_tz\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__21041\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_3_cascade_\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__21038\,
            I => \b2v_inst11.N_26_i_1_cascade_\
        );

    \I__3326\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21032\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__21029\,
            I => \b2v_inst11.un1_dutycycle_53_axb_9_1\
        );

    \I__3323\ : InMux
    port map (
            O => \N__21026\,
            I => \N__21020\
        );

    \I__3322\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21020\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__21020\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__21017\,
            I => \N__21013\
        );

    \I__3319\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21008\
        );

    \I__3318\ : InMux
    port map (
            O => \N__21013\,
            I => \N__21008\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__21008\,
            I => \b2v_inst11.dutycycleZ1Z_4\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__21005\,
            I => \N__21001\
        );

    \I__3315\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20998\
        );

    \I__3314\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20995\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__20998\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__20995\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__3311\ : InMux
    port map (
            O => \N__20990\,
            I => \b2v_inst20.counter_1_cry_26\
        );

    \I__3310\ : InMux
    port map (
            O => \N__20987\,
            I => \b2v_inst20.counter_1_cry_27\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20984\,
            I => \b2v_inst20.counter_1_cry_28\
        );

    \I__3308\ : InMux
    port map (
            O => \N__20981\,
            I => \b2v_inst20.counter_1_cry_29\
        );

    \I__3307\ : InMux
    port map (
            O => \N__20978\,
            I => \b2v_inst20.counter_1_cry_30\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__3305\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20966\
        );

    \I__3304\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20966\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__20966\,
            I => \b2v_inst20.counterZ0Z_28\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__3301\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20954\
        );

    \I__3300\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20954\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__20954\,
            I => \b2v_inst20.counterZ0Z_29\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__20951\,
            I => \N__20947\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__20950\,
            I => \N__20944\
        );

    \I__3296\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20939\
        );

    \I__3295\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20939\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__20939\,
            I => \b2v_inst20.counterZ0Z_30\
        );

    \I__3293\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20930\
        );

    \I__3292\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20930\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__20930\,
            I => \b2v_inst20.counterZ0Z_31\
        );

    \I__3290\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__20924\,
            I => \b2v_inst20.un4_counter_7_and\
        );

    \I__3288\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__20918\,
            I => \b2v_inst11.un1_dutycycle_53_9_1_1\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__20915\,
            I => \b2v_inst11.dutycycleZ1Z_5_cascade_\
        );

    \I__3285\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20908\
        );

    \I__3284\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20905\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__20908\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__20905\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__3281\ : InMux
    port map (
            O => \N__20900\,
            I => \b2v_inst20.counter_1_cry_18\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__20897\,
            I => \N__20893\
        );

    \I__3279\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__3278\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20887\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__20890\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__20887\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__3275\ : InMux
    port map (
            O => \N__20882\,
            I => \b2v_inst20.counter_1_cry_19\
        );

    \I__3274\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20875\
        );

    \I__3273\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20872\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__20875\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__20872\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__3270\ : InMux
    port map (
            O => \N__20867\,
            I => \b2v_inst20.counter_1_cry_20\
        );

    \I__3269\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20860\
        );

    \I__3268\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20857\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__20860\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__20857\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__3265\ : InMux
    port map (
            O => \N__20852\,
            I => \b2v_inst20.counter_1_cry_21\
        );

    \I__3264\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20845\
        );

    \I__3263\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20842\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__20845\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__20842\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__3260\ : InMux
    port map (
            O => \N__20837\,
            I => \b2v_inst20.counter_1_cry_22\
        );

    \I__3259\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20830\
        );

    \I__3258\ : InMux
    port map (
            O => \N__20833\,
            I => \N__20827\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__20830\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__20827\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__3255\ : InMux
    port map (
            O => \N__20822\,
            I => \b2v_inst20.counter_1_cry_23\
        );

    \I__3254\ : InMux
    port map (
            O => \N__20819\,
            I => \N__20815\
        );

    \I__3253\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20812\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__20815\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__20812\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__3250\ : InMux
    port map (
            O => \N__20807\,
            I => \bfn_6_5_0_\
        );

    \I__3249\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20800\
        );

    \I__3248\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20797\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__20800\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__20797\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__3245\ : InMux
    port map (
            O => \N__20792\,
            I => \b2v_inst20.counter_1_cry_25\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__20789\,
            I => \N__20785\
        );

    \I__3243\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20782\
        );

    \I__3242\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20779\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__20782\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__20779\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__3239\ : InMux
    port map (
            O => \N__20774\,
            I => \b2v_inst20.counter_1_cry_9\
        );

    \I__3238\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20767\
        );

    \I__3237\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20764\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__20767\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__20764\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__3234\ : InMux
    port map (
            O => \N__20759\,
            I => \b2v_inst20.counter_1_cry_10\
        );

    \I__3233\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20752\
        );

    \I__3232\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20749\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__20752\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__20749\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__3229\ : InMux
    port map (
            O => \N__20744\,
            I => \b2v_inst20.counter_1_cry_11\
        );

    \I__3228\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20737\
        );

    \I__3227\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20734\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__20737\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__20734\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__3224\ : InMux
    port map (
            O => \N__20729\,
            I => \b2v_inst20.counter_1_cry_12\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__20726\,
            I => \N__20722\
        );

    \I__3222\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20719\
        );

    \I__3221\ : InMux
    port map (
            O => \N__20722\,
            I => \N__20716\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__20719\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__20716\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__3218\ : InMux
    port map (
            O => \N__20711\,
            I => \b2v_inst20.counter_1_cry_13\
        );

    \I__3217\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20704\
        );

    \I__3216\ : InMux
    port map (
            O => \N__20707\,
            I => \N__20701\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__20704\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__20701\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__3213\ : InMux
    port map (
            O => \N__20696\,
            I => \b2v_inst20.counter_1_cry_14\
        );

    \I__3212\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20689\
        );

    \I__3211\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20686\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__20689\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__20686\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__3208\ : InMux
    port map (
            O => \N__20681\,
            I => \b2v_inst20.counter_1_cry_15\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__20678\,
            I => \N__20674\
        );

    \I__3206\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20671\
        );

    \I__3205\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20668\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__20671\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__20668\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__3202\ : InMux
    port map (
            O => \N__20663\,
            I => \bfn_6_4_0_\
        );

    \I__3201\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20656\
        );

    \I__3200\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20653\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__20656\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__20653\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__3197\ : InMux
    port map (
            O => \N__20648\,
            I => \b2v_inst20.counter_1_cry_17\
        );

    \I__3196\ : InMux
    port map (
            O => \N__20645\,
            I => \b2v_inst20.counter_1_cry_1\
        );

    \I__3195\ : InMux
    port map (
            O => \N__20642\,
            I => \b2v_inst20.counter_1_cry_2\
        );

    \I__3194\ : InMux
    port map (
            O => \N__20639\,
            I => \b2v_inst20.counter_1_cry_3\
        );

    \I__3193\ : InMux
    port map (
            O => \N__20636\,
            I => \b2v_inst20.counter_1_cry_4\
        );

    \I__3192\ : InMux
    port map (
            O => \N__20633\,
            I => \b2v_inst20.counter_1_cry_5\
        );

    \I__3191\ : InMux
    port map (
            O => \N__20630\,
            I => \b2v_inst20.counter_1_cry_6\
        );

    \I__3190\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20623\
        );

    \I__3189\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20620\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__20623\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__20620\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__3186\ : InMux
    port map (
            O => \N__20615\,
            I => \b2v_inst20.counter_1_cry_7\
        );

    \I__3185\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20608\
        );

    \I__3184\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20605\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__20608\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__20605\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__3181\ : InMux
    port map (
            O => \N__20600\,
            I => \bfn_6_3_0_\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__20597\,
            I => \N__20594\
        );

    \I__3179\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__20591\,
            I => \b2v_inst11.mult1_un159_sum_cry_2_s\
        );

    \I__3177\ : InMux
    port map (
            O => \N__20588\,
            I => \b2v_inst11.mult1_un159_sum_cry_1\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__3175\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20579\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__20579\,
            I => \b2v_inst11.mult1_un159_sum_cry_3_s\
        );

    \I__3173\ : InMux
    port map (
            O => \N__20576\,
            I => \b2v_inst11.mult1_un159_sum_cry_2\
        );

    \I__3172\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20570\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__20570\,
            I => \b2v_inst11.mult1_un159_sum_cry_4_s\
        );

    \I__3170\ : InMux
    port map (
            O => \N__20567\,
            I => \b2v_inst11.mult1_un159_sum_cry_3\
        );

    \I__3169\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20561\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__20561\,
            I => \b2v_inst11.mult1_un159_sum_cry_5_s\
        );

    \I__3167\ : InMux
    port map (
            O => \N__20558\,
            I => \b2v_inst11.mult1_un159_sum_cry_4\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__3165\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__20549\,
            I => \b2v_inst11.mult1_un166_sum_axb_6\
        );

    \I__3163\ : InMux
    port map (
            O => \N__20546\,
            I => \b2v_inst11.mult1_un159_sum_cry_5\
        );

    \I__3162\ : InMux
    port map (
            O => \N__20543\,
            I => \b2v_inst11.mult1_un159_sum_cry_6\
        );

    \I__3161\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20536\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__20539\,
            I => \N__20532\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20527\
        );

    \I__3158\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20524\
        );

    \I__3157\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20517\
        );

    \I__3156\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20517\
        );

    \I__3155\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20517\
        );

    \I__3154\ : Odrv12
    port map (
            O => \N__20527\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__20524\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__20517\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__20510\,
            I => \N__20507\
        );

    \I__3150\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20504\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20501\
        );

    \I__3148\ : Odrv4
    port map (
            O => \N__20501\,
            I => \b2v_inst11.mult1_un124_sum_i_0_8\
        );

    \I__3147\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__20495\,
            I => \b2v_inst11.mult1_un159_sum_i\
        );

    \I__3145\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20489\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20486\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__20486\,
            I => \b2v_inst11.mult1_un117_sum_i\
        );

    \I__3142\ : InMux
    port map (
            O => \N__20483\,
            I => \b2v_inst11.mult1_un124_sum_cry_2\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__20480\,
            I => \N__20477\
        );

    \I__3140\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20474\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__20474\,
            I => \b2v_inst11.mult1_un117_sum_cry_3_s\
        );

    \I__3138\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__20468\,
            I => \b2v_inst11.mult1_un124_sum_cry_4_s\
        );

    \I__3136\ : InMux
    port map (
            O => \N__20465\,
            I => \b2v_inst11.mult1_un124_sum_cry_3\
        );

    \I__3135\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__20459\,
            I => \b2v_inst11.mult1_un117_sum_cry_4_s\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__20456\,
            I => \N__20453\
        );

    \I__3132\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20450\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__20450\,
            I => \b2v_inst11.mult1_un124_sum_cry_5_s\
        );

    \I__3130\ : InMux
    port map (
            O => \N__20447\,
            I => \b2v_inst11.mult1_un124_sum_cry_4\
        );

    \I__3129\ : InMux
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__20441\,
            I => \N__20437\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__20440\,
            I => \N__20433\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__20437\,
            I => \N__20429\
        );

    \I__3125\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20424\
        );

    \I__3124\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20424\
        );

    \I__3123\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20421\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__20429\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__20424\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__20421\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__3118\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__20408\,
            I => \b2v_inst11.mult1_un117_sum_cry_5_s\
        );

    \I__3116\ : InMux
    port map (
            O => \N__20405\,
            I => \b2v_inst11.mult1_un124_sum_cry_5\
        );

    \I__3115\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20399\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__20399\,
            I => \b2v_inst11.mult1_un117_sum_cry_6_s\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20392\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__20395\,
            I => \N__20388\
        );

    \I__3111\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20381\
        );

    \I__3110\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20381\
        );

    \I__3109\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20381\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__20381\,
            I => \b2v_inst11.mult1_un117_sum_i_0_8\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__3106\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20372\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__20372\,
            I => \b2v_inst11.mult1_un131_sum_axb_8\
        );

    \I__3104\ : InMux
    port map (
            O => \N__20369\,
            I => \b2v_inst11.mult1_un124_sum_cry_6\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__3102\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__20360\,
            I => \b2v_inst11.mult1_un124_sum_axb_8\
        );

    \I__3100\ : InMux
    port map (
            O => \N__20357\,
            I => \b2v_inst11.mult1_un124_sum_cry_7\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__20354\,
            I => \b2v_inst11.mult1_un124_sum_s_8_cascade_\
        );

    \I__3098\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20347\
        );

    \I__3097\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20344\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__20347\,
            I => \b2v_inst11.mult1_un124_sum_cry_6_s\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__20344\,
            I => \b2v_inst11.mult1_un124_sum_cry_6_s\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__3093\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__20333\,
            I => \b2v_inst11.mult1_un131_sum_axb_7_l_fx\
        );

    \I__3091\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20324\
        );

    \I__3089\ : Sp12to4
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__3088\ : Odrv12
    port map (
            O => \N__20321\,
            I => \b2v_inst11.g3_0\
        );

    \I__3087\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__20315\,
            I => \b2v_inst11.mult1_un124_sum_i\
        );

    \I__3085\ : InMux
    port map (
            O => \N__20312\,
            I => \b2v_inst11.mult1_un131_sum_cry_2\
        );

    \I__3084\ : InMux
    port map (
            O => \N__20309\,
            I => \b2v_inst11.mult1_un131_sum_cry_3\
        );

    \I__3083\ : InMux
    port map (
            O => \N__20306\,
            I => \b2v_inst11.mult1_un131_sum_cry_4\
        );

    \I__3082\ : InMux
    port map (
            O => \N__20303\,
            I => \b2v_inst11.mult1_un131_sum_cry_5\
        );

    \I__3081\ : InMux
    port map (
            O => \N__20300\,
            I => \b2v_inst11.mult1_un131_sum_cry_6\
        );

    \I__3080\ : InMux
    port map (
            O => \N__20297\,
            I => \b2v_inst11.mult1_un131_sum_cry_7\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__20294\,
            I => \b2v_inst11.mult1_un131_sum_s_8_cascade_\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__3077\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__20285\,
            I => \b2v_inst11.mult1_un124_sum_i_8\
        );

    \I__3075\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__20279\,
            I => \b2v_inst11.un85_clk_100khz_2\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__3072\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20270\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__20270\,
            I => \b2v_inst11.un85_clk_100khz_1\
        );

    \I__3070\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20264\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__20264\,
            I => \N__20261\
        );

    \I__3068\ : Odrv12
    port map (
            O => \N__20261\,
            I => \b2v_inst11.mult1_un96_sum_i\
        );

    \I__3067\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__20255\,
            I => \b2v_inst11.mult1_un131_sum_i_8\
        );

    \I__3065\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__20249\,
            I => \b2v_inst11.un85_clk_100khz_3\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__20246\,
            I => \N__20242\
        );

    \I__3062\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20235\
        );

    \I__3061\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20235\
        );

    \I__3060\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20232\
        );

    \I__3059\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20229\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20226\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__20232\,
            I => \N__20222\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__20229\,
            I => \N__20219\
        );

    \I__3055\ : Span4Mux_h
    port map (
            O => \N__20226\,
            I => \N__20216\
        );

    \I__3054\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20213\
        );

    \I__3053\ : Span4Mux_h
    port map (
            O => \N__20222\,
            I => \N__20210\
        );

    \I__3052\ : Odrv12
    port map (
            O => \N__20219\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__20216\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__20213\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__20210\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__3048\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20198\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__20198\,
            I => \b2v_inst11.mult1_un103_sum_i_8\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__3045\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__20189\,
            I => \b2v_inst11.mult1_un40_sum_i_5\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__20186\,
            I => \b2v_inst11.mult1_un40_sum_i_5_cascade_\
        );

    \I__3042\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20179\
        );

    \I__3041\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20176\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__20179\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__20176\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__3038\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20166\
        );

    \I__3037\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20163\
        );

    \I__3036\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20160\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__20166\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__20163\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__20160\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__3031\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__20147\,
            I => \b2v_inst11.un1_dutycycle_53_i_29\
        );

    \I__3029\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__20138\,
            I => \N__20135\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__20135\,
            I => \N__20131\
        );

    \I__3025\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20128\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__20131\,
            I => \b2v_inst16.count_rst\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__20128\,
            I => \b2v_inst16.count_rst\
        );

    \I__3022\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20120\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__3020\ : Span4Mux_h
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__3019\ : Span4Mux_v
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__20111\,
            I => \b2v_inst16.count_4_10\
        );

    \I__3017\ : CEMux
    port map (
            O => \N__20108\,
            I => \N__20100\
        );

    \I__3016\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20097\
        );

    \I__3015\ : CEMux
    port map (
            O => \N__20106\,
            I => \N__20090\
        );

    \I__3014\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20080\
        );

    \I__3013\ : CEMux
    port map (
            O => \N__20104\,
            I => \N__20080\
        );

    \I__3012\ : CEMux
    port map (
            O => \N__20103\,
            I => \N__20072\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__20100\,
            I => \N__20069\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__20097\,
            I => \N__20066\
        );

    \I__3009\ : CEMux
    port map (
            O => \N__20096\,
            I => \N__20063\
        );

    \I__3008\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20056\
        );

    \I__3007\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20056\
        );

    \I__3006\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20056\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__20090\,
            I => \N__20053\
        );

    \I__3004\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20050\
        );

    \I__3003\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20045\
        );

    \I__3002\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20045\
        );

    \I__3001\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20040\
        );

    \I__3000\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20040\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__20080\,
            I => \N__20033\
        );

    \I__2998\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20022\
        );

    \I__2997\ : CEMux
    port map (
            O => \N__20078\,
            I => \N__20022\
        );

    \I__2996\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20022\
        );

    \I__2995\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20022\
        );

    \I__2994\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20022\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__20072\,
            I => \N__20019\
        );

    \I__2992\ : Span4Mux_s1_v
    port map (
            O => \N__20069\,
            I => \N__20016\
        );

    \I__2991\ : Span4Mux_v
    port map (
            O => \N__20066\,
            I => \N__20013\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__20063\,
            I => \N__20008\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N__20008\
        );

    \I__2988\ : Span4Mux_s1_v
    port map (
            O => \N__20053\,
            I => \N__20003\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__20050\,
            I => \N__20003\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__20045\,
            I => \N__20000\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__19997\
        );

    \I__2984\ : InMux
    port map (
            O => \N__20039\,
            I => \N__19988\
        );

    \I__2983\ : CEMux
    port map (
            O => \N__20038\,
            I => \N__19988\
        );

    \I__2982\ : InMux
    port map (
            O => \N__20037\,
            I => \N__19988\
        );

    \I__2981\ : InMux
    port map (
            O => \N__20036\,
            I => \N__19988\
        );

    \I__2980\ : Span4Mux_s3_h
    port map (
            O => \N__20033\,
            I => \N__19985\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__19982\
        );

    \I__2978\ : Span4Mux_v
    port map (
            O => \N__20019\,
            I => \N__19965\
        );

    \I__2977\ : Span4Mux_s1_h
    port map (
            O => \N__20016\,
            I => \N__19965\
        );

    \I__2976\ : Span4Mux_v
    port map (
            O => \N__20013\,
            I => \N__19965\
        );

    \I__2975\ : Span4Mux_s1_v
    port map (
            O => \N__20008\,
            I => \N__19965\
        );

    \I__2974\ : Span4Mux_v
    port map (
            O => \N__20003\,
            I => \N__19965\
        );

    \I__2973\ : Span4Mux_s1_v
    port map (
            O => \N__20000\,
            I => \N__19965\
        );

    \I__2972\ : Span4Mux_s1_h
    port map (
            O => \N__19997\,
            I => \N__19965\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19965\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__19985\,
            I => \b2v_inst16.count_en\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__19982\,
            I => \b2v_inst16.count_en\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__19965\,
            I => \b2v_inst16.count_en\
        );

    \I__2967\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__19955\,
            I => \N__19951\
        );

    \I__2965\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19948\
        );

    \I__2964\ : Sp12to4
    port map (
            O => \N__19951\,
            I => \N__19943\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19943\
        );

    \I__2962\ : Span12Mux_s9_v
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__19940\,
            I => \b2v_inst16.countZ0Z_10\
        );

    \I__2960\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__2958\ : Span4Mux_s3_v
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__19928\,
            I => \b2v_inst11.mult1_un110_sum_i\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__2955\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__19919\,
            I => \b2v_inst11.mult1_un117_sum_i_8\
        );

    \I__2953\ : IoInMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__2951\ : Odrv12
    port map (
            O => \N__19910\,
            I => vccst_en
        );

    \I__2950\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__19904\,
            I => \b2v_inst11.un85_clk_100khz_4\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__2947\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__19895\,
            I => \b2v_inst11.mult1_un47_sum_cry_4_s\
        );

    \I__2945\ : InMux
    port map (
            O => \N__19892\,
            I => \b2v_inst11.mult1_un47_sum_cry_3\
        );

    \I__2944\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__19886\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_s\
        );

    \I__2942\ : InMux
    port map (
            O => \N__19883\,
            I => \b2v_inst11.mult1_un47_sum_cry_4\
        );

    \I__2941\ : InMux
    port map (
            O => \N__19880\,
            I => \b2v_inst11.mult1_un47_sum_cry_5\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__2939\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__19871\,
            I => \b2v_inst11.mult1_un47_sum_l_fx_6\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__2936\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__19862\,
            I => \b2v_inst11.mult1_un47_sum_i\
        );

    \I__2934\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__19853\,
            I => \b2v_inst11.un1_dutycycle_53_axb_12\
        );

    \I__2931\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19842\
        );

    \I__2929\ : InMux
    port map (
            O => \N__19846\,
            I => \N__19835\
        );

    \I__2928\ : InMux
    port map (
            O => \N__19845\,
            I => \N__19835\
        );

    \I__2927\ : Span4Mux_h
    port map (
            O => \N__19842\,
            I => \N__19832\
        );

    \I__2926\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19827\
        );

    \I__2925\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19827\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19824\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__19832\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__19827\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__19824\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__19817\,
            I => \N__19813\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__19816\,
            I => \N__19808\
        );

    \I__2918\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19805\
        );

    \I__2917\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19798\
        );

    \I__2916\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19798\
        );

    \I__2915\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19798\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__19805\,
            I => \N__19795\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__19798\,
            I => \N__19792\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__19795\,
            I => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__19792\,
            I => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2910\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__19784\,
            I => \N__19780\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__19783\,
            I => \N__19775\
        );

    \I__2907\ : Span4Mux_v
    port map (
            O => \N__19780\,
            I => \N__19772\
        );

    \I__2906\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19767\
        );

    \I__2905\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19767\
        );

    \I__2904\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19764\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__19772\,
            I => \N__19759\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__19767\,
            I => \N__19759\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__19764\,
            I => \b2v_inst11.count_RNIZ0Z_8\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__19759\,
            I => \b2v_inst11.count_RNIZ0Z_8\
        );

    \I__2899\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__19742\,
            I => \b2v_inst11.curr_state_4_0\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__2893\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__19733\,
            I => \b2v_inst11.mult1_un47_sum_s_4_sf\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__2890\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__19724\,
            I => \b2v_inst11.mult1_un40_sum_i_l_ofx_4\
        );

    \I__2888\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__19718\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_11\
        );

    \I__2886\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__19709\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_7\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\
        );

    \I__2882\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__19700\,
            I => \b2v_inst11.dutycycle_RNI_8Z0Z_6\
        );

    \I__2880\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19692\
        );

    \I__2879\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19687\
        );

    \I__2878\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19687\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__19692\,
            I => \b2v_inst11.mult1_un47_sum_cry_3_s\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__19687\,
            I => \b2v_inst11.mult1_un47_sum_cry_3_s\
        );

    \I__2875\ : InMux
    port map (
            O => \N__19682\,
            I => \b2v_inst11.mult1_un47_sum_cry_2\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__19679\,
            I => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9_cascade_\
        );

    \I__2873\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19672\
        );

    \I__2872\ : InMux
    port map (
            O => \N__19675\,
            I => \N__19669\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__19672\,
            I => \b2v_inst11.dutycycleZ1Z_9\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__19669\,
            I => \b2v_inst11.dutycycleZ1Z_9\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \b2v_inst11.un1_dutycycle_53_30_a1_0_cascade_\
        );

    \I__2868\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__19658\,
            I => \b2v_inst11.un1_dutycycle_53_44_2\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__19655\,
            I => \b2v_inst11.un1_dutycycle_53_5_1_cascade_\
        );

    \I__2865\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19645\
        );

    \I__2864\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19645\
        );

    \I__2863\ : InMux
    port map (
            O => \N__19650\,
            I => \N__19642\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__19645\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_6\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__19642\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_6\
        );

    \I__2860\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19633\
        );

    \I__2859\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19630\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__19633\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_4\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__19630\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_4\
        );

    \I__2856\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__19622\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_8\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__19619\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_8_cascade_\
        );

    \I__2853\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__19613\,
            I => \b2v_inst11.un1_dutycycle_53_9_1\
        );

    \I__2851\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__19607\,
            I => \b2v_inst11.un1_dutycycle_53_axb_7\
        );

    \I__2849\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__19601\,
            I => \b2v_inst20.un4_counter_6_and\
        );

    \I__2847\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__19595\,
            I => \b2v_inst11.un1_dutycycle_53_39_d_0_0\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__19592\,
            I => \b2v_inst11.dutycycle_RNITSFK3Z0Z_10_cascade_\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__19589\,
            I => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10_cascade_\
        );

    \I__2843\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__19583\,
            I => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__2840\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19571\
        );

    \I__2839\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19571\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__19571\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \b2v_inst11.dutycycleZ0Z_1_cascade_\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__19565\,
            I => \b2v_inst11.dutycycle_RNITSFK3Z0Z_9_cascade_\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__2834\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__19556\,
            I => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9\
        );

    \I__2832\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__19550\,
            I => \b2v_inst20.un4_counter_4_and\
        );

    \I__2830\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__19544\,
            I => \b2v_inst20.un4_counter_5_and\
        );

    \I__2828\ : InMux
    port map (
            O => \N__19541\,
            I => \bfn_5_5_0_\
        );

    \I__2827\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19534\
        );

    \I__2826\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19531\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__19534\,
            I => \b2v_inst11.un1_dutycycle_53_axb_11_1\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__19531\,
            I => \b2v_inst11.un1_dutycycle_53_axb_11_1\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__19526\,
            I => \b2v_inst11.un1_dutycycle_53_39_0_1_0_cascade_\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__19523\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_\
        );

    \I__2821\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19516\
        );

    \I__2820\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19513\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19510\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19507\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__19507\,
            I => \N__19501\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__19504\,
            I => \b2v_inst16.curr_state_2_0\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__19501\,
            I => \b2v_inst16.curr_state_2_0\
        );

    \I__2813\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__19493\,
            I => \b2v_inst20.un4_counter_2_and\
        );

    \I__2811\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19487\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__19487\,
            I => \b2v_inst20.un4_counter_3_and\
        );

    \I__2809\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19476\
        );

    \I__2808\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19476\
        );

    \I__2807\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19471\
        );

    \I__2806\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19471\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N_411\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__19471\,
            I => \N_411\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__19466\,
            I => \b2v_inst200.m6_i_0_cascade_\
        );

    \I__2802\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19458\
        );

    \I__2801\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19455\
        );

    \I__2800\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19452\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__19458\,
            I => \N__19447\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__19455\,
            I => \N__19447\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__19452\,
            I => \N__19442\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__19447\,
            I => \N__19434\
        );

    \I__2795\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19429\
        );

    \I__2794\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19429\
        );

    \I__2793\ : Span12Mux_s5_v
    port map (
            O => \N__19442\,
            I => \N__19426\
        );

    \I__2792\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19423\
        );

    \I__2791\ : InMux
    port map (
            O => \N__19440\,
            I => \N__19418\
        );

    \I__2790\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19418\
        );

    \I__2789\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19413\
        );

    \I__2788\ : InMux
    port map (
            O => \N__19437\,
            I => \N__19413\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__19434\,
            I => \N__19408\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__19429\,
            I => \N__19408\
        );

    \I__2785\ : Odrv12
    port map (
            O => \N__19426\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__19423\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__19418\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__19413\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__19408\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__2780\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__19394\,
            I => \b2v_inst200.curr_state_3_0\
        );

    \I__2778\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__19388\,
            I => \b2v_inst200.curr_stateZ0Z_2\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__19385\,
            I => \b2v_inst200.i4_mux_cascade_\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__19382\,
            I => \b2v_inst200.curr_state_i_2_cascade_\
        );

    \I__2774\ : IoInMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__2772\ : IoSpan4Mux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__2771\ : Span4Mux_s0_h
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__19364\,
            I => hda_sdo_atp
        );

    \I__2768\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19357\
        );

    \I__2767\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__19357\,
            I => \b2v_inst200.N_3031_i\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__19354\,
            I => \b2v_inst200.N_3031_i\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__19349\,
            I => \N__19345\
        );

    \I__2763\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19337\
        );

    \I__2762\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19337\
        );

    \I__2761\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19337\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__19337\,
            I => \b2v_inst200.N_205\
        );

    \I__2759\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19325\
        );

    \I__2758\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19325\
        );

    \I__2757\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19325\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__19325\,
            I => \b2v_inst200.curr_state_i_2\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__19322\,
            I => \b2v_inst200.N_205_cascade_\
        );

    \I__2754\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__19316\,
            I => \b2v_inst200.HDA_SDO_ATP_0\
        );

    \I__2752\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19305\
        );

    \I__2751\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19305\
        );

    \I__2750\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19300\
        );

    \I__2749\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19300\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__19305\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__19300\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__19295\,
            I => \N__19291\
        );

    \I__2745\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19287\
        );

    \I__2744\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19284\
        );

    \I__2743\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19281\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__19287\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__19284\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__19281\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__19274\,
            I => \N__19268\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__19273\,
            I => \N__19265\
        );

    \I__2737\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19258\
        );

    \I__2736\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19258\
        );

    \I__2735\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19258\
        );

    \I__2734\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19255\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__19258\,
            I => \b2v_inst200.N_282\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__19255\,
            I => \b2v_inst200.N_282\
        );

    \I__2731\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__19247\,
            I => \b2v_inst200.curr_state_3_1\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__19244\,
            I => \N__19240\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__19243\,
            I => \N__19236\
        );

    \I__2727\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19229\
        );

    \I__2726\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19229\
        );

    \I__2725\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19229\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__19229\,
            I => \G_2814\
        );

    \I__2723\ : InMux
    port map (
            O => \N__19226\,
            I => \b2v_inst11.mult1_un166_sum_cry_5\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__2721\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__2719\ : Odrv12
    port map (
            O => \N__19214\,
            I => \b2v_inst11.un85_clk_100khz_0\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__19211\,
            I => \b2v_inst200.N_58_cascade_\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__19208\,
            I => \b2v_inst200.curr_stateZ0Z_0_cascade_\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__19205\,
            I => \b2v_inst200.curr_stateZ0Z_1_cascade_\
        );

    \I__2715\ : InMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__19199\,
            I => \b2v_inst200.N_56\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__2712\ : InMux
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__19184\,
            I => gpio_fpga_soc_1
        );

    \I__2708\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__19178\,
            I => \b2v_inst200.m6_i_0\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__19175\,
            I => \N__19170\
        );

    \I__2705\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19166\
        );

    \I__2704\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19161\
        );

    \I__2703\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19161\
        );

    \I__2702\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19158\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__19166\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__19161\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__19158\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__2697\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__19145\,
            I => \b2v_inst11.mult1_un110_sum_cry_5_s\
        );

    \I__2695\ : InMux
    port map (
            O => \N__19142\,
            I => \b2v_inst11.mult1_un117_sum_cry_5\
        );

    \I__2694\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__19136\,
            I => \b2v_inst11.mult1_un110_sum_cry_6_s\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \N__19129\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__19132\,
            I => \N__19125\
        );

    \I__2690\ : InMux
    port map (
            O => \N__19129\,
            I => \N__19118\
        );

    \I__2689\ : InMux
    port map (
            O => \N__19128\,
            I => \N__19118\
        );

    \I__2688\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19118\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__19118\,
            I => \b2v_inst11.mult1_un110_sum_i_0_8\
        );

    \I__2686\ : InMux
    port map (
            O => \N__19115\,
            I => \b2v_inst11.mult1_un117_sum_cry_6\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__2684\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__19106\,
            I => \b2v_inst11.mult1_un117_sum_axb_8\
        );

    \I__2682\ : InMux
    port map (
            O => \N__19103\,
            I => \b2v_inst11.mult1_un117_sum_cry_7\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__19100\,
            I => \b2v_inst11.mult1_un117_sum_s_8_cascade_\
        );

    \I__2680\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__19088\,
            I => \b2v_inst11.mult1_un103_sum_cry_4_s\
        );

    \I__2676\ : InMux
    port map (
            O => \N__19085\,
            I => \b2v_inst11.mult1_un110_sum_cry_4\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__2674\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__19070\,
            I => \b2v_inst11.mult1_un103_sum_cry_5_s\
        );

    \I__2670\ : InMux
    port map (
            O => \N__19067\,
            I => \b2v_inst11.mult1_un110_sum_cry_5\
        );

    \I__2669\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__19055\,
            I => \b2v_inst11.mult1_un103_sum_cry_6_s\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__19052\,
            I => \N__19048\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__19051\,
            I => \N__19044\
        );

    \I__2663\ : InMux
    port map (
            O => \N__19048\,
            I => \N__19037\
        );

    \I__2662\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19037\
        );

    \I__2661\ : InMux
    port map (
            O => \N__19044\,
            I => \N__19037\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__19037\,
            I => \b2v_inst11.mult1_un103_sum_i_0_8\
        );

    \I__2659\ : InMux
    port map (
            O => \N__19034\,
            I => \b2v_inst11.mult1_un110_sum_cry_6\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__2657\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19025\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__19019\,
            I => \b2v_inst11.mult1_un110_sum_axb_8\
        );

    \I__2653\ : InMux
    port map (
            O => \N__19016\,
            I => \b2v_inst11.mult1_un110_sum_cry_7\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__19013\,
            I => \b2v_inst11.mult1_un110_sum_s_8_cascade_\
        );

    \I__2651\ : InMux
    port map (
            O => \N__19010\,
            I => \b2v_inst11.mult1_un117_sum_cry_2\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__2649\ : InMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__19001\,
            I => \b2v_inst11.mult1_un110_sum_cry_3_s\
        );

    \I__2647\ : InMux
    port map (
            O => \N__18998\,
            I => \b2v_inst11.mult1_un117_sum_cry_3\
        );

    \I__2646\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__18992\,
            I => \b2v_inst11.mult1_un110_sum_cry_4_s\
        );

    \I__2644\ : InMux
    port map (
            O => \N__18989\,
            I => \b2v_inst11.mult1_un117_sum_cry_4\
        );

    \I__2643\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__18983\,
            I => \N__18980\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__18980\,
            I => \b2v_inst11.mult1_un68_sum_i_8\
        );

    \I__2640\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__2638\ : Span12Mux_s10_h
    port map (
            O => \N__18971\,
            I => \N__18966\
        );

    \I__2637\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18963\
        );

    \I__2636\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18960\
        );

    \I__2635\ : Odrv12
    port map (
            O => \N__18966\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__18963\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__18960\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__2631\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__18944\,
            I => \b2v_inst11.N_5994_i\
        );

    \I__2628\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18938\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__18935\,
            I => \N__18930\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18927\
        );

    \I__2624\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18924\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__18930\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__18927\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__18924\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__2620\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__18911\,
            I => \b2v_inst11.mult1_un61_sum_i_8\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__2616\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__18902\,
            I => \b2v_inst11.N_5995_i\
        );

    \I__2614\ : InMux
    port map (
            O => \N__18899\,
            I => \bfn_4_13_0_\
        );

    \I__2613\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__18893\,
            I => \b2v_inst11.mult1_un110_sum_i_8\
        );

    \I__2611\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__18881\,
            I => \b2v_inst11.mult1_un103_sum_i\
        );

    \I__2607\ : InMux
    port map (
            O => \N__18878\,
            I => \b2v_inst11.mult1_un110_sum_cry_2\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__2605\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__2603\ : Span4Mux_h
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__18863\,
            I => \b2v_inst11.mult1_un103_sum_cry_3_s\
        );

    \I__2601\ : InMux
    port map (
            O => \N__18860\,
            I => \b2v_inst11.mult1_un110_sum_cry_3\
        );

    \I__2600\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__18851\,
            I => \N__18848\
        );

    \I__2597\ : Span4Mux_v
    port map (
            O => \N__18848\,
            I => \N__18843\
        );

    \I__2596\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18840\
        );

    \I__2595\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18837\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__18843\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__18840\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__18837\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__2591\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__18827\,
            I => \b2v_inst11.N_5986_i\
        );

    \I__2589\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__2586\ : Span4Mux_v
    port map (
            O => \N__18815\,
            I => \N__18810\
        );

    \I__2585\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18807\
        );

    \I__2584\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18804\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__18810\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__18807\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__18804\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__2580\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__18794\,
            I => \b2v_inst11.N_5987_i\
        );

    \I__2578\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__18788\,
            I => \N__18783\
        );

    \I__2576\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18780\
        );

    \I__2575\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18777\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__18783\,
            I => \N__18774\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__18780\,
            I => \N__18771\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18768\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__18774\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__18771\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__18768\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__2567\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__18755\,
            I => \b2v_inst11.N_5988_i\
        );

    \I__2565\ : InMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__18749\,
            I => \N__18744\
        );

    \I__2563\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18741\
        );

    \I__2562\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18738\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__18744\,
            I => \N__18731\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__18741\,
            I => \N__18731\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__18738\,
            I => \N__18731\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__18731\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__18728\,
            I => \N__18725\
        );

    \I__2556\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__18722\,
            I => \b2v_inst11.N_5989_i\
        );

    \I__2554\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__18713\,
            I => \N__18710\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__18710\,
            I => \b2v_inst11.mult1_un96_sum_i_8\
        );

    \I__2550\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__18704\,
            I => \N__18700\
        );

    \I__2548\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18696\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__18700\,
            I => \N__18693\
        );

    \I__2546\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18690\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__18696\,
            I => \N__18687\
        );

    \I__2544\ : Span4Mux_s0_h
    port map (
            O => \N__18693\,
            I => \N__18682\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__18690\,
            I => \N__18682\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__18687\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__18682\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__2539\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__18671\,
            I => \b2v_inst11.N_5990_i\
        );

    \I__2537\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18665\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__18665\,
            I => \N__18662\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__18662\,
            I => \b2v_inst11.mult1_un89_sum_i_8\
        );

    \I__2534\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18655\
        );

    \I__2533\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18652\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__18655\,
            I => \N__18648\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__18652\,
            I => \N__18645\
        );

    \I__2530\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18642\
        );

    \I__2529\ : Span4Mux_s3_v
    port map (
            O => \N__18648\,
            I => \N__18639\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__18645\,
            I => \N__18634\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__18642\,
            I => \N__18634\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__18639\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__18634\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__2523\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__18623\,
            I => \b2v_inst11.N_5991_i\
        );

    \I__2521\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18612\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__18616\,
            I => \N__18609\
        );

    \I__2518\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18606\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__18612\,
            I => \N__18603\
        );

    \I__2516\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18600\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18597\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__18603\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__18600\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__18597\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__2511\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__2509\ : Span4Mux_h
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__18581\,
            I => \b2v_inst11.mult1_un82_sum_i_8\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__2506\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__18572\,
            I => \b2v_inst11.N_5992_i\
        );

    \I__2504\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__18560\,
            I => \b2v_inst11.mult1_un75_sum_i_8\
        );

    \I__2500\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18553\
        );

    \I__2499\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18550\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18547\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18544\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__18547\,
            I => \N__18538\
        );

    \I__2495\ : Span4Mux_s2_v
    port map (
            O => \N__18544\,
            I => \N__18538\
        );

    \I__2494\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18535\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__18538\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__18535\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__2490\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__18524\,
            I => \b2v_inst11.N_5993_i\
        );

    \I__2488\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__18515\,
            I => \b2v_inst11.mult1_un75_sum_i\
        );

    \I__2485\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18505\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__18508\,
            I => \N__18501\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__18505\,
            I => \N__18497\
        );

    \I__2481\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18492\
        );

    \I__2480\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18492\
        );

    \I__2479\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18489\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__18497\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__18492\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__18489\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__2475\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18475\
        );

    \I__2473\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18468\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__18475\,
            I => \N__18465\
        );

    \I__2471\ : InMux
    port map (
            O => \N__18474\,
            I => \N__18462\
        );

    \I__2470\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18455\
        );

    \I__2469\ : InMux
    port map (
            O => \N__18472\,
            I => \N__18455\
        );

    \I__2468\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18455\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__18468\,
            I => \N__18452\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__18465\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__18462\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__18455\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__18452\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__2462\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__18440\,
            I => \b2v_inst11.N_5980_i\
        );

    \I__2460\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__18434\,
            I => \N__18429\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__18433\,
            I => \N__18426\
        );

    \I__2457\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18423\
        );

    \I__2456\ : Span4Mux_v
    port map (
            O => \N__18429\,
            I => \N__18420\
        );

    \I__2455\ : InMux
    port map (
            O => \N__18426\,
            I => \N__18417\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__18423\,
            I => \N__18414\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__18420\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__18417\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__18414\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__2450\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__18404\,
            I => \b2v_inst11.N_5981_i\
        );

    \I__2448\ : InMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__18395\,
            I => \N__18391\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__18394\,
            I => \N__18388\
        );

    \I__2444\ : Span4Mux_h
    port map (
            O => \N__18391\,
            I => \N__18384\
        );

    \I__2443\ : InMux
    port map (
            O => \N__18388\,
            I => \N__18381\
        );

    \I__2442\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18378\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__18384\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__18381\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__18378\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__2437\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__18365\,
            I => \b2v_inst11.N_5982_i\
        );

    \I__2435\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__18359\,
            I => \N__18355\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__18358\,
            I => \N__18351\
        );

    \I__2432\ : Span4Mux_v
    port map (
            O => \N__18355\,
            I => \N__18348\
        );

    \I__2431\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18345\
        );

    \I__2430\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18342\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__18348\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__18345\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__18342\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__2425\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__18329\,
            I => \b2v_inst11.N_5983_i\
        );

    \I__2423\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18323\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__18320\,
            I => \N__18315\
        );

    \I__2420\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18312\
        );

    \I__2419\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18309\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__18315\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__18312\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__18309\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__18302\,
            I => \N__18299\
        );

    \I__2414\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__18296\,
            I => \b2v_inst11.N_5984_i\
        );

    \I__2412\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__18287\,
            I => \N__18282\
        );

    \I__2409\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18279\
        );

    \I__2408\ : InMux
    port map (
            O => \N__18285\,
            I => \N__18276\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__18282\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__18279\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__18276\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__2403\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18263\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__18263\,
            I => \b2v_inst11.N_5985_i\
        );

    \I__2401\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__18254\,
            I => \b2v_inst11.mult1_un61_sum_axb_8\
        );

    \I__2398\ : InMux
    port map (
            O => \N__18251\,
            I => \b2v_inst11.mult1_un54_sum_cry_6\
        );

    \I__2397\ : InMux
    port map (
            O => \N__18248\,
            I => \b2v_inst11.mult1_un54_sum_cry_7\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__18245\,
            I => \N__18240\
        );

    \I__2395\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18237\
        );

    \I__2394\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18232\
        );

    \I__2393\ : InMux
    port map (
            O => \N__18240\,
            I => \N__18232\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__18237\,
            I => \N__18228\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__18232\,
            I => \N__18225\
        );

    \I__2390\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18222\
        );

    \I__2389\ : Span4Mux_s3_h
    port map (
            O => \N__18228\,
            I => \N__18219\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__18225\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__18222\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__18219\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__2384\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__18206\,
            I => \b2v_inst11.mult1_un47_sum_l_fx_3\
        );

    \I__2382\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__18194\,
            I => vpp_ok
        );

    \I__2378\ : IoInMux
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__2376\ : IoSpan4Mux
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__2375\ : Span4Mux_s1_h
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__18179\,
            I => \N__18176\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__18176\,
            I => vddq_en
        );

    \I__2372\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__2370\ : Span4Mux_s3_h
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__18164\,
            I => \b2v_inst11.mult1_un54_sum_i\
        );

    \I__2368\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__18158\,
            I => \N__18154\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__18157\,
            I => \N__18150\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__18154\,
            I => \N__18146\
        );

    \I__2364\ : InMux
    port map (
            O => \N__18153\,
            I => \N__18141\
        );

    \I__2363\ : InMux
    port map (
            O => \N__18150\,
            I => \N__18141\
        );

    \I__2362\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18138\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__18146\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__18141\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__18138\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__2358\ : InMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__2356\ : Span4Mux_s3_h
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__18122\,
            I => \b2v_inst11.mult1_un61_sum_i\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__18119\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_6_cascade_\
        );

    \I__2353\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__18113\,
            I => \b2v_inst11.dutycycle_RNI_9Z0Z_7\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__18110\,
            I => \b2v_inst11.un1_dutycycle_53_46_0_cascade_\
        );

    \I__2350\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__18101\,
            I => \b2v_inst11.un1_dutycycle_53_axb_11_1_0\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__2346\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__18089\,
            I => \b2v_inst11.mult1_un54_sum_cry_3_s\
        );

    \I__2343\ : InMux
    port map (
            O => \N__18086\,
            I => \b2v_inst11.mult1_un54_sum_cry_2\
        );

    \I__2342\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__18077\,
            I => \b2v_inst11.mult1_un54_sum_cry_4_s\
        );

    \I__2339\ : InMux
    port map (
            O => \N__18074\,
            I => \b2v_inst11.mult1_un54_sum_cry_3\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__2337\ : InMux
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__18062\,
            I => \b2v_inst11.mult1_un54_sum_cry_5_s\
        );

    \I__2334\ : InMux
    port map (
            O => \N__18059\,
            I => \b2v_inst11.mult1_un54_sum_cry_4\
        );

    \I__2333\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__18050\,
            I => \b2v_inst11.mult1_un54_sum_cry_6_s\
        );

    \I__2330\ : InMux
    port map (
            O => \N__18047\,
            I => \b2v_inst11.mult1_un54_sum_cry_5\
        );

    \I__2329\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__18041\,
            I => \b2v_inst11.un1_dutycycle_53_55_1_tz\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__18038\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_11_cascade_\
        );

    \I__2326\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__18032\,
            I => \b2v_inst11.un1_dutycycle_53_50_a0_1\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__18029\,
            I => \b2v_inst11.un1_dutycycle_53_50_a0_1_cascade_\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__18026\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_6_cascade_\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__18023\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_12_cascade_\
        );

    \I__2321\ : InMux
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__18017\,
            I => \b2v_inst11.un1_dutycycle_53_4_1\
        );

    \I__2319\ : InMux
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__18011\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_12\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__18008\,
            I => \b2v_inst11.un1_dutycycle_53_4_1_cascade_\
        );

    \I__2316\ : InMux
    port map (
            O => \N__18005\,
            I => \N__17999\
        );

    \I__2315\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17999\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__17999\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_8\
        );

    \I__2313\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__2310\ : Odrv4
    port map (
            O => \N__17987\,
            I => \b2v_inst16.curr_state_2_1\
        );

    \I__2309\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__2307\ : Span4Mux_v
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__17975\,
            I => \b2v_inst16.curr_state_7_0_1\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__17972\,
            I => \b2v_inst11.un1_dutycycle_53_44_0_2_cascade_\
        );

    \I__2304\ : InMux
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__17966\,
            I => \b2v_inst11.un2_count_clk_17_0_a2_1_4\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__17963\,
            I => \b2v_inst11.N_355_cascade_\
        );

    \I__2301\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17954\
        );

    \I__2300\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17954\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__17951\,
            I => \b2v_inst16.count_rst_1\
        );

    \I__2297\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17945\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__17945\,
            I => \b2v_inst16.count_4_12\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__17942\,
            I => \N__17938\
        );

    \I__2294\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17935\
        );

    \I__2293\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17932\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__17935\,
            I => \N__17929\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__17932\,
            I => \b2v_inst16.countZ0Z_13\
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__17929\,
            I => \b2v_inst16.countZ0Z_13\
        );

    \I__2289\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17918\
        );

    \I__2288\ : InMux
    port map (
            O => \N__17923\,
            I => \N__17918\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__17915\,
            I => \b2v_inst16.count_rst_2\
        );

    \I__2285\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__17909\,
            I => \b2v_inst16.count_4_13\
        );

    \I__2283\ : SRMux
    port map (
            O => \N__17906\,
            I => \N__17900\
        );

    \I__2282\ : SRMux
    port map (
            O => \N__17905\,
            I => \N__17896\
        );

    \I__2281\ : SRMux
    port map (
            O => \N__17904\,
            I => \N__17893\
        );

    \I__2280\ : SRMux
    port map (
            O => \N__17903\,
            I => \N__17889\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__17900\,
            I => \N__17885\
        );

    \I__2278\ : SRMux
    port map (
            O => \N__17899\,
            I => \N__17882\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__17896\,
            I => \N__17877\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__17893\,
            I => \N__17877\
        );

    \I__2275\ : SRMux
    port map (
            O => \N__17892\,
            I => \N__17874\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__17889\,
            I => \N__17871\
        );

    \I__2273\ : SRMux
    port map (
            O => \N__17888\,
            I => \N__17868\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__17885\,
            I => \N__17863\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__17882\,
            I => \N__17863\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__17877\,
            I => \N__17860\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__17874\,
            I => \N__17857\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__17871\,
            I => \N__17852\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__17868\,
            I => \N__17852\
        );

    \I__2266\ : Span4Mux_h
    port map (
            O => \N__17863\,
            I => \N__17849\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__17860\,
            I => \b2v_inst16.N_3079_i\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__17857\,
            I => \b2v_inst16.N_3079_i\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__17852\,
            I => \b2v_inst16.N_3079_i\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__17849\,
            I => \b2v_inst16.N_3079_i\
        );

    \I__2261\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__17831\,
            I => \b2v_inst16.count_4_3\
        );

    \I__2257\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__17825\,
            I => \b2v_inst16.count_rst_8\
        );

    \I__2255\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17818\
        );

    \I__2254\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17815\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__17818\,
            I => \N__17811\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__17815\,
            I => \N__17808\
        );

    \I__2251\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17804\
        );

    \I__2250\ : Span4Mux_s3_h
    port map (
            O => \N__17811\,
            I => \N__17801\
        );

    \I__2249\ : Span4Mux_s3_h
    port map (
            O => \N__17808\,
            I => \N__17798\
        );

    \I__2248\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17795\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__17804\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__17801\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__17798\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__17795\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__2243\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17780\
        );

    \I__2242\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17780\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__17780\,
            I => \b2v_inst11.dutycycleZ1Z_7\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__17777\,
            I => \b2v_inst11.dutycycleZ1Z_3_cascade_\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__17774\,
            I => \b2v_inst11.un1_dutycycle_53_axb_7_1_cascade_\
        );

    \I__2238\ : IoInMux
    port map (
            O => \N__17771\,
            I => \N__17768\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__17768\,
            I => \N__17765\
        );

    \I__2236\ : Span4Mux_s3_h
    port map (
            O => \N__17765\,
            I => \N__17762\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__17762\,
            I => \N__17759\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__17759\,
            I => \N__17756\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__17753\,
            I => vpp_en
        );

    \I__2231\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17747\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__17747\,
            I => \b2v_inst16.delayed_vddq_pwrgd_eZ0Z_0\
        );

    \I__2229\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17738\
        );

    \I__2228\ : CEMux
    port map (
            O => \N__17743\,
            I => \N__17738\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__17735\,
            I => \b2v_inst16.delayed_vddq_pwrgd_en\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__17732\,
            I => \N__17718\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__17731\,
            I => \N__17705\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__17730\,
            I => \N__17701\
        );

    \I__2222\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17695\
        );

    \I__2221\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17692\
        );

    \I__2220\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17683\
        );

    \I__2219\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17683\
        );

    \I__2218\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17683\
        );

    \I__2217\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17683\
        );

    \I__2216\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17675\
        );

    \I__2215\ : InMux
    port map (
            O => \N__17722\,
            I => \N__17675\
        );

    \I__2214\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17675\
        );

    \I__2213\ : InMux
    port map (
            O => \N__17718\,
            I => \N__17662\
        );

    \I__2212\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17662\
        );

    \I__2211\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17662\
        );

    \I__2210\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17662\
        );

    \I__2209\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17662\
        );

    \I__2208\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17662\
        );

    \I__2207\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17653\
        );

    \I__2206\ : InMux
    port map (
            O => \N__17711\,
            I => \N__17653\
        );

    \I__2205\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17653\
        );

    \I__2204\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17653\
        );

    \I__2203\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17642\
        );

    \I__2202\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17642\
        );

    \I__2201\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17642\
        );

    \I__2200\ : InMux
    port map (
            O => \N__17701\,
            I => \N__17642\
        );

    \I__2199\ : InMux
    port map (
            O => \N__17700\,
            I => \N__17642\
        );

    \I__2198\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17639\
        );

    \I__2197\ : InMux
    port map (
            O => \N__17698\,
            I => \N__17636\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__17695\,
            I => \N__17633\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17628\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__17683\,
            I => \N__17628\
        );

    \I__2193\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17625\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__17675\,
            I => \N__17620\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__17662\,
            I => \N__17620\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__17653\,
            I => \N__17615\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__17642\,
            I => \N__17615\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__17639\,
            I => \N__17611\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__17636\,
            I => \N__17608\
        );

    \I__2186\ : Span4Mux_s2_v
    port map (
            O => \N__17633\,
            I => \N__17601\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__17628\,
            I => \N__17601\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17601\
        );

    \I__2183\ : Span4Mux_s3_h
    port map (
            O => \N__17620\,
            I => \N__17598\
        );

    \I__2182\ : Span4Mux_s3_h
    port map (
            O => \N__17615\,
            I => \N__17595\
        );

    \I__2181\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17592\
        );

    \I__2180\ : Odrv12
    port map (
            O => \N__17611\,
            I => \b2v_inst16.N_26\
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__17608\,
            I => \b2v_inst16.N_26\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__17601\,
            I => \b2v_inst16.N_26\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__17598\,
            I => \b2v_inst16.N_26\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__17595\,
            I => \b2v_inst16.N_26\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__17592\,
            I => \b2v_inst16.N_26\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__17579\,
            I => \N__17572\
        );

    \I__2173\ : InMux
    port map (
            O => \N__17578\,
            I => \N__17561\
        );

    \I__2172\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17550\
        );

    \I__2171\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17550\
        );

    \I__2170\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17550\
        );

    \I__2169\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17550\
        );

    \I__2168\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17550\
        );

    \I__2167\ : InMux
    port map (
            O => \N__17570\,
            I => \N__17547\
        );

    \I__2166\ : InMux
    port map (
            O => \N__17569\,
            I => \N__17544\
        );

    \I__2165\ : InMux
    port map (
            O => \N__17568\,
            I => \N__17532\
        );

    \I__2164\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17532\
        );

    \I__2163\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17532\
        );

    \I__2162\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17532\
        );

    \I__2161\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17529\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__17561\,
            I => \N__17524\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__17550\,
            I => \N__17524\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__17547\,
            I => \N__17519\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__17544\,
            I => \N__17519\
        );

    \I__2156\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17516\
        );

    \I__2155\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17511\
        );

    \I__2154\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17511\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__17532\,
            I => \N__17508\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__17529\,
            I => \N__17503\
        );

    \I__2151\ : Span4Mux_s0_v
    port map (
            O => \N__17524\,
            I => \N__17503\
        );

    \I__2150\ : Span12Mux_s2_v
    port map (
            O => \N__17519\,
            I => \N__17500\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__17516\,
            I => \b2v_inst16.N_416\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__17511\,
            I => \b2v_inst16.N_416\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__17508\,
            I => \b2v_inst16.N_416\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__17503\,
            I => \b2v_inst16.N_416\
        );

    \I__2145\ : Odrv12
    port map (
            O => \N__17500\,
            I => \b2v_inst16.N_416\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__17489\,
            I => \N__17485\
        );

    \I__2143\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17482\
        );

    \I__2142\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17479\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__17482\,
            I => \N__17476\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__17479\,
            I => \N__17473\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__17476\,
            I => \b2v_inst16.un4_count_1_cry_2_THRU_CO\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__17473\,
            I => \b2v_inst16.un4_count_1_cry_2_THRU_CO\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__17468\,
            I => \b2v_inst16.N_26_cascade_\
        );

    \I__2136\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__17462\,
            I => \N__17459\
        );

    \I__2134\ : Span4Mux_s3_h
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__17456\,
            I => \b2v_inst16.count_4_i_a3_10_0\
        );

    \I__2132\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17449\
        );

    \I__2131\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17446\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__17449\,
            I => \N__17443\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__17446\,
            I => \b2v_inst16.countZ0Z_14\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__17443\,
            I => \b2v_inst16.countZ0Z_14\
        );

    \I__2127\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17432\
        );

    \I__2126\ : InMux
    port map (
            O => \N__17437\,
            I => \N__17432\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__2124\ : Odrv12
    port map (
            O => \N__17429\,
            I => \b2v_inst16.count_rst_3\
        );

    \I__2123\ : InMux
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__17423\,
            I => \b2v_inst16.count_4_14\
        );

    \I__2121\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17416\
        );

    \I__2120\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17413\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__17416\,
            I => \N__17410\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__17413\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__17410\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__2115\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17396\
        );

    \I__2114\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17396\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__17396\,
            I => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\
        );

    \I__2112\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17390\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__17390\,
            I => \b2v_inst11.count_0_15\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__2109\ : InMux
    port map (
            O => \N__17384\,
            I => \N__17378\
        );

    \I__2108\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17378\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__17378\,
            I => \b2v_inst11.count_1_7\
        );

    \I__2106\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__17372\,
            I => \b2v_inst11.count_0_7\
        );

    \I__2104\ : IoInMux
    port map (
            O => \N__17369\,
            I => \N__17366\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__2102\ : Span4Mux_s3_h
    port map (
            O => \N__17363\,
            I => \N__17360\
        );

    \I__2101\ : Sp12to4
    port map (
            O => \N__17360\,
            I => \N__17357\
        );

    \I__2100\ : Odrv12
    port map (
            O => \N__17357\,
            I => \b2v_inst200.count_enZ0\
        );

    \I__2099\ : IoInMux
    port map (
            O => \N__17354\,
            I => \N__17351\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__17351\,
            I => \N__17348\
        );

    \I__2097\ : IoSpan4Mux
    port map (
            O => \N__17348\,
            I => \N__17345\
        );

    \I__2096\ : Span4Mux_s0_h
    port map (
            O => \N__17345\,
            I => \N__17341\
        );

    \I__2095\ : IoInMux
    port map (
            O => \N__17344\,
            I => \N__17338\
        );

    \I__2094\ : Sp12to4
    port map (
            O => \N__17341\,
            I => \N__17334\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__17338\,
            I => \N__17331\
        );

    \I__2092\ : IoInMux
    port map (
            O => \N__17337\,
            I => \N__17328\
        );

    \I__2091\ : Span12Mux_s8_h
    port map (
            O => \N__17334\,
            I => \N__17325\
        );

    \I__2090\ : IoSpan4Mux
    port map (
            O => \N__17331\,
            I => \N__17322\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__17328\,
            I => \N__17319\
        );

    \I__2088\ : Odrv12
    port map (
            O => \N__17325\,
            I => pch_pwrok
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__17322\,
            I => pch_pwrok
        );

    \I__2086\ : Odrv12
    port map (
            O => \N__17319\,
            I => pch_pwrok
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__17312\,
            I => \b2v_inst11.un79_clk_100khzlt6_cascade_\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__17309\,
            I => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__17306\,
            I => \b2v_inst11.un79_clk_100khzlto15_7_cascade_\
        );

    \I__2082\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__17300\,
            I => \b2v_inst11.un79_clk_100khzlto15_3\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \b2v_inst11.count_RNIZ0Z_8_cascade_\
        );

    \I__2079\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17288\
        );

    \I__2078\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17288\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__17288\,
            I => \N__17285\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__17285\,
            I => \b2v_inst11.N_8\
        );

    \I__2075\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17276\
        );

    \I__2074\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17276\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__17276\,
            I => \b2v_inst11.count_1_14\
        );

    \I__2072\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17270\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__17270\,
            I => \b2v_inst11.count_0_14\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2069\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17258\
        );

    \I__2068\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17258\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__17258\,
            I => \b2v_inst11.count_1_6\
        );

    \I__2066\ : InMux
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__17252\,
            I => \b2v_inst11.count_0_6\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__17249\,
            I => \N__17246\
        );

    \I__2063\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17240\
        );

    \I__2062\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17240\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__17240\,
            I => \b2v_inst11.count_1_3\
        );

    \I__2060\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17234\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__17234\,
            I => \b2v_inst11.count_0_3\
        );

    \I__2058\ : InMux
    port map (
            O => \N__17231\,
            I => \N__17225\
        );

    \I__2057\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17225\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__17222\,
            I => \b2v_inst11.count_1_13\
        );

    \I__2054\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__17216\,
            I => \b2v_inst11.count_0_13\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__17213\,
            I => \N__17210\
        );

    \I__2051\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17204\
        );

    \I__2050\ : InMux
    port map (
            O => \N__17209\,
            I => \N__17204\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__17204\,
            I => \b2v_inst11.count_1_4\
        );

    \I__2048\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__17198\,
            I => \b2v_inst11.count_0_4\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__2045\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17186\
        );

    \I__2044\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17186\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__17186\,
            I => \b2v_inst11.count_1_5\
        );

    \I__2042\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__17180\,
            I => \b2v_inst11.count_0_5\
        );

    \I__2040\ : SRMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__17174\,
            I => \N__17171\
        );

    \I__2038\ : Odrv12
    port map (
            O => \N__17171\,
            I => \b2v_inst11.pwm_out_1_sqmuxa\
        );

    \I__2037\ : IoInMux
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17162\
        );

    \I__2035\ : Odrv12
    port map (
            O => \N__17162\,
            I => pwrbtn_led
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__17159\,
            I => \b2v_inst11.curr_state_3_0_cascade_\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__17156\,
            I => \b2v_inst11.curr_stateZ0Z_0_cascade_\
        );

    \I__2032\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17132\
        );

    \I__2031\ : InMux
    port map (
            O => \N__17152\,
            I => \N__17132\
        );

    \I__2030\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17132\
        );

    \I__2029\ : InMux
    port map (
            O => \N__17150\,
            I => \N__17123\
        );

    \I__2028\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17123\
        );

    \I__2027\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17123\
        );

    \I__2026\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17123\
        );

    \I__2025\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17114\
        );

    \I__2024\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17114\
        );

    \I__2023\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17114\
        );

    \I__2022\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17114\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__17142\,
            I => \N__17110\
        );

    \I__2020\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17102\
        );

    \I__2019\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17102\
        );

    \I__2018\ : InMux
    port map (
            O => \N__17139\,
            I => \N__17102\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__17132\,
            I => \N__17095\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17095\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__17114\,
            I => \N__17095\
        );

    \I__2014\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17088\
        );

    \I__2013\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17088\
        );

    \I__2012\ : InMux
    port map (
            O => \N__17109\,
            I => \N__17088\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__17102\,
            I => \N__17085\
        );

    \I__2010\ : Span4Mux_s2_v
    port map (
            O => \N__17095\,
            I => \N__17082\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__17088\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__17085\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__17082\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__17075\,
            I => \b2v_inst11.count_0_sqmuxa_i_cascade_\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__17072\,
            I => \b2v_inst11.count_1_0_cascade_\
        );

    \I__2004\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17066\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__17066\,
            I => \b2v_inst11.count_0_0\
        );

    \I__2002\ : InMux
    port map (
            O => \N__17063\,
            I => \N__17057\
        );

    \I__2001\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17057\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__17057\,
            I => \b2v_inst11.pwm_outZ0\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__17054\,
            I => \N__17050\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__17053\,
            I => \N__17047\
        );

    \I__1997\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17042\
        );

    \I__1996\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17042\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__17042\,
            I => \b2v_inst11.g0_i_o3_0\
        );

    \I__1994\ : InMux
    port map (
            O => \N__17039\,
            I => \b2v_inst11.mult1_un103_sum_cry_2\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__1992\ : InMux
    port map (
            O => \N__17033\,
            I => \N__17030\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__17030\,
            I => \b2v_inst11.mult1_un96_sum_cry_3_s\
        );

    \I__1990\ : InMux
    port map (
            O => \N__17027\,
            I => \b2v_inst11.mult1_un103_sum_cry_3\
        );

    \I__1989\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__17021\,
            I => \b2v_inst11.mult1_un96_sum_cry_4_s\
        );

    \I__1987\ : InMux
    port map (
            O => \N__17018\,
            I => \b2v_inst11.mult1_un103_sum_cry_4\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__17015\,
            I => \N__17010\
        );

    \I__1985\ : InMux
    port map (
            O => \N__17014\,
            I => \N__17006\
        );

    \I__1984\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17001\
        );

    \I__1983\ : InMux
    port map (
            O => \N__17010\,
            I => \N__17001\
        );

    \I__1982\ : InMux
    port map (
            O => \N__17009\,
            I => \N__16998\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__17006\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__17001\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__16998\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__1977\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__16985\,
            I => \b2v_inst11.mult1_un96_sum_cry_5_s\
        );

    \I__1975\ : InMux
    port map (
            O => \N__16982\,
            I => \b2v_inst11.mult1_un103_sum_cry_5\
        );

    \I__1974\ : InMux
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__16976\,
            I => \b2v_inst11.mult1_un96_sum_cry_6_s\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__16973\,
            I => \N__16969\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__16972\,
            I => \N__16965\
        );

    \I__1970\ : InMux
    port map (
            O => \N__16969\,
            I => \N__16958\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16968\,
            I => \N__16958\
        );

    \I__1968\ : InMux
    port map (
            O => \N__16965\,
            I => \N__16958\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__16958\,
            I => \b2v_inst11.mult1_un96_sum_i_0_8\
        );

    \I__1966\ : InMux
    port map (
            O => \N__16955\,
            I => \b2v_inst11.mult1_un103_sum_cry_6\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__16952\,
            I => \N__16949\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16946\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__16946\,
            I => \b2v_inst11.mult1_un103_sum_axb_8\
        );

    \I__1962\ : InMux
    port map (
            O => \N__16943\,
            I => \b2v_inst11.mult1_un103_sum_cry_7\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__16940\,
            I => \N__16935\
        );

    \I__1960\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16931\
        );

    \I__1959\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16926\
        );

    \I__1958\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16926\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16923\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__16931\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__16926\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__16923\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__1953\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__16913\,
            I => \b2v_inst11.mult1_un75_sum_cry_6_s\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__16910\,
            I => \N__16906\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__16909\,
            I => \N__16902\
        );

    \I__1949\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16895\
        );

    \I__1948\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16895\
        );

    \I__1947\ : InMux
    port map (
            O => \N__16902\,
            I => \N__16895\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__16895\,
            I => \b2v_inst11.mult1_un75_sum_i_0_8\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__1944\ : InMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__16886\,
            I => \b2v_inst11.mult1_un89_sum_axb_8\
        );

    \I__1942\ : InMux
    port map (
            O => \N__16883\,
            I => \b2v_inst11.mult1_un82_sum_cry_6\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \N__16877\
        );

    \I__1940\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16874\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__16874\,
            I => \b2v_inst11.mult1_un82_sum_axb_8\
        );

    \I__1938\ : InMux
    port map (
            O => \N__16871\,
            I => \b2v_inst11.mult1_un82_sum_cry_7\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__16868\,
            I => \N__16864\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__16867\,
            I => \N__16860\
        );

    \I__1935\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16853\
        );

    \I__1934\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16853\
        );

    \I__1933\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16853\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__16853\,
            I => \b2v_inst11.mult1_un54_sum_i_8\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__16850\,
            I => \N__16845\
        );

    \I__1930\ : InMux
    port map (
            O => \N__16849\,
            I => \N__16841\
        );

    \I__1929\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16836\
        );

    \I__1928\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16836\
        );

    \I__1927\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16833\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__16841\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__16836\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__16833\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__1923\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__16823\,
            I => \b2v_inst11.mult1_un68_sum_i\
        );

    \I__1921\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__16817\,
            I => \b2v_inst11.mult1_un82_sum_i\
        );

    \I__1919\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__1917\ : Span4Mux_s1_h
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__16805\,
            I => \b2v_inst11.mult1_un89_sum_i\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__16802\,
            I => \N__16798\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__16801\,
            I => \N__16794\
        );

    \I__1913\ : InMux
    port map (
            O => \N__16798\,
            I => \N__16787\
        );

    \I__1912\ : InMux
    port map (
            O => \N__16797\,
            I => \N__16787\
        );

    \I__1911\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16787\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__16787\,
            I => \b2v_inst11.mult1_un82_sum_i_0_8\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__16784\,
            I => \N__16780\
        );

    \I__1908\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16772\
        );

    \I__1907\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16772\
        );

    \I__1906\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16769\
        );

    \I__1905\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16764\
        );

    \I__1904\ : InMux
    port map (
            O => \N__16777\,
            I => \N__16764\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__16772\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__16769\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__16764\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__1899\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__16751\,
            I => \b2v_inst11.mult1_un68_sum_axb_8\
        );

    \I__1897\ : InMux
    port map (
            O => \N__16748\,
            I => \b2v_inst11.mult1_un61_sum_cry_6\
        );

    \I__1896\ : InMux
    port map (
            O => \N__16745\,
            I => \b2v_inst11.mult1_un61_sum_cry_7\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__16742\,
            I => \b2v_inst11.mult1_un61_sum_s_8_cascade_\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__16739\,
            I => \N__16735\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__16738\,
            I => \N__16731\
        );

    \I__1892\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16724\
        );

    \I__1891\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16724\
        );

    \I__1890\ : InMux
    port map (
            O => \N__16731\,
            I => \N__16724\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__16724\,
            I => \b2v_inst11.mult1_un61_sum_i_0_8\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__1887\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__16715\,
            I => \b2v_inst11.mult1_un82_sum_cry_3_s\
        );

    \I__1885\ : InMux
    port map (
            O => \N__16712\,
            I => \b2v_inst11.mult1_un82_sum_cry_2\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__16709\,
            I => \N__16706\
        );

    \I__1883\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__16703\,
            I => \b2v_inst11.mult1_un75_sum_cry_3_s\
        );

    \I__1881\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16697\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__16697\,
            I => \b2v_inst11.mult1_un82_sum_cry_4_s\
        );

    \I__1879\ : InMux
    port map (
            O => \N__16694\,
            I => \b2v_inst11.mult1_un82_sum_cry_3\
        );

    \I__1878\ : InMux
    port map (
            O => \N__16691\,
            I => \N__16688\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__16688\,
            I => \b2v_inst11.mult1_un75_sum_cry_4_s\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__1875\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__16679\,
            I => \b2v_inst11.mult1_un82_sum_cry_5_s\
        );

    \I__1873\ : InMux
    port map (
            O => \N__16676\,
            I => \b2v_inst11.mult1_un82_sum_cry_4\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__1871\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__16667\,
            I => \b2v_inst11.mult1_un75_sum_cry_5_s\
        );

    \I__1869\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__16661\,
            I => \b2v_inst11.mult1_un82_sum_cry_6_s\
        );

    \I__1867\ : InMux
    port map (
            O => \N__16658\,
            I => \b2v_inst11.mult1_un82_sum_cry_5\
        );

    \I__1866\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16649\
        );

    \I__1865\ : InMux
    port map (
            O => \N__16654\,
            I => \N__16649\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__16649\,
            I => \b2v_inst200.count_3_13\
        );

    \I__1863\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16637\
        );

    \I__1862\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16637\
        );

    \I__1861\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16637\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__16637\,
            I => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\
        );

    \I__1859\ : InMux
    port map (
            O => \N__16634\,
            I => \N__16631\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__16631\,
            I => \b2v_inst200.un2_count_1_axb_13\
        );

    \I__1857\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16625\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__16622\,
            I => \N__16617\
        );

    \I__1854\ : InMux
    port map (
            O => \N__16621\,
            I => \N__16612\
        );

    \I__1853\ : InMux
    port map (
            O => \N__16620\,
            I => \N__16612\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__16617\,
            I => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__16612\,
            I => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\
        );

    \I__1850\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16603\
        );

    \I__1849\ : InMux
    port map (
            O => \N__16606\,
            I => \N__16600\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__16603\,
            I => \b2v_inst200.count_3_5\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__16600\,
            I => \b2v_inst200.count_3_5\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__1845\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16588\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__16591\,
            I => \N__16585\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__16588\,
            I => \N__16582\
        );

    \I__1842\ : InMux
    port map (
            O => \N__16585\,
            I => \N__16579\
        );

    \I__1841\ : Odrv12
    port map (
            O => \N__16582\,
            I => \b2v_inst200.countZ0Z_7\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__16579\,
            I => \b2v_inst200.countZ0Z_7\
        );

    \I__1839\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16540\
        );

    \I__1838\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16540\
        );

    \I__1837\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16540\
        );

    \I__1836\ : InMux
    port map (
            O => \N__16571\,
            I => \N__16540\
        );

    \I__1835\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16529\
        );

    \I__1834\ : InMux
    port map (
            O => \N__16569\,
            I => \N__16529\
        );

    \I__1833\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16529\
        );

    \I__1832\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16529\
        );

    \I__1831\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16529\
        );

    \I__1830\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16524\
        );

    \I__1829\ : InMux
    port map (
            O => \N__16564\,
            I => \N__16524\
        );

    \I__1828\ : InMux
    port map (
            O => \N__16563\,
            I => \N__16515\
        );

    \I__1827\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16515\
        );

    \I__1826\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16515\
        );

    \I__1825\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16515\
        );

    \I__1824\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16502\
        );

    \I__1823\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16502\
        );

    \I__1822\ : InMux
    port map (
            O => \N__16557\,
            I => \N__16502\
        );

    \I__1821\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16502\
        );

    \I__1820\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16502\
        );

    \I__1819\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16502\
        );

    \I__1818\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16491\
        );

    \I__1817\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16491\
        );

    \I__1816\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16491\
        );

    \I__1815\ : InMux
    port map (
            O => \N__16550\,
            I => \N__16491\
        );

    \I__1814\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16491\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__16540\,
            I => \N__16482\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__16529\,
            I => \N__16479\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__16524\,
            I => \N__16476\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__16515\,
            I => \N__16473\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__16502\,
            I => \N__16470\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__16491\,
            I => \N__16467\
        );

    \I__1807\ : CEMux
    port map (
            O => \N__16490\,
            I => \N__16442\
        );

    \I__1806\ : CEMux
    port map (
            O => \N__16489\,
            I => \N__16442\
        );

    \I__1805\ : CEMux
    port map (
            O => \N__16488\,
            I => \N__16442\
        );

    \I__1804\ : CEMux
    port map (
            O => \N__16487\,
            I => \N__16442\
        );

    \I__1803\ : CEMux
    port map (
            O => \N__16486\,
            I => \N__16442\
        );

    \I__1802\ : CEMux
    port map (
            O => \N__16485\,
            I => \N__16442\
        );

    \I__1801\ : Glb2LocalMux
    port map (
            O => \N__16482\,
            I => \N__16442\
        );

    \I__1800\ : Glb2LocalMux
    port map (
            O => \N__16479\,
            I => \N__16442\
        );

    \I__1799\ : Glb2LocalMux
    port map (
            O => \N__16476\,
            I => \N__16442\
        );

    \I__1798\ : Glb2LocalMux
    port map (
            O => \N__16473\,
            I => \N__16442\
        );

    \I__1797\ : Glb2LocalMux
    port map (
            O => \N__16470\,
            I => \N__16442\
        );

    \I__1796\ : Glb2LocalMux
    port map (
            O => \N__16467\,
            I => \N__16442\
        );

    \I__1795\ : GlobalMux
    port map (
            O => \N__16442\,
            I => \N__16439\
        );

    \I__1794\ : gio2CtrlBuf
    port map (
            O => \N__16439\,
            I => \b2v_inst200.count_en_g\
        );

    \I__1793\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__16433\,
            I => \b2v_inst200.un25_clk_100khz_3\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__16430\,
            I => \N__16427\
        );

    \I__1790\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16424\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__16424\,
            I => \b2v_inst11.mult1_un61_sum_cry_3_s\
        );

    \I__1788\ : InMux
    port map (
            O => \N__16421\,
            I => \b2v_inst11.mult1_un61_sum_cry_2\
        );

    \I__1787\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16415\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__16415\,
            I => \b2v_inst11.mult1_un61_sum_cry_4_s\
        );

    \I__1785\ : InMux
    port map (
            O => \N__16412\,
            I => \b2v_inst11.mult1_un61_sum_cry_3\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__1783\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__16403\,
            I => \b2v_inst11.mult1_un61_sum_cry_5_s\
        );

    \I__1781\ : InMux
    port map (
            O => \N__16400\,
            I => \b2v_inst11.mult1_un61_sum_cry_4\
        );

    \I__1780\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__16394\,
            I => \b2v_inst11.mult1_un61_sum_cry_6_s\
        );

    \I__1778\ : InMux
    port map (
            O => \N__16391\,
            I => \b2v_inst11.mult1_un61_sum_cry_5\
        );

    \I__1777\ : InMux
    port map (
            O => \N__16388\,
            I => \N__16382\
        );

    \I__1776\ : InMux
    port map (
            O => \N__16387\,
            I => \N__16382\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__16382\,
            I => \b2v_inst200.count_3_9\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__16379\,
            I => \b2v_inst200.countZ0Z_12_cascade_\
        );

    \I__1773\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16367\
        );

    \I__1772\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16367\
        );

    \I__1771\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16367\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__16367\,
            I => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\
        );

    \I__1769\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__16361\,
            I => \b2v_inst200.un2_count_1_axb_5\
        );

    \I__1767\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16355\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__16352\,
            I => \b2v_inst200.count_3_11\
        );

    \I__1764\ : InMux
    port map (
            O => \N__16349\,
            I => \N__16346\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__16346\,
            I => \N__16342\
        );

    \I__1762\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16339\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__16342\,
            I => \b2v_inst200.count_1_11\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__16339\,
            I => \b2v_inst200.count_1_11\
        );

    \I__1759\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__1757\ : Span4Mux_s1_h
    port map (
            O => \N__16328\,
            I => \N__16324\
        );

    \I__1756\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16321\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__16324\,
            I => \b2v_inst200.countZ0Z_11\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__16321\,
            I => \b2v_inst200.countZ0Z_11\
        );

    \I__1753\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16313\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__16313\,
            I => \N__16310\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__16310\,
            I => \b2v_inst200.un2_count_1_axb_3\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__16307\,
            I => \N__16304\
        );

    \I__1749\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16300\
        );

    \I__1748\ : InMux
    port map (
            O => \N__16303\,
            I => \N__16297\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__16300\,
            I => \N__16292\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__16297\,
            I => \N__16292\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__16292\,
            I => \b2v_inst200.countZ0Z_14\
        );

    \I__1744\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16286\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__16286\,
            I => \b2v_inst200.un25_clk_100khz_4\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__16283\,
            I => \b2v_inst200.un25_clk_100khz_5_cascade_\
        );

    \I__1741\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16277\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__16277\,
            I => \N__16274\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__16274\,
            I => \b2v_inst200.un25_clk_100khz_14\
        );

    \I__1738\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16265\
        );

    \I__1737\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16265\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__16265\,
            I => \b2v_inst200.count_3_3\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__16262\,
            I => \N__16259\
        );

    \I__1734\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16256\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__16256\,
            I => \N__16252\
        );

    \I__1732\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16249\
        );

    \I__1731\ : Span12Mux_v
    port map (
            O => \N__16252\,
            I => \N__16246\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__16249\,
            I => \N__16243\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__16246\,
            I => \b2v_inst200.countZ0Z_4\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__16243\,
            I => \b2v_inst200.countZ0Z_4\
        );

    \I__1727\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16229\
        );

    \I__1726\ : InMux
    port map (
            O => \N__16237\,
            I => \N__16229\
        );

    \I__1725\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16229\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__16229\,
            I => \N__16226\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__16226\,
            I => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\
        );

    \I__1722\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16220\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__16220\,
            I => \b2v_inst200.un25_clk_100khz_2\
        );

    \I__1720\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16208\
        );

    \I__1719\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16208\
        );

    \I__1718\ : InMux
    port map (
            O => \N__16215\,
            I => \N__16208\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__16208\,
            I => \b2v_inst200.count_1_8\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__16205\,
            I => \N__16202\
        );

    \I__1715\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16196\
        );

    \I__1714\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16196\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__16196\,
            I => \b2v_inst200.count_3_8\
        );

    \I__1712\ : InMux
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__16190\,
            I => \b2v_inst200.un2_count_1_axb_8\
        );

    \I__1710\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__16184\,
            I => \b2v_inst200.un2_count_1_axb_15\
        );

    \I__1708\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16175\
        );

    \I__1707\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16175\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__16175\,
            I => \b2v_inst200.count_3_15\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__16172\,
            I => \N__16167\
        );

    \I__1704\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16160\
        );

    \I__1703\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16160\
        );

    \I__1702\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16160\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__16160\,
            I => \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__16157\,
            I => \N__16153\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__16156\,
            I => \N__16150\
        );

    \I__1698\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16147\
        );

    \I__1697\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16144\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__16147\,
            I => \b2v_inst200.countZ0Z_6\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__16144\,
            I => \b2v_inst200.countZ0Z_6\
        );

    \I__1694\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16136\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__16136\,
            I => \b2v_inst200.un25_clk_100khz_7\
        );

    \I__1692\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16130\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__16130\,
            I => \N__16127\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__16124\,
            I => \b2v_inst200.un25_clk_100khz_13\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__16121\,
            I => \b2v_inst200.un25_clk_100khz_6_cascade_\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__16118\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_\
        );

    \I__1686\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16111\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__16114\,
            I => \N__16107\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__16111\,
            I => \N__16101\
        );

    \I__1683\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16098\
        );

    \I__1682\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16095\
        );

    \I__1681\ : InMux
    port map (
            O => \N__16106\,
            I => \N__16088\
        );

    \I__1680\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16088\
        );

    \I__1679\ : InMux
    port map (
            O => \N__16104\,
            I => \N__16088\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__16101\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__16098\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__16095\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__16088\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__1674\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16076\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__16076\,
            I => \b2v_inst200.count_3_0\
        );

    \I__1672\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16070\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__16070\,
            I => \b2v_inst200.un2_count_1_axb_9\
        );

    \I__1670\ : InMux
    port map (
            O => \N__16067\,
            I => \N__16064\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__16064\,
            I => \b2v_inst200.count_3_12\
        );

    \I__1668\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16055\
        );

    \I__1667\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16055\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__16055\,
            I => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\
        );

    \I__1665\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16049\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__16049\,
            I => \b2v_inst200.countZ0Z_12\
        );

    \I__1663\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__16043\,
            I => \b2v_inst200.count_3_6\
        );

    \I__1661\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16036\
        );

    \I__1660\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16033\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__16036\,
            I => \b2v_inst200.count_1_6\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__16033\,
            I => \b2v_inst200.count_1_6\
        );

    \I__1657\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__16025\,
            I => \b2v_inst200.count_3_7\
        );

    \I__1655\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16018\
        );

    \I__1654\ : InMux
    port map (
            O => \N__16021\,
            I => \N__16015\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__16018\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__16015\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__1651\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__1649\ : Span4Mux_h
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__16001\,
            I => \b2v_inst200.count_0_17\
        );

    \I__1647\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__15995\,
            I => \N__15991\
        );

    \I__1645\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15988\
        );

    \I__1644\ : Span4Mux_h
    port map (
            O => \N__15991\,
            I => \N__15985\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__15988\,
            I => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__15985\,
            I => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\
        );

    \I__1641\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__15977\,
            I => \N__15973\
        );

    \I__1639\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15970\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__15973\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__15970\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__15965\,
            I => \N__15961\
        );

    \I__1635\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15958\
        );

    \I__1634\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15955\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__15958\,
            I => \N__15950\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__15955\,
            I => \N__15950\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__15950\,
            I => \b2v_inst200.count_1_10\
        );

    \I__1630\ : InMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__15941\,
            I => \b2v_inst200.count_3_10\
        );

    \I__1627\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15935\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__15935\,
            I => \N__15932\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__15932\,
            I => \b2v_inst200.count_1_0\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__1623\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15922\
        );

    \I__1622\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15919\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__15922\,
            I => \N__15916\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__15919\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__15916\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__1618\ : InMux
    port map (
            O => \N__15911\,
            I => \N__15906\
        );

    \I__1617\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15901\
        );

    \I__1616\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15901\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__15906\,
            I => \N__15898\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__15901\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1613\ : Odrv4
    port map (
            O => \N__15898\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1612\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15887\
        );

    \I__1611\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15887\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__15884\,
            I => \b2v_inst16.un4_count_1_cry_10_THRU_CO\
        );

    \I__1608\ : InMux
    port map (
            O => \N__15881\,
            I => \b2v_inst16.un4_count_1_cry_10\
        );

    \I__1607\ : InMux
    port map (
            O => \N__15878\,
            I => \b2v_inst16.un4_count_1_cry_11\
        );

    \I__1606\ : InMux
    port map (
            O => \N__15875\,
            I => \b2v_inst16.un4_count_1_cry_12\
        );

    \I__1605\ : InMux
    port map (
            O => \N__15872\,
            I => \b2v_inst16.un4_count_1_cry_13\
        );

    \I__1604\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15866\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15862\
        );

    \I__1602\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15859\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__15862\,
            I => \b2v_inst16.countZ0Z_15\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__15859\,
            I => \b2v_inst16.countZ0Z_15\
        );

    \I__1599\ : InMux
    port map (
            O => \N__15854\,
            I => \b2v_inst16.un4_count_1_cry_14\
        );

    \I__1598\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15847\
        );

    \I__1597\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15844\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__15847\,
            I => \b2v_inst16.count_rst_4\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__15844\,
            I => \b2v_inst16.count_rst_4\
        );

    \I__1594\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15836\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__15836\,
            I => \b2v_inst200.count_3_14\
        );

    \I__1592\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15829\
        );

    \I__1591\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15826\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__15829\,
            I => \N__15821\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__15826\,
            I => \N__15821\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__15821\,
            I => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\
        );

    \I__1587\ : InMux
    port map (
            O => \N__15818\,
            I => \b2v_inst16.un4_count_1_cry_1\
        );

    \I__1586\ : InMux
    port map (
            O => \N__15815\,
            I => \b2v_inst16.un4_count_1_cry_2\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__15812\,
            I => \N__15809\
        );

    \I__1584\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15804\
        );

    \I__1583\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15801\
        );

    \I__1582\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15798\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__15804\,
            I => \N__15795\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__15801\,
            I => \N__15790\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__15798\,
            I => \N__15790\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__15795\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__15790\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1576\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15779\
        );

    \I__1575\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15779\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__15776\,
            I => \b2v_inst16.un4_count_1_cry_3_THRU_CO\
        );

    \I__1572\ : InMux
    port map (
            O => \N__15773\,
            I => \b2v_inst16.un4_count_1_cry_3\
        );

    \I__1571\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15765\
        );

    \I__1570\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15762\
        );

    \I__1569\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15759\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__15765\,
            I => \N__15756\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__15762\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__15759\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__15756\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1564\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15743\
        );

    \I__1563\ : InMux
    port map (
            O => \N__15748\,
            I => \N__15743\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__15743\,
            I => \N__15740\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__15740\,
            I => \b2v_inst16.un4_count_1_cry_4_THRU_CO\
        );

    \I__1560\ : InMux
    port map (
            O => \N__15737\,
            I => \b2v_inst16.un4_count_1_cry_4\
        );

    \I__1559\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15730\
        );

    \I__1558\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15727\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__15730\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__15727\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1555\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15716\
        );

    \I__1554\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15716\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__15716\,
            I => \b2v_inst16.count_rst_11\
        );

    \I__1552\ : InMux
    port map (
            O => \N__15713\,
            I => \b2v_inst16.un4_count_1_cry_5\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__15710\,
            I => \N__15705\
        );

    \I__1550\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15701\
        );

    \I__1549\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15698\
        );

    \I__1548\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15695\
        );

    \I__1547\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15692\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__15701\,
            I => \N__15689\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__15698\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__15695\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__15692\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__15689\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1541\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15676\
        );

    \I__1540\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15673\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__15676\,
            I => \N__15668\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__15673\,
            I => \N__15668\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__15668\,
            I => \b2v_inst16.un4_count_1_cry_6_THRU_CO\
        );

    \I__1536\ : InMux
    port map (
            O => \N__15665\,
            I => \b2v_inst16.un4_count_1_cry_6\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__15662\,
            I => \N__15658\
        );

    \I__1534\ : InMux
    port map (
            O => \N__15661\,
            I => \N__15653\
        );

    \I__1533\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15650\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15645\
        );

    \I__1531\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15645\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__15653\,
            I => \N__15642\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__15650\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__15645\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__15642\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__15635\,
            I => \N__15631\
        );

    \I__1525\ : InMux
    port map (
            O => \N__15634\,
            I => \N__15628\
        );

    \I__1524\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15625\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__15628\,
            I => \N__15622\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__15625\,
            I => \b2v_inst16.un4_count_1_cry_7_THRU_CO\
        );

    \I__1521\ : Odrv4
    port map (
            O => \N__15622\,
            I => \b2v_inst16.un4_count_1_cry_7_THRU_CO\
        );

    \I__1520\ : InMux
    port map (
            O => \N__15617\,
            I => \b2v_inst16.un4_count_1_cry_7\
        );

    \I__1519\ : InMux
    port map (
            O => \N__15614\,
            I => \N__15609\
        );

    \I__1518\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15606\
        );

    \I__1517\ : InMux
    port map (
            O => \N__15612\,
            I => \N__15603\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__15609\,
            I => \N__15598\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__15606\,
            I => \N__15598\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__15603\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__15598\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__15593\,
            I => \N__15589\
        );

    \I__1511\ : InMux
    port map (
            O => \N__15592\,
            I => \N__15586\
        );

    \I__1510\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15583\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__15586\,
            I => \N__15578\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__15583\,
            I => \N__15578\
        );

    \I__1507\ : Span4Mux_s1_h
    port map (
            O => \N__15578\,
            I => \N__15575\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__15575\,
            I => \b2v_inst16.un4_count_1_cry_8_THRU_CO\
        );

    \I__1505\ : InMux
    port map (
            O => \N__15572\,
            I => \bfn_2_4_0_\
        );

    \I__1504\ : InMux
    port map (
            O => \N__15569\,
            I => \b2v_inst16.un4_count_1_cry_9\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__15566\,
            I => \b2v_inst16.countZ0Z_2_cascade_\
        );

    \I__1502\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__15560\,
            I => \b2v_inst16.count_4_i_a3_8_0\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__15557\,
            I => \b2v_inst16.count_4_i_a3_9_0_cascade_\
        );

    \I__1499\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15551\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__15551\,
            I => \b2v_inst16.count_4_i_a3_7_0\
        );

    \I__1497\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15545\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__15545\,
            I => \b2v_inst16.count_rst_5\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__15542\,
            I => \b2v_inst16.countZ0Z_0_cascade_\
        );

    \I__1494\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15534\
        );

    \I__1493\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15531\
        );

    \I__1492\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15528\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__15534\,
            I => \b2v_inst16.N_414\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__15531\,
            I => \b2v_inst16.N_414\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__15528\,
            I => \b2v_inst16.N_414\
        );

    \I__1488\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15518\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__15518\,
            I => \b2v_inst16.count_4_0\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__15515\,
            I => \N__15512\
        );

    \I__1485\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15506\
        );

    \I__1484\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15506\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__15506\,
            I => \b2v_inst16.count_4_2\
        );

    \I__1482\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15494\
        );

    \I__1481\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15494\
        );

    \I__1480\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15491\
        );

    \I__1479\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15486\
        );

    \I__1478\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15486\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__15494\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__15491\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__15486\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__15479\,
            I => \N__15474\
        );

    \I__1473\ : InMux
    port map (
            O => \N__15478\,
            I => \N__15469\
        );

    \I__1472\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15469\
        );

    \I__1471\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15466\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__15469\,
            I => \b2v_inst16.countZ0Z_1\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__15466\,
            I => \b2v_inst16.countZ0Z_1\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__1467\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__15455\,
            I => \b2v_inst16.un4_count_1_axb_2\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__15452\,
            I => \N__15448\
        );

    \I__1464\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15440\
        );

    \I__1463\ : InMux
    port map (
            O => \N__15448\,
            I => \N__15440\
        );

    \I__1462\ : InMux
    port map (
            O => \N__15447\,
            I => \N__15440\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__15440\,
            I => \b2v_inst16.un4_count_1_cry_1_c_RNIAGMEZ0\
        );

    \I__1460\ : InMux
    port map (
            O => \N__15437\,
            I => \b2v_inst11.un1_count_cry_14\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__15434\,
            I => \b2v_inst16.count_rst_9_cascade_\
        );

    \I__1458\ : CascadeMux
    port map (
            O => \N__15431\,
            I => \b2v_inst16.countZ0Z_4_cascade_\
        );

    \I__1457\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__15425\,
            I => \b2v_inst16.count_4_4\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__15422\,
            I => \b2v_inst16.count_rst_10_cascade_\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__15419\,
            I => \b2v_inst16.countZ0Z_5_cascade_\
        );

    \I__1453\ : InMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__15413\,
            I => \b2v_inst16.count_4_5\
        );

    \I__1451\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15407\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__15407\,
            I => \b2v_inst16.count_4_7\
        );

    \I__1449\ : InMux
    port map (
            O => \N__15404\,
            I => \b2v_inst11.un1_count_cry_6\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__15401\,
            I => \N__15398\
        );

    \I__1447\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15392\
        );

    \I__1446\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15392\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__15392\,
            I => \N__15389\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__15389\,
            I => \b2v_inst11.count_1_8\
        );

    \I__1443\ : InMux
    port map (
            O => \N__15386\,
            I => \b2v_inst11.un1_count_cry_7\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__15383\,
            I => \N__15380\
        );

    \I__1441\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15374\
        );

    \I__1440\ : InMux
    port map (
            O => \N__15379\,
            I => \N__15374\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__15374\,
            I => \N__15371\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__15371\,
            I => \b2v_inst11.count_1_9\
        );

    \I__1437\ : InMux
    port map (
            O => \N__15368\,
            I => \bfn_1_16_0_\
        );

    \I__1436\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15359\
        );

    \I__1435\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15359\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__15359\,
            I => \N__15356\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__15356\,
            I => \b2v_inst11.count_1_10\
        );

    \I__1432\ : InMux
    port map (
            O => \N__15353\,
            I => \b2v_inst11.un1_count_cry_9\
        );

    \I__1431\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15344\
        );

    \I__1430\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15344\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__15344\,
            I => \N__15341\
        );

    \I__1428\ : Odrv4
    port map (
            O => \N__15341\,
            I => \b2v_inst11.count_1_11\
        );

    \I__1427\ : InMux
    port map (
            O => \N__15338\,
            I => \b2v_inst11.un1_count_cry_10\
        );

    \I__1426\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15329\
        );

    \I__1425\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15329\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__15326\,
            I => \b2v_inst11.count_1_12\
        );

    \I__1422\ : InMux
    port map (
            O => \N__15323\,
            I => \b2v_inst11.un1_count_cry_11\
        );

    \I__1421\ : InMux
    port map (
            O => \N__15320\,
            I => \b2v_inst11.un1_count_cry_12\
        );

    \I__1420\ : InMux
    port map (
            O => \N__15317\,
            I => \b2v_inst11.un1_count_cry_13\
        );

    \I__1419\ : InMux
    port map (
            O => \N__15314\,
            I => \N__15311\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__15311\,
            I => \b2v_inst11.count_0_2\
        );

    \I__1417\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15305\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__15305\,
            I => \b2v_inst11.count_0_12\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__15302\,
            I => \N__15298\
        );

    \I__1414\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15293\
        );

    \I__1413\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15293\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__15293\,
            I => \b2v_inst11.count_1_2\
        );

    \I__1411\ : InMux
    port map (
            O => \N__15290\,
            I => \b2v_inst11.un1_count_cry_1_cZ0\
        );

    \I__1410\ : InMux
    port map (
            O => \N__15287\,
            I => \b2v_inst11.un1_count_cry_2\
        );

    \I__1409\ : InMux
    port map (
            O => \N__15284\,
            I => \b2v_inst11.un1_count_cry_3\
        );

    \I__1408\ : InMux
    port map (
            O => \N__15281\,
            I => \b2v_inst11.un1_count_cry_4\
        );

    \I__1407\ : InMux
    port map (
            O => \N__15278\,
            I => \b2v_inst11.un1_count_cry_5\
        );

    \I__1406\ : InMux
    port map (
            O => \N__15275\,
            I => \N__15272\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__15272\,
            I => \b2v_inst11.count_0_9\
        );

    \I__1404\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15266\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__15266\,
            I => \b2v_inst11.count_0_10\
        );

    \I__1402\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__15260\,
            I => \b2v_inst11.count_0_11\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \b2v_inst11.count_1_1_cascade_\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__15254\,
            I => \b2v_inst11.countZ0Z_1_cascade_\
        );

    \I__1398\ : InMux
    port map (
            O => \N__15251\,
            I => \N__15248\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__15248\,
            I => \b2v_inst11.count_0_1\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__1395\ : InMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__15239\,
            I => \b2v_inst11.mult1_un89_sum_cry_3_s\
        );

    \I__1393\ : InMux
    port map (
            O => \N__15236\,
            I => \b2v_inst11.mult1_un96_sum_cry_3\
        );

    \I__1392\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__15230\,
            I => \b2v_inst11.mult1_un89_sum_cry_4_s\
        );

    \I__1390\ : InMux
    port map (
            O => \N__15227\,
            I => \b2v_inst11.mult1_un96_sum_cry_4\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__1388\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15218\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__15218\,
            I => \b2v_inst11.mult1_un89_sum_cry_5_s\
        );

    \I__1386\ : InMux
    port map (
            O => \N__15215\,
            I => \b2v_inst11.mult1_un96_sum_cry_5\
        );

    \I__1385\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15209\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__15209\,
            I => \b2v_inst11.mult1_un89_sum_cry_6_s\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__15206\,
            I => \N__15202\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__15205\,
            I => \N__15198\
        );

    \I__1381\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15191\
        );

    \I__1380\ : InMux
    port map (
            O => \N__15201\,
            I => \N__15191\
        );

    \I__1379\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15191\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__15191\,
            I => \b2v_inst11.mult1_un89_sum_i_0_8\
        );

    \I__1377\ : InMux
    port map (
            O => \N__15188\,
            I => \b2v_inst11.mult1_un96_sum_cry_6\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__15185\,
            I => \N__15182\
        );

    \I__1375\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15179\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__15179\,
            I => \b2v_inst11.mult1_un96_sum_axb_8\
        );

    \I__1373\ : InMux
    port map (
            O => \N__15176\,
            I => \b2v_inst11.mult1_un96_sum_cry_7\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__15173\,
            I => \b2v_inst11.mult1_un96_sum_s_8_cascade_\
        );

    \I__1371\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__15167\,
            I => \b2v_inst11.count_0_8\
        );

    \I__1369\ : InMux
    port map (
            O => \N__15164\,
            I => \b2v_inst11.mult1_un89_sum_cry_2\
        );

    \I__1368\ : InMux
    port map (
            O => \N__15161\,
            I => \b2v_inst11.mult1_un89_sum_cry_3\
        );

    \I__1367\ : InMux
    port map (
            O => \N__15158\,
            I => \b2v_inst11.mult1_un89_sum_cry_4\
        );

    \I__1366\ : InMux
    port map (
            O => \N__15155\,
            I => \b2v_inst11.mult1_un89_sum_cry_5\
        );

    \I__1365\ : InMux
    port map (
            O => \N__15152\,
            I => \b2v_inst11.mult1_un89_sum_cry_6\
        );

    \I__1364\ : InMux
    port map (
            O => \N__15149\,
            I => \b2v_inst11.mult1_un89_sum_cry_7\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__15146\,
            I => \b2v_inst11.mult1_un89_sum_s_8_cascade_\
        );

    \I__1362\ : InMux
    port map (
            O => \N__15143\,
            I => \b2v_inst11.mult1_un96_sum_cry_2\
        );

    \I__1361\ : InMux
    port map (
            O => \N__15140\,
            I => \b2v_inst11.mult1_un75_sum_cry_2\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__15137\,
            I => \N__15134\
        );

    \I__1359\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15131\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__15131\,
            I => \b2v_inst11.mult1_un68_sum_cry_3_s\
        );

    \I__1357\ : InMux
    port map (
            O => \N__15128\,
            I => \b2v_inst11.mult1_un75_sum_cry_3\
        );

    \I__1356\ : InMux
    port map (
            O => \N__15125\,
            I => \N__15122\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__15122\,
            I => \b2v_inst11.mult1_un68_sum_cry_4_s\
        );

    \I__1354\ : InMux
    port map (
            O => \N__15119\,
            I => \b2v_inst11.mult1_un75_sum_cry_4\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__15116\,
            I => \N__15113\
        );

    \I__1352\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__15110\,
            I => \b2v_inst11.mult1_un68_sum_cry_5_s\
        );

    \I__1350\ : InMux
    port map (
            O => \N__15107\,
            I => \b2v_inst11.mult1_un75_sum_cry_5\
        );

    \I__1349\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__15101\,
            I => \b2v_inst11.mult1_un68_sum_cry_6_s\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__15098\,
            I => \N__15094\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__15097\,
            I => \N__15090\
        );

    \I__1345\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15083\
        );

    \I__1344\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15083\
        );

    \I__1343\ : InMux
    port map (
            O => \N__15090\,
            I => \N__15083\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__15083\,
            I => \b2v_inst11.mult1_un68_sum_i_0_8\
        );

    \I__1341\ : InMux
    port map (
            O => \N__15080\,
            I => \b2v_inst11.mult1_un75_sum_cry_6\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__1339\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__15071\,
            I => \b2v_inst11.mult1_un75_sum_axb_8\
        );

    \I__1337\ : InMux
    port map (
            O => \N__15068\,
            I => \b2v_inst11.mult1_un75_sum_cry_7\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__15065\,
            I => \b2v_inst11.mult1_un75_sum_s_8_cascade_\
        );

    \I__1335\ : InMux
    port map (
            O => \N__15062\,
            I => \b2v_inst11.mult1_un68_sum_cry_2\
        );

    \I__1334\ : InMux
    port map (
            O => \N__15059\,
            I => \b2v_inst11.mult1_un68_sum_cry_3\
        );

    \I__1333\ : InMux
    port map (
            O => \N__15056\,
            I => \b2v_inst11.mult1_un68_sum_cry_4\
        );

    \I__1332\ : InMux
    port map (
            O => \N__15053\,
            I => \b2v_inst11.mult1_un68_sum_cry_5\
        );

    \I__1331\ : InMux
    port map (
            O => \N__15050\,
            I => \b2v_inst11.mult1_un68_sum_cry_6\
        );

    \I__1330\ : InMux
    port map (
            O => \N__15047\,
            I => \b2v_inst11.mult1_un68_sum_cry_7\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__15044\,
            I => \b2v_inst11.mult1_un68_sum_s_8_cascade_\
        );

    \I__1328\ : InMux
    port map (
            O => \N__15041\,
            I => \b2v_inst200.un2_count_1_cry_9\
        );

    \I__1327\ : InMux
    port map (
            O => \N__15038\,
            I => \b2v_inst200.un2_count_1_cry_10\
        );

    \I__1326\ : InMux
    port map (
            O => \N__15035\,
            I => \b2v_inst200.un2_count_1_cry_11\
        );

    \I__1325\ : InMux
    port map (
            O => \N__15032\,
            I => \b2v_inst200.un2_count_1_cry_12\
        );

    \I__1324\ : InMux
    port map (
            O => \N__15029\,
            I => \b2v_inst200.un2_count_1_cry_13\
        );

    \I__1323\ : InMux
    port map (
            O => \N__15026\,
            I => \b2v_inst200.un2_count_1_cry_14\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__1321\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15017\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__1319\ : Odrv12
    port map (
            O => \N__15014\,
            I => \b2v_inst200.un2_count_1_axb_16\
        );

    \I__1318\ : InMux
    port map (
            O => \N__15011\,
            I => \N__15002\
        );

    \I__1317\ : InMux
    port map (
            O => \N__15010\,
            I => \N__15002\
        );

    \I__1316\ : InMux
    port map (
            O => \N__15009\,
            I => \N__15002\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__1314\ : Odrv12
    port map (
            O => \N__14999\,
            I => \b2v_inst200.count_1_16\
        );

    \I__1313\ : InMux
    port map (
            O => \N__14996\,
            I => \b2v_inst200.un2_count_1_cry_15\
        );

    \I__1312\ : InMux
    port map (
            O => \N__14993\,
            I => \bfn_1_8_0_\
        );

    \I__1311\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14986\
        );

    \I__1310\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14983\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__14986\,
            I => \N__14980\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__14983\,
            I => \b2v_inst200.un2_count_1_axb_1\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__14980\,
            I => \b2v_inst200.un2_count_1_axb_1\
        );

    \I__1306\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14971\
        );

    \I__1305\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14968\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__14971\,
            I => \N__14965\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__14968\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__14965\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__1301\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14956\
        );

    \I__1300\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14953\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__14956\,
            I => \N__14950\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__14953\,
            I => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\
        );

    \I__1297\ : Odrv4
    port map (
            O => \N__14950\,
            I => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14945\,
            I => \b2v_inst200.un2_count_1_cry_1\
        );

    \I__1295\ : InMux
    port map (
            O => \N__14942\,
            I => \b2v_inst200.un2_count_1_cry_2\
        );

    \I__1294\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14935\
        );

    \I__1293\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14932\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__14935\,
            I => \N__14929\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__14932\,
            I => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__14929\,
            I => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\
        );

    \I__1289\ : InMux
    port map (
            O => \N__14924\,
            I => \b2v_inst200.un2_count_1_cry_3\
        );

    \I__1288\ : InMux
    port map (
            O => \N__14921\,
            I => \b2v_inst200.un2_count_1_cry_4\
        );

    \I__1287\ : InMux
    port map (
            O => \N__14918\,
            I => \b2v_inst200.un2_count_1_cry_5_cZ0\
        );

    \I__1286\ : InMux
    port map (
            O => \N__14915\,
            I => \b2v_inst200.un2_count_1_cry_6\
        );

    \I__1285\ : InMux
    port map (
            O => \N__14912\,
            I => \b2v_inst200.un2_count_1_cry_7\
        );

    \I__1284\ : InMux
    port map (
            O => \N__14909\,
            I => \bfn_1_7_0_\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__14906\,
            I => \b2v_inst200.count_RNIZ0Z_1_cascade_\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__14903\,
            I => \b2v_inst200.un2_count_1_axb_1_cascade_\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \N__14897\
        );

    \I__1280\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14893\
        );

    \I__1279\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14890\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__14893\,
            I => \b2v_inst200.count_3_1\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__14890\,
            I => \b2v_inst200.count_3_1\
        );

    \I__1276\ : InMux
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__14879\,
            I => \b2v_inst200.count_3_2\
        );

    \I__1273\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__14870\,
            I => \b2v_inst200.count_3_4\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__14867\,
            I => \b2v_inst200.un25_clk_100khz_1_cascade_\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__1268\ : InMux
    port map (
            O => \N__14861\,
            I => \N__14857\
        );

    \I__1267\ : InMux
    port map (
            O => \N__14860\,
            I => \N__14854\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__14857\,
            I => \b2v_inst200.countZ0Z_16\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__14854\,
            I => \b2v_inst200.countZ0Z_16\
        );

    \I__1264\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14846\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__14846\,
            I => \b2v_inst200.un25_clk_100khz_0\
        );

    \I__1262\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14840\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__14840\,
            I => \b2v_inst200.count_RNIZ0Z_1\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__14837\,
            I => \b2v_inst16.countZ0Z_1_cascade_\
        );

    \I__1259\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14831\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__14831\,
            I => \b2v_inst16.count_4_1\
        );

    \I__1257\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__14825\,
            I => \b2v_inst16.count_4_11\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__14822\,
            I => \b2v_inst16.count_rst_0_cascade_\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__14819\,
            I => \b2v_inst16.countZ0Z_11_cascade_\
        );

    \I__1253\ : InMux
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__14813\,
            I => \b2v_inst16.count_4_8\
        );

    \I__1251\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__14807\,
            I => \b2v_inst16.count_4_6\
        );

    \I__1249\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__14801\,
            I => \b2v_inst16.count_4_15\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__14798\,
            I => \b2v_inst16.count_rst_12_cascade_\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__14795\,
            I => \b2v_inst16.count_rst_13_cascade_\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__14792\,
            I => \b2v_inst16.count_rst_14_cascade_\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__14789\,
            I => \b2v_inst16.countZ0Z_9_cascade_\
        );

    \I__1243\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__14783\,
            I => \b2v_inst16.count_4_9\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__14780\,
            I => \b2v_inst16.count_rst_6_cascade_\
        );

    \IN_MUX_bfv_11_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_1_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst6.un2_count_1_cry_8\,
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst5.un2_count_1_cry_7\,
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst36.un2_count_1_cry_7\,
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_8\,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_16\,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => b2v_inst20_un4_counter_7,
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_8\,
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_16\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_24\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst16.un4_count_1_cry_8\,
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un3_count_off_1_cry_8\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_15_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_94_cry_7\,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_cry_8\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \b2v_inst200.count_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17369\,
            GLOBALBUFFEROUTPUT => \b2v_inst200.count_en_g\
        );

    \N_606_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__31250\,
            GLOBALBUFFEROUTPUT => \N_606_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__15679\,
            in1 => \N__17721\,
            in2 => \N__15710\,
            in3 => \N__17565\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNINJ2K1_7_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15410\,
            in1 => \_gnd_net_\,
            in2 => \N__14798\,
            in3 => \N__20093\,
            lcout => \b2v_inst16.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__15634\,
            in1 => \N__17722\,
            in2 => \N__15662\,
            in3 => \N__17566\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14816\,
            in2 => \N__14795\,
            in3 => \N__20094\,
            lcout => \b2v_inst16.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__15612\,
            in1 => \N__17723\,
            in2 => \N__15593\,
            in3 => \N__17567\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIRP4K1_9_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14786\,
            in2 => \N__14792\,
            in3 => \N__20095\,
            lcout => \b2v_inst16.countZ0Z_9\,
            ltout => \b2v_inst16.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_9_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__17729\,
            in1 => \N__17568\,
            in2 => \N__14789\,
            in3 => \N__15592\,
            lcout => \b2v_inst16.count_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36421\,
            ce => \N__20108\,
            sr => \N__17888\
        );

    \b2v_inst16.count_11_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__17542\,
            in1 => \N__15893\,
            in2 => \N__17731\,
            in3 => \N__15909\,
            lcout => \b2v_inst16.count_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36469\,
            ce => \N__20096\,
            sr => \N__17906\
        );

    \b2v_inst16.count_RNI_1_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__15478\,
            in1 => \N__17700\,
            in2 => \_gnd_net_\,
            in3 => \N__15499\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI2J651_1_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14834\,
            in2 => \N__14780\,
            in3 => \N__20085\,
            lcout => \b2v_inst16.countZ0Z_1\,
            ltout => \b2v_inst16.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_1_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17704\,
            in2 => \N__14837\,
            in3 => \N__15500\,
            lcout => \b2v_inst16.count_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36469\,
            ce => \N__20096\,
            sr => \N__17906\
        );

    \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__17541\,
            in1 => \N__15892\,
            in2 => \N__17730\,
            in3 => \N__15910\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIDGU31_11_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__20086\,
            in1 => \N__14828\,
            in2 => \N__14822\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.countZ0Z_11\,
            ltout => \b2v_inst16.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_11_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15657\,
            in1 => \N__15614\,
            in2 => \N__14819\,
            in3 => \N__15477\,
            lcout => \b2v_inst16.count_4_i_a3_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_8_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__17543\,
            in1 => \N__15656\,
            in2 => \N__15635\,
            in3 => \N__17708\,
            lcout => \b2v_inst16.count_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36469\,
            ce => \N__20096\,
            sr => \N__17906\
        );

    \b2v_inst16.count_RNILG1K1_6_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20089\,
            in1 => \N__14810\,
            in2 => \_gnd_net_\,
            in3 => \N__15721\,
            lcout => \b2v_inst16.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_6_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36422\,
            ce => \N__20104\,
            sr => \N__17903\
        );

    \b2v_inst16.count_RNILS241_15_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20105\,
            in1 => \N__15851\,
            in2 => \_gnd_net_\,
            in3 => \N__14804\,
            lcout => \b2v_inst16.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_15_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15850\,
            lcout => \b2v_inst16.count_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36422\,
            ce => \N__20104\,
            sr => \N__17903\
        );

    \b2v_inst16.count_RNI_0_0_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15502\,
            in1 => \N__17699\,
            in2 => \_gnd_net_\,
            in3 => \N__15538\,
            lcout => \b2v_inst16.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_0_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15537\,
            in2 => \_gnd_net_\,
            in3 => \N__15503\,
            lcout => \b2v_inst16.N_416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI1QV41_2_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14885\,
            in1 => \N__16564\,
            in2 => \_gnd_net_\,
            in3 => \N__14960\,
            lcout => \b2v_inst200.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50251_4_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16565\,
            in1 => \N__14876\,
            in2 => \_gnd_net_\,
            in3 => \N__14939\,
            lcout => \b2v_inst200.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9S71_16_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15009\,
            in1 => \N__14860\,
            in2 => \_gnd_net_\,
            in3 => \N__16561\,
            lcout => \b2v_inst200.un2_count_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_16_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15011\,
            lcout => \b2v_inst200.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36401\,
            ce => \N__16485\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNID13N_0_1_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000111"
        )
    port map (
            in0 => \N__14843\,
            in1 => \N__16563\,
            in2 => \N__14900\,
            in3 => \N__14974\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIOAVU1_1_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14849\,
            in1 => \N__16334\,
            in2 => \N__14867\,
            in3 => \N__16105\,
            lcout => \b2v_inst200.un25_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9S71_0_16_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__15010\,
            in1 => \N__15976\,
            in2 => \N__14864\,
            in3 => \N__16562\,
            lcout => \b2v_inst200.un25_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_1_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16104\,
            in2 => \_gnd_net_\,
            in3 => \N__14989\,
            lcout => \b2v_inst200.count_RNIZ0Z_1\,
            ltout => \b2v_inst200.count_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNID13N_1_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14896\,
            in2 => \N__14906\,
            in3 => \N__16560\,
            lcout => \b2v_inst200.un2_count_1_axb_1\,
            ltout => \b2v_inst200.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_1_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14903\,
            in3 => \N__16106\,
            lcout => \b2v_inst200.count_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36401\,
            ce => \N__16485\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_11_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16349\,
            lcout => \b2v_inst200.count_3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36490\,
            ce => \N__16488\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_14_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15833\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36490\,
            ce => \N__16488\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_2_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14959\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36490\,
            ce => \N__16488\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_4_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14938\,
            lcout => \b2v_inst200.count_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36490\,
            ce => \N__16488\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_6_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16040\,
            lcout => \b2v_inst200.count_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36490\,
            ce => \N__16488\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_7_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16022\,
            lcout => \b2v_inst200.count_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36490\,
            ce => \N__16488\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_10_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15964\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36490\,
            ce => \N__16488\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_1_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14990\,
            in2 => \N__16114\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14975\,
            in2 => \_gnd_net_\,
            in3 => \N__14945\,
            lcout => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_1\,
            carryout => \b2v_inst200.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16316\,
            in2 => \_gnd_net_\,
            in3 => \N__14942\,
            lcout => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_2\,
            carryout => \b2v_inst200.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16255\,
            in2 => \_gnd_net_\,
            in3 => \N__14924\,
            lcout => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_3\,
            carryout => \b2v_inst200.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16364\,
            in2 => \_gnd_net_\,
            in3 => \N__14921\,
            lcout => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_4\,
            carryout => \b2v_inst200.un2_count_1_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19437\,
            in1 => \_gnd_net_\,
            in2 => \N__16156\,
            in3 => \N__14918\,
            lcout => \b2v_inst200.count_1_6\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_5_cZ0\,
            carryout => \b2v_inst200.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16591\,
            in3 => \N__14915\,
            lcout => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_6\,
            carryout => \b2v_inst200.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19438\,
            in1 => \N__16193\,
            in2 => \_gnd_net_\,
            in3 => \N__14912\,
            lcout => \b2v_inst200.count_1_8\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_7\,
            carryout => \b2v_inst200.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16073\,
            in2 => \_gnd_net_\,
            in3 => \N__14909\,
            lcout => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19439\,
            in1 => \_gnd_net_\,
            in2 => \N__15929\,
            in3 => \N__15041\,
            lcout => \b2v_inst200.count_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_9\,
            carryout => \b2v_inst200.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19441\,
            in1 => \N__16327\,
            in2 => \_gnd_net_\,
            in3 => \N__15038\,
            lcout => \b2v_inst200.count_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_10\,
            carryout => \b2v_inst200.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16052\,
            in2 => \_gnd_net_\,
            in3 => \N__15035\,
            lcout => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_11\,
            carryout => \b2v_inst200.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16634\,
            in2 => \_gnd_net_\,
            in3 => \N__15032\,
            lcout => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_12\,
            carryout => \b2v_inst200.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16303\,
            in2 => \_gnd_net_\,
            in3 => \N__15029\,
            lcout => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_13\,
            carryout => \b2v_inst200.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16187\,
            in2 => \_gnd_net_\,
            in3 => \N__15026\,
            lcout => \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_14\,
            carryout => \b2v_inst200.un2_count_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19440\,
            in1 => \_gnd_net_\,
            in2 => \N__15023\,
            in3 => \N__14996\,
            lcout => \b2v_inst200.count_1_16\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_15\,
            carryout => \b2v_inst200.un2_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__15980\,
            in1 => \N__19446\,
            in2 => \_gnd_net_\,
            in3 => \N__14993\,
            lcout => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_17_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15994\,
            lcout => \b2v_inst200.count_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36542\,
            ce => \N__16490\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_0_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16115\,
            in2 => \_gnd_net_\,
            in3 => \N__19445\,
            lcout => \b2v_inst200.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21314\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18131\,
            in2 => \N__16738\,
            in3 => \N__15062\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16734\,
            in2 => \N__16430\,
            in3 => \N__15059\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16418\,
            in2 => \N__18157\,
            in3 => \N__15056\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18153\,
            in2 => \N__16409\,
            in3 => \N__15053\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18500\,
            in1 => \N__16397\,
            in2 => \N__16739\,
            in3 => \N__15050\,
            lcout => \b2v_inst11.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16757\,
            in3 => \N__15047\,
            lcout => \b2v_inst11.mult1_un68_sum_s_8\,
            ltout => \b2v_inst11.mult1_un68_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15044\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21346\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16826\,
            in2 => \N__15097\,
            in3 => \N__15140\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15093\,
            in2 => \N__15137\,
            in3 => \N__15128\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15125\,
            in2 => \N__18508\,
            in3 => \N__15119\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18504\,
            in2 => \N__15116\,
            in3 => \N__15107\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16844\,
            in1 => \N__15104\,
            in2 => \N__15098\,
            in3 => \N__15080\,
            lcout => \b2v_inst11.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15077\,
            in3 => \N__15068\,
            lcout => \b2v_inst11.mult1_un75_sum_s_8\,
            ltout => \b2v_inst11.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15065\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21419\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16820\,
            in2 => \N__16801\,
            in3 => \N__15164\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16797\,
            in2 => \N__16721\,
            in3 => \N__15161\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16700\,
            in2 => \N__16784\,
            in3 => \N__15158\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16783\,
            in2 => \N__16685\,
            in3 => \N__15155\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16934\,
            in1 => \N__16664\,
            in2 => \N__16802\,
            in3 => \N__15152\,
            lcout => \b2v_inst11.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16892\,
            in3 => \N__15149\,
            lcout => \b2v_inst11.mult1_un89_sum_s_8\,
            ltout => \b2v_inst11.mult1_un89_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15146\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21455\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16814\,
            in2 => \N__15205\,
            in3 => \N__15143\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15201\,
            in2 => \N__15245\,
            in3 => \N__15236\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15233\,
            in2 => \N__16940\,
            in3 => \N__15227\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16938\,
            in2 => \N__15224\,
            in3 => \N__15215\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17009\,
            in1 => \N__15212\,
            in2 => \N__15206\,
            in3 => \N__15188\,
            lcout => \b2v_inst11.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15185\,
            in3 => \N__15176\,
            lcout => \b2v_inst11.mult1_un96_sum_s_8\,
            ltout => \b2v_inst11.mult1_un96_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15173\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI0AHN_8_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30732\,
            in1 => \N__15170\,
            in2 => \_gnd_net_\,
            in3 => \N__15397\,
            lcout => \b2v_inst11.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_8_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15401\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36580\,
            ce => \N__32182\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI2DIN_9_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30731\,
            in1 => \N__15275\,
            in2 => \_gnd_net_\,
            in3 => \N__15379\,
            lcout => \b2v_inst11.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_9_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15383\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36580\,
            ce => \N__32182\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIB49T_10_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15365\,
            in1 => \N__15269\,
            in2 => \_gnd_net_\,
            in3 => \N__30733\,
            lcout => \b2v_inst11.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_10_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15364\,
            lcout => \b2v_inst11.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36580\,
            ce => \N__32182\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIK61M_11_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15350\,
            in1 => \N__15263\,
            in2 => \_gnd_net_\,
            in3 => \N__30734\,
            lcout => \b2v_inst11.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_11_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15349\,
            lcout => \b2v_inst11.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36580\,
            ce => \N__32182\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_1_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__18432\,
            in1 => \N__18471\,
            in2 => \_gnd_net_\,
            in3 => \N__17109\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI14G9_1_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30729\,
            in1 => \_gnd_net_\,
            in2 => \N__15257\,
            in3 => \N__15251\,
            lcout => \b2v_inst11.countZ0Z_1\,
            ltout => \b2v_inst11.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_1_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18473\,
            in2 => \N__15254\,
            in3 => \N__17113\,
            lcout => \b2v_inst11.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__32181\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_0_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__18472\,
            in1 => \_gnd_net_\,
            in2 => \N__17142\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__32181\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIKNAN_2_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15314\,
            in2 => \N__15302\,
            in3 => \N__30728\,
            lcout => \b2v_inst11.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_2_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15301\,
            lcout => \b2v_inst11.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__32181\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIM92M_12_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15335\,
            in1 => \N__15308\,
            in2 => \_gnd_net_\,
            in3 => \N__30730\,
            lcout => \b2v_inst11.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_12_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15334\,
            lcout => \b2v_inst11.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__32181\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18478\,
            in2 => \N__18433\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \b2v_inst11.un1_count_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__17146\,
            in1 => \_gnd_net_\,
            in2 => \N__18394\,
            in3 => \N__15290\,
            lcout => \b2v_inst11.count_1_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_1_cZ0\,
            carryout => \b2v_inst11.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17139\,
            in1 => \N__18354\,
            in2 => \_gnd_net_\,
            in3 => \N__15287\,
            lcout => \b2v_inst11.count_1_3\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_2\,
            carryout => \b2v_inst11.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17143\,
            in1 => \N__18319\,
            in2 => \_gnd_net_\,
            in3 => \N__15284\,
            lcout => \b2v_inst11.count_1_4\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_3\,
            carryout => \b2v_inst11.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17140\,
            in1 => \N__18286\,
            in2 => \_gnd_net_\,
            in3 => \N__15281\,
            lcout => \b2v_inst11.count_1_5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_4\,
            carryout => \b2v_inst11.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17144\,
            in1 => \N__18847\,
            in2 => \_gnd_net_\,
            in3 => \N__15278\,
            lcout => \b2v_inst11.count_1_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_5\,
            carryout => \b2v_inst11.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17141\,
            in1 => \N__18814\,
            in2 => \_gnd_net_\,
            in3 => \N__15404\,
            lcout => \b2v_inst11.count_1_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_6\,
            carryout => \b2v_inst11.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__18787\,
            in2 => \_gnd_net_\,
            in3 => \N__15386\,
            lcout => \b2v_inst11.count_1_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_7\,
            carryout => \b2v_inst11.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17147\,
            in1 => \N__18748\,
            in2 => \_gnd_net_\,
            in3 => \N__15368\,
            lcout => \b2v_inst11.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \b2v_inst11.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17152\,
            in1 => \N__18699\,
            in2 => \_gnd_net_\,
            in3 => \N__15353\,
            lcout => \b2v_inst11.count_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_9\,
            carryout => \b2v_inst11.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17148\,
            in1 => \N__18651\,
            in2 => \_gnd_net_\,
            in3 => \N__15338\,
            lcout => \b2v_inst11.count_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_10\,
            carryout => \b2v_inst11.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17151\,
            in1 => \N__18615\,
            in2 => \_gnd_net_\,
            in3 => \N__15323\,
            lcout => \b2v_inst11.count_1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_11\,
            carryout => \b2v_inst11.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17149\,
            in1 => \N__18556\,
            in2 => \_gnd_net_\,
            in3 => \N__15320\,
            lcout => \b2v_inst11.count_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_12\,
            carryout => \b2v_inst11.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17153\,
            in1 => \N__18970\,
            in2 => \_gnd_net_\,
            in3 => \N__15317\,
            lcout => \b2v_inst11.count_1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_13\,
            carryout => \b2v_inst11.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17150\,
            in1 => \N__18934\,
            in2 => \_gnd_net_\,
            in3 => \N__15437\,
            lcout => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__17571\,
            in1 => \N__15784\,
            in2 => \N__15812\,
            in3 => \N__17713\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIHAVJ1_4_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15428\,
            in2 => \N__15434\,
            in3 => \N__20087\,
            lcout => \b2v_inst16.countZ0Z_4\,
            ltout => \b2v_inst16.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_4_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17575\,
            in1 => \N__17716\,
            in2 => \N__15431\,
            in3 => \N__15785\,
            lcout => \b2v_inst16.count_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36420\,
            ce => \N__20106\,
            sr => \N__17899\
        );

    \b2v_inst16.count_3_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__17715\,
            in1 => \N__17577\,
            in2 => \N__17489\,
            in3 => \N__17822\,
            lcout => \b2v_inst16.count_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36420\,
            ce => \N__20106\,
            sr => \N__17899\
        );

    \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__15768\,
            in1 => \N__17714\,
            in2 => \N__17579\,
            in3 => \N__15748\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15416\,
            in2 => \N__15422\,
            in3 => \N__20088\,
            lcout => \b2v_inst16.countZ0Z_5\,
            ltout => \b2v_inst16.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_5_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17576\,
            in1 => \N__17717\,
            in2 => \N__15419\,
            in3 => \N__15749\,
            lcout => \b2v_inst16.count_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36420\,
            ce => \N__20106\,
            sr => \N__17899\
        );

    \b2v_inst16.count_7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__17578\,
            in1 => \N__15704\,
            in2 => \N__17732\,
            in3 => \N__15680\,
            lcout => \b2v_inst16.count_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36420\,
            ce => \N__20106\,
            sr => \N__17899\
        );

    \b2v_inst16.count_2_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__17711\,
            in1 => \N__15447\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36468\,
            ce => \N__20038\,
            sr => \N__17904\
        );

    \b2v_inst16.count_RNID4TJ1_2_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15451\,
            in1 => \N__17712\,
            in2 => \N__15515\,
            in3 => \N__20039\,
            lcout => OPEN,
            ltout => \b2v_inst16.countZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNID4TJ1_2_2_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19958\,
            in1 => \N__15865\,
            in2 => \N__15566\,
            in3 => \N__15734\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_4_i_a3_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI2T6K2_13_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15554\,
            in1 => \N__15563\,
            in2 => \N__15557\,
            in3 => \N__17465\,
            lcout => \b2v_inst16.N_414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_4_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15769\,
            in1 => \N__15808\,
            in2 => \_gnd_net_\,
            in3 => \N__15708\,
            lcout => \b2v_inst16.count_4_i_a3_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI1I651_0_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15548\,
            in1 => \N__15521\,
            in2 => \_gnd_net_\,
            in3 => \N__20036\,
            lcout => \b2v_inst16.countZ0Z_0\,
            ltout => \b2v_inst16.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_0_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__17710\,
            in1 => \_gnd_net_\,
            in2 => \N__15542\,
            in3 => \N__15539\,
            lcout => \b2v_inst16.count_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36468\,
            ce => \N__20038\,
            sr => \N__17904\
        );

    \b2v_inst16.count_RNID4TJ1_0_2_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__15511\,
            in1 => \N__17709\,
            in2 => \N__15452\,
            in3 => \N__20037\,
            lcout => \b2v_inst16.un4_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_1_c_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15501\,
            in2 => \N__15479\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15461\,
            in3 => \N__15818\,
            lcout => \b2v_inst16.un4_count_1_cry_1_c_RNIAGMEZ0\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_1\,
            carryout => \b2v_inst16.un4_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17821\,
            in2 => \_gnd_net_\,
            in3 => \N__15815\,
            lcout => \b2v_inst16.un4_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_2\,
            carryout => \b2v_inst16.un4_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15807\,
            in2 => \_gnd_net_\,
            in3 => \N__15773\,
            lcout => \b2v_inst16.un4_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_3\,
            carryout => \b2v_inst16.un4_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15770\,
            in2 => \_gnd_net_\,
            in3 => \N__15737\,
            lcout => \b2v_inst16.un4_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_4\,
            carryout => \b2v_inst16.un4_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17682\,
            in1 => \N__15733\,
            in2 => \_gnd_net_\,
            in3 => \N__15713\,
            lcout => \b2v_inst16.count_rst_11\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_5\,
            carryout => \b2v_inst16.un4_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15709\,
            in2 => \_gnd_net_\,
            in3 => \N__15665\,
            lcout => \b2v_inst16.un4_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_6\,
            carryout => \b2v_inst16.un4_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15661\,
            in2 => \_gnd_net_\,
            in3 => \N__15617\,
            lcout => \b2v_inst16.un4_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_7\,
            carryout => \b2v_inst16.un4_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15613\,
            in2 => \_gnd_net_\,
            in3 => \N__15572\,
            lcout => \b2v_inst16.un4_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_4_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17727\,
            in1 => \N__19954\,
            in2 => \_gnd_net_\,
            in3 => \N__15569\,
            lcout => \b2v_inst16.count_rst\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_9\,
            carryout => \b2v_inst16.un4_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15911\,
            in2 => \_gnd_net_\,
            in3 => \N__15881\,
            lcout => \b2v_inst16.un4_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_10\,
            carryout => \b2v_inst16.un4_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17724\,
            in1 => \N__17420\,
            in2 => \_gnd_net_\,
            in3 => \N__15878\,
            lcout => \b2v_inst16.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_11\,
            carryout => \b2v_inst16.un4_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_12_c_RNIHM041_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17728\,
            in1 => \N__17941\,
            in2 => \_gnd_net_\,
            in3 => \N__15875\,
            lcout => \b2v_inst16.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_12\,
            carryout => \b2v_inst16.un4_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17725\,
            in1 => \N__17453\,
            in2 => \_gnd_net_\,
            in3 => \N__15872\,
            lcout => \b2v_inst16.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_13\,
            carryout => \b2v_inst16.un4_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__15869\,
            in1 => \N__17726\,
            in2 => \_gnd_net_\,
            in3 => \N__15854\,
            lcout => \b2v_inst16.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_10_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20134\,
            lcout => \b2v_inst16.count_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36619\,
            ce => \N__20103\,
            sr => \N__17905\
        );

    \b2v_inst16.curr_state_1_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__27735\,
            in1 => \N__17564\,
            in2 => \_gnd_net_\,
            in3 => \N__27770\,
            lcout => \b2v_inst16.curr_state_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36438\,
            ce => \N__32177\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__33576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27736\,
            lcout => \b2v_inst16.curr_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36438\,
            ce => \N__32177\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73Q71_14_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16558\,
            in1 => \N__15839\,
            in2 => \_gnd_net_\,
            in3 => \N__15832\,
            lcout => \b2v_inst200.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI96451_6_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16046\,
            in1 => \N__16039\,
            in2 => \_gnd_net_\,
            in3 => \N__16555\,
            lcout => \b2v_inst200.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9551_7_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16556\,
            in1 => \N__16028\,
            in2 => \_gnd_net_\,
            in3 => \N__16021\,
            lcout => \b2v_inst200.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDCT71_17_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16010\,
            in1 => \N__15998\,
            in2 => \_gnd_net_\,
            in3 => \N__16559\,
            lcout => \b2v_inst200.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIOMPC1_10_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16557\,
            in1 => \_gnd_net_\,
            in2 => \N__15965\,
            in3 => \N__15947\,
            lcout => \b2v_inst200.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_0_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16079\,
            in1 => \N__16554\,
            in2 => \_gnd_net_\,
            in3 => \N__15938\,
            lcout => \b2v_inst200.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_8_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16217\,
            lcout => \b2v_inst200.count_3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36470\,
            ce => \N__16486\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_15_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16171\,
            lcout => \b2v_inst200.count_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36470\,
            ce => \N__16486\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDC651_0_8_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__16573\,
            in1 => \N__15925\,
            in2 => \N__16205\,
            in3 => \N__16216\,
            lcout => \b2v_inst200.un25_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDC651_8_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16215\,
            in1 => \N__16201\,
            in2 => \_gnd_net_\,
            in3 => \N__16571\,
            lcout => \b2v_inst200.un2_count_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI2KKU_15_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16572\,
            in1 => \_gnd_net_\,
            in2 => \N__16172\,
            in3 => \N__16180\,
            lcout => \b2v_inst200.un2_count_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI2KKU_0_15_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001010000"
        )
    port map (
            in0 => \N__16181\,
            in1 => \N__16170\,
            in2 => \N__16157\,
            in3 => \N__16574\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI5RUP8_8_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16139\,
            in1 => \N__16133\,
            in2 => \N__16121\,
            in3 => \N__16280\,
            lcout => \b2v_inst200.count_RNI5RUP8Z0Z_8\,
            ltout => \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16118\,
            in3 => \N__16110\,
            lcout => \b2v_inst200.count_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36470\,
            ce => \N__16486\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_12_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16061\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36491\,
            ce => \N__16487\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_9_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36491\,
            ce => \N__16487\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIFF751_9_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16567\,
            in1 => \N__16387\,
            in2 => \_gnd_net_\,
            in3 => \N__16374\,
            lcout => \b2v_inst200.un2_count_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3TN71_12_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16067\,
            in1 => \N__16060\,
            in2 => \_gnd_net_\,
            in3 => \N__16569\,
            lcout => \b2v_inst200.countZ0Z_12\,
            ltout => \b2v_inst200.countZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIFF751_0_9_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__16570\,
            in1 => \N__16388\,
            in2 => \N__16379\,
            in3 => \N__16376\,
            lcout => \b2v_inst200.un25_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73351_5_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16607\,
            in1 => \N__16566\,
            in2 => \_gnd_net_\,
            in3 => \N__16620\,
            lcout => \b2v_inst200.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_5_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36491\,
            ce => \N__16487\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI1QM71_11_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16358\,
            in1 => \N__16345\,
            in2 => \_gnd_net_\,
            in3 => \N__16568\,
            lcout => \b2v_inst200.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3T051_3_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16550\,
            in1 => \N__16270\,
            in2 => \_gnd_net_\,
            in3 => \N__16236\,
            lcout => \b2v_inst200.un2_count_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_3_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36531\,
            ce => \N__16489\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50P71_0_13_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__16553\,
            in1 => \N__16655\,
            in2 => \N__16307\,
            in3 => \N__16646\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIUF4N4_3_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16289\,
            in1 => \N__16223\,
            in2 => \N__16283\,
            in3 => \N__16436\,
            lcout => \b2v_inst200.un25_clk_100khz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3T051_0_3_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__16552\,
            in1 => \N__16271\,
            in2 => \N__16262\,
            in3 => \N__16238\,
            lcout => \b2v_inst200.un25_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_13_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16645\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36531\,
            ce => \N__16489\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50P71_13_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16551\,
            in1 => \N__16654\,
            in2 => \_gnd_net_\,
            in3 => \N__16644\,
            lcout => \b2v_inst200.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73351_0_5_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__16628\,
            in1 => \N__16606\,
            in2 => \N__16595\,
            in3 => \N__16549\,
            lcout => \b2v_inst200.un25_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21275\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18173\,
            in2 => \N__16867\,
            in3 => \N__16421\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16863\,
            in2 => \N__18098\,
            in3 => \N__16412\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18083\,
            in2 => \N__18245\,
            in3 => \N__16400\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18243\,
            in2 => \N__18071\,
            in3 => \N__16391\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18149\,
            in1 => \N__18056\,
            in2 => \N__16868\,
            in3 => \N__16748\,
            lcout => \b2v_inst11.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18260\,
            in2 => \_gnd_net_\,
            in3 => \N__16745\,
            lcout => \b2v_inst11.mult1_un61_sum_s_8\,
            ltout => \b2v_inst11.mult1_un61_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16742\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21379\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18521\,
            in2 => \N__16909\,
            in3 => \N__16712\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16905\,
            in2 => \N__16709\,
            in3 => \N__16694\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16691\,
            in2 => \N__16850\,
            in3 => \N__16676\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16848\,
            in2 => \N__16673\,
            in3 => \N__16658\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16779\,
            in1 => \N__16916\,
            in2 => \N__16910\,
            in3 => \N__16883\,
            lcout => \b2v_inst11.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16880\,
            in3 => \N__16871\,
            lcout => \b2v_inst11.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18244\,
            lcout => \b2v_inst11.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16849\,
            lcout => \b2v_inst11.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21313\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21383\,
            lcout => \b2v_inst11.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21418\,
            lcout => \b2v_inst11.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16777\,
            lcout => \b2v_inst11.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un82_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17014\,
            lcout => \b2v_inst11.mult1_un96_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21496\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20267\,
            in2 => \N__16972\,
            in3 => \N__17039\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16968\,
            in2 => \N__17036\,
            in3 => \N__17027\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17024\,
            in2 => \N__17015\,
            in3 => \N__17018\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17013\,
            in2 => \N__16991\,
            in3 => \N__16982\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20225\,
            in1 => \N__16979\,
            in2 => \N__16973\,
            in3 => \N__16955\,
            lcout => \b2v_inst11.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16952\,
            in3 => \N__16943\,
            lcout => \b2v_inst11.mult1_un103_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16939\,
            lcout => \b2v_inst11.mult1_un89_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNI2EHH1_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__17063\,
            in1 => \N__19812\,
            in2 => \N__17054\,
            in3 => \N__17294\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19841\,
            in2 => \N__19816\,
            in3 => \N__19779\,
            lcout => OPEN,
            ltout => \b2v_inst11.curr_state_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIJK34_0_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19754\,
            in2 => \N__17159\,
            in3 => \N__30577\,
            lcout => \b2v_inst11.curr_stateZ0Z_0\,
            ltout => \b2v_inst11.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIOCA3_0_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__30578\,
            in1 => \_gnd_net_\,
            in2 => \N__17156\,
            in3 => \N__19778\,
            lcout => \b2v_inst11.count_0_sqmuxa_i\,
            ltout => \b2v_inst11.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_0_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__18474\,
            in1 => \_gnd_net_\,
            in2 => \N__17075\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI03G9_0_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30579\,
            in1 => \_gnd_net_\,
            in2 => \N__17072\,
            in3 => \N__17069\,
            lcout => \b2v_inst11.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__17062\,
            in1 => \N__19811\,
            in2 => \N__17053\,
            in3 => \N__17293\,
            lcout => \b2v_inst11.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36575\,
            ce => 'H',
            sr => \N__17177\
        );

    \b2v_inst11.curr_state_RNIKEBL_0_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32223\,
            in2 => \_gnd_net_\,
            in3 => \N__19840\,
            lcout => \b2v_inst11.g0_i_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIMQBN_3_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30693\,
            in1 => \N__17237\,
            in2 => \_gnd_net_\,
            in3 => \N__17245\,
            lcout => \b2v_inst11.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_3_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17249\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36581\,
            ce => \N__32180\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOC3M_13_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__17231\,
            in1 => \N__17219\,
            in2 => \N__30726\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_13_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17230\,
            lcout => \b2v_inst11.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36581\,
            ce => \N__32180\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOTCN_4_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30692\,
            in1 => \N__17201\,
            in2 => \_gnd_net_\,
            in3 => \N__17209\,
            lcout => \b2v_inst11.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_4_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17213\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36581\,
            ce => \N__32180\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQ0EN_5_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30694\,
            in1 => \N__17183\,
            in2 => \_gnd_net_\,
            in3 => \N__17191\,
            lcout => \b2v_inst11.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_5_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17195\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36581\,
            ce => \N__32180\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNO_0_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19846\,
            in2 => \N__19783\,
            in3 => \N__30700\,
            lcout => \b2v_inst11.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_2_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18318\,
            in2 => \N__18358\,
            in3 => \N__18387\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_5_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__18285\,
            in1 => \N__18846\,
            in2 => \N__17312\,
            in3 => \N__18813\,
            lcout => \b2v_inst11.un79_clk_100khzlto15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_10_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18703\,
            in1 => \N__18543\,
            in2 => \N__18616\,
            in3 => \N__18659\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_15_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__18969\,
            in1 => \_gnd_net_\,
            in2 => \N__17309\,
            in3 => \N__18933\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_8_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18747\,
            in1 => \N__18786\,
            in2 => \N__17306\,
            in3 => \N__17303\,
            lcout => \b2v_inst11.count_RNIZ0Z_8\,
            ltout => \b2v_inst11.count_RNIZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNICRLO_0_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30701\,
            in1 => \N__32222\,
            in2 => \N__17297\,
            in3 => \N__19845\,
            lcout => \b2v_inst11.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQF4M_14_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17282\,
            in1 => \N__17273\,
            in2 => \_gnd_net_\,
            in3 => \N__30691\,
            lcout => \b2v_inst11.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_14_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17281\,
            lcout => \b2v_inst11.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36602\,
            ce => \N__32179\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIS3FN_6_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30698\,
            in1 => \N__17255\,
            in2 => \_gnd_net_\,
            in3 => \N__17263\,
            lcout => \b2v_inst11.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_6_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17267\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36602\,
            ce => \N__32179\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNISI5M_15_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17393\,
            in1 => \N__30690\,
            in2 => \_gnd_net_\,
            in3 => \N__17401\,
            lcout => \b2v_inst11.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_15_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17405\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36602\,
            ce => \N__32179\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIU6GN_7_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30699\,
            in1 => \N__17375\,
            in2 => \_gnd_net_\,
            in3 => \N__17383\,
            lcout => \b2v_inst11.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_7_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17387\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36602\,
            ce => \N__32179\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19482\,
            in2 => \_gnd_net_\,
            in3 => \N__19461\,
            lcout => \b2v_inst200.N_282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI_0_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17698\,
            lcout => \b2v_inst16.N_3079_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_en_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19481\,
            in2 => \_gnd_net_\,
            in3 => \N__32219\,
            lcout => \b2v_inst200.count_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIKEBL_1_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__17614\,
            in1 => \N__27720\,
            in2 => \_gnd_net_\,
            in3 => \N__32220\,
            lcout => \b2v_inst16.count_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_0_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29492\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIUCAD1_1_0_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27721\,
            in1 => \N__17569\,
            in2 => \_gnd_net_\,
            in3 => \N__27759\,
            lcout => \b2v_inst16.curr_state_7_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.delayed_vddq_pwrgd_e_0_RNI8HF43_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__17744\,
            in1 => \N__17750\,
            in2 => \N__27734\,
            in3 => \N__33653\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.delayed_vddq_pwrgd_e_0_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011111111"
        )
    port map (
            in0 => \N__19520\,
            in1 => \N__27722\,
            in2 => \N__30689\,
            in3 => \N__33578\,
            lcout => \b2v_inst16.delayed_vddq_pwrgd_eZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36208\,
            ce => \N__17743\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIIRL22_0_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32221\,
            lcout => \b2v_inst16.delayed_vddq_pwrgd_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIMPKG1_0_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27688\,
            in2 => \_gnd_net_\,
            in3 => \N__30627\,
            lcout => \b2v_inst16.N_26\,
            ltout => \b2v_inst16.N_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__17570\,
            in1 => \N__17488\,
            in2 => \N__17468\,
            in3 => \N__17814\,
            lcout => \b2v_inst16.count_rst_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNILO901_0_13_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__17419\,
            in1 => \N__17452\,
            in2 => \N__17942\,
            in3 => \N__17807\,
            lcout => \b2v_inst16.count_4_i_a3_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIJP141_14_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17426\,
            in1 => \N__20077\,
            in2 => \_gnd_net_\,
            in3 => \N__17437\,
            lcout => \b2v_inst16.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_14_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17438\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36291\,
            ce => \N__20078\,
            sr => \N__17892\
        );

    \b2v_inst16.count_RNIFJV31_12_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17948\,
            in1 => \N__20075\,
            in2 => \_gnd_net_\,
            in3 => \N__17959\,
            lcout => \b2v_inst16.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_12_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36291\,
            ce => \N__20078\,
            sr => \N__17892\
        );

    \b2v_inst16.count_RNILO901_13_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17912\,
            in1 => \N__20076\,
            in2 => \_gnd_net_\,
            in3 => \N__17923\,
            lcout => \b2v_inst16.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_13_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36291\,
            ce => \N__20078\,
            sr => \N__17892\
        );

    \b2v_inst16.count_RNIF7UJ1_3_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17840\,
            in1 => \N__20079\,
            in2 => \_gnd_net_\,
            in3 => \N__17828\,
            lcout => \b2v_inst16.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_7_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__33884\,
            in1 => \N__25346\,
            in2 => \N__22841\,
            in3 => \N__17786\,
            lcout => \b2v_inst11.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36314\,
            ce => 'H',
            sr => \N__31031\
        );

    \b2v_inst11.dutycycle_RNIRH7VD_7_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__17785\,
            in1 => \N__33883\,
            in2 => \N__22840\,
            in3 => \N__25345\,
            lcout => \b2v_inst11.dutycycleZ1Z_3\,
            ltout => \b2v_inst11.dutycycleZ1Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_7_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17777\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_7Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_7_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22631\,
            in2 => \_gnd_net_\,
            in3 => \N__22877\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011010010"
        )
    port map (
            in0 => \N__29972\,
            in1 => \N__22775\,
            in2 => \N__17774\,
            in3 => \N__19715\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_3_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20330\,
            in1 => \N__23437\,
            in2 => \N__30185\,
            in3 => \N__24629\,
            lcout => \b2v_inst11.g3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIN8NR1_1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__17996\,
            in1 => \N__17984\,
            in2 => \_gnd_net_\,
            in3 => \N__30631\,
            lcout => \b2v_inst16.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_10_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22769\,
            in2 => \N__22659\,
            in3 => \N__23563\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_44_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_6_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__19538\,
            in1 => \N__18035\,
            in2 => \N__17972\,
            in3 => \N__29968\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_11_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_13_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22635\,
            in1 => \N__24955\,
            in2 => \N__23099\,
            in3 => \N__23564\,
            lcout => \b2v_inst11.un2_count_clk_17_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_6_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22768\,
            in1 => \N__25414\,
            in2 => \_gnd_net_\,
            in3 => \N__29967\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__25415\,
            in1 => \N__23436\,
            in2 => \_gnd_net_\,
            in3 => \N__24628\,
            lcout => \b2v_inst11.N_355\,
            ltout => \b2v_inst11.N_355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_15_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__22770\,
            in1 => \N__17969\,
            in2 => \N__17963\,
            in3 => \N__24712\,
            lcout => \b2v_inst11.N_363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_8_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001111"
        )
    port map (
            in0 => \N__24598\,
            in1 => \N__25422\,
            in2 => \N__25140\,
            in3 => \N__23572\,
            lcout => \b2v_inst11.un1_dutycycle_53_55_1_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_11_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101011111"
        )
    port map (
            in0 => \N__25080\,
            in1 => \N__22779\,
            in2 => \N__22658\,
            in3 => \N__25216\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_6Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_8_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__19721\,
            in1 => \N__18044\,
            in2 => \N__18038\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_10_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24597\,
            in2 => \N__22657\,
            in3 => \N__23571\,
            lcout => \b2v_inst11.un1_dutycycle_53_50_a0_1\,
            ltout => \b2v_inst11.un1_dutycycle_53_50_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_6_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__22780\,
            in1 => \N__29965\,
            in2 => \N__18029\,
            in3 => \N__18116\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_6_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000100"
        )
    port map (
            in0 => \N__19636\,
            in1 => \N__19616\,
            in2 => \N__18026\,
            in3 => \N__24644\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_12_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23573\,
            in2 => \N__22665\,
            in3 => \N__25085\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_12\,
            ltout => \b2v_inst11.dutycycle_RNI_1Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_6_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__19651\,
            in1 => \N__18020\,
            in2 => \N__18023\,
            in3 => \N__18005\,
            lcout => \b2v_inst11.dutycycle_RNI_8Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_6_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__29961\,
            in1 => \N__24630\,
            in2 => \_gnd_net_\,
            in3 => \N__25426\,
            lcout => \b2v_inst11.un1_dutycycle_53_4_1\,
            ltout => \b2v_inst11.un1_dutycycle_53_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_6_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18014\,
            in2 => \N__18008\,
            in3 => \N__18004\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_7Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_13_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000111100"
        )
    port map (
            in0 => \N__24956\,
            in1 => \N__25086\,
            in2 => \N__18119\,
            in3 => \N__19652\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_7_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__25425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25139\,
            lcout => \b2v_inst11.dutycycle_RNI_9Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_11_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22666\,
            in3 => \N__25217\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_46_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_14_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011110000"
        )
    port map (
            in0 => \N__23091\,
            in1 => \N__19661\,
            in2 => \N__18110\,
            in3 => \N__18107\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21236\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19868\,
            in3 => \N__18086\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19696\,
            in2 => \N__18212\,
            in3 => \N__18074\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32052\,
            in2 => \N__19901\,
            in3 => \N__18059\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19889\,
            in2 => \N__32059\,
            in3 => \N__18047\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18231\,
            in1 => \N__20171\,
            in2 => \N__19877\,
            in3 => \N__18251\,
            lcout => \b2v_inst11.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20183\,
            in2 => \N__20195\,
            in3 => \N__18248\,
            lcout => \b2v_inst11.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__19695\,
            in1 => \N__19697\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un1_vddq_en_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33646\,
            in2 => \_gnd_net_\,
            in3 => \N__18203\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21497\,
            lcout => \b2v_inst11.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21232\,
            lcout => \b2v_inst11.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18161\,
            lcout => \b2v_inst11.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21274\,
            lcout => \b2v_inst11.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_5_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35182\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21347\,
            lcout => \b2v_inst11.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18512\,
            lcout => \b2v_inst11.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18482\,
            in1 => \N__18443\,
            in2 => \N__19223\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5980_i\,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18407\,
            in2 => \N__20276\,
            in3 => \N__18437\,
            lcout => \b2v_inst11.N_5981_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_0\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20282\,
            in2 => \N__18371\,
            in3 => \N__18401\,
            lcout => \b2v_inst11.N_5982_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_1\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18362\,
            in1 => \N__20252\,
            in2 => \N__18335\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5983_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_2\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18326\,
            in1 => \N__19907\,
            in2 => \N__18302\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5984_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_3\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18293\,
            in1 => \N__20258\,
            in2 => \N__18269\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5985_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_4\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18830\,
            in2 => \N__20291\,
            in3 => \N__18857\,
            lcout => \b2v_inst11.N_5986_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_5\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18824\,
            in1 => \N__18797\,
            in2 => \N__19925\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5987_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_6\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18896\,
            in2 => \N__18761\,
            in3 => \N__18791\,
            lcout => \b2v_inst11.N_5988_i\,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20201\,
            in2 => \N__18728\,
            in3 => \N__18752\,
            lcout => \b2v_inst11.N_5989_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_8\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18719\,
            in2 => \N__18677\,
            in3 => \N__18707\,
            lcout => \b2v_inst11.N_5990_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_9\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18668\,
            in2 => \N__18629\,
            in3 => \N__18658\,
            lcout => \b2v_inst11.N_5991_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_10\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18620\,
            in1 => \N__18590\,
            in2 => \N__18578\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5992_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_11\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18569\,
            in2 => \N__18530\,
            in3 => \N__18557\,
            lcout => \b2v_inst11.N_5993_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_12\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18986\,
            in2 => \N__18953\,
            in3 => \N__18977\,
            lcout => \b2v_inst11.N_5994_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_13\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18941\,
            in1 => \N__18917\,
            in2 => \N__18908\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5995_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_14\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18899\,
            lcout => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20241\,
            lcout => \b2v_inst11.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19174\,
            lcout => \b2v_inst11.mult1_un110_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21110\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18890\,
            in2 => \N__19051\,
            in3 => \N__18878\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19047\,
            in2 => \N__18875\,
            in3 => \N__18860\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19097\,
            in2 => \N__20246\,
            in3 => \N__19085\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20245\,
            in2 => \N__19082\,
            in3 => \N__19067\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19169\,
            in1 => \N__19064\,
            in2 => \N__19052\,
            in3 => \N__19034\,
            lcout => \b2v_inst11.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19031\,
            in3 => \N__19016\,
            lcout => \b2v_inst11.mult1_un110_sum_s_8\,
            ltout => \b2v_inst11.mult1_un110_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19013\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21140\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19937\,
            in2 => \N__19132\,
            in3 => \N__19010\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19128\,
            in2 => \N__19007\,
            in3 => \N__18998\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18995\,
            in2 => \N__19175\,
            in3 => \N__18989\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19173\,
            in2 => \N__19151\,
            in3 => \N__19142\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20432\,
            in1 => \N__19139\,
            in2 => \N__19133\,
            in3 => \N__19115\,
            lcout => \b2v_inst11.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19112\,
            in3 => \N__19103\,
            lcout => \b2v_inst11.mult1_un117_sum_s_8\,
            ltout => \b2v_inst11.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19100\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30183\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20498\,
            in2 => \N__19243\,
            in3 => \N__20530\,
            lcout => \G_2814\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_0\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19239\,
            in2 => \N__20597\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20531\,
            in2 => \N__20585\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20573\,
            in2 => \N__20539\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20564\,
            in2 => \N__19244\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20555\,
            in3 => \N__19226\,
            lcout => \b2v_inst11.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__19484\,
            in1 => \N__19463\,
            in2 => \_gnd_net_\,
            in3 => \N__19181\,
            lcout => OPEN,
            ltout => \b2v_inst200.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNILNOU4_0_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19397\,
            in2 => \N__19211\,
            in3 => \N__30575\,
            lcout => \b2v_inst200.curr_stateZ0Z_0\,
            ltout => \b2v_inst200.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19208\,
            in3 => \N__19361\,
            lcout => \N_411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNIMK8L4_1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19250\,
            in1 => \N__19202\,
            in2 => \_gnd_net_\,
            in3 => \N__30576\,
            lcout => \b2v_inst200.curr_stateZ0Z_1\,
            ltout => \b2v_inst200.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI_1_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19205\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.N_3031_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__29488\,
            in1 => \N__19310\,
            in2 => \N__19273\,
            in3 => \N__19294\,
            lcout => \b2v_inst200.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010011101"
        )
    port map (
            in0 => \N__19311\,
            in1 => \N__19290\,
            in2 => \N__19196\,
            in3 => \N__29487\,
            lcout => \b2v_inst200.m6_i_0\,
            ltout => \b2v_inst200.m6_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_0_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19483\,
            in2 => \N__19466\,
            in3 => \N__19462\,
            lcout => \b2v_inst200.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36209\,
            ce => \N__32173\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_2_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000110011"
        )
    port map (
            in0 => \N__29491\,
            in1 => \N__19271\,
            in2 => \N__19349\,
            in3 => \N__19332\,
            lcout => \b2v_inst200.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36368\,
            ce => \N__32175\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__19334\,
            in1 => \N__19344\,
            in2 => \N__19274\,
            in3 => \N__29489\,
            lcout => OPEN,
            ltout => \b2v_inst200.i4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNINL8L4_2_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19391\,
            in2 => \N__19385\,
            in3 => \N__30632\,
            lcout => \b2v_inst200.curr_state_i_2\,
            ltout => \b2v_inst200.curr_state_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__30633\,
            in1 => \N__19319\,
            in2 => \N__19382\,
            in3 => \N__19348\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI_0_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19312\,
            in2 => \_gnd_net_\,
            in3 => \N__19360\,
            lcout => \b2v_inst200.N_205\,
            ltout => \b2v_inst200.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_ATP_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__19333\,
            in1 => \_gnd_net_\,
            in2 => \N__19322\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.HDA_SDO_ATP_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36368\,
            ce => \N__32175\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_1_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__29490\,
            in1 => \N__19313\,
            in2 => \N__19295\,
            in3 => \N__19272\,
            lcout => \b2v_inst200.curr_state_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36368\,
            ce => \N__32175\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_RNO_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20770\,
            in1 => \N__20611\,
            in2 => \N__20789\,
            in3 => \N__20626\,
            lcout => \b2v_inst20.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_RNO_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20707\,
            in1 => \N__20740\,
            in2 => \N__20726\,
            in3 => \N__20755\,
            lcout => \b2v_inst20.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_RNO_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20692\,
            in1 => \N__20659\,
            in2 => \N__20678\,
            in3 => \N__20911\,
            lcout => \b2v_inst20.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_RNO_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20878\,
            in1 => \N__20848\,
            in2 => \N__20897\,
            in3 => \N__20863\,
            lcout => \b2v_inst20.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_0_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__28178\,
            in1 => \N__28130\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIUCAD1_0_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__19519\,
            in1 => \N__33577\,
            in2 => \_gnd_net_\,
            in3 => \N__30543\,
            lcout => \b2v_inst16.curr_state_RNIUCAD1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22334\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => \b2v_inst20.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_1_c_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22220\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_0\,
            carryout => \b2v_inst20.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19496\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_1\,
            carryout => \b2v_inst20.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19490\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_2\,
            carryout => \b2v_inst20.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19553\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_3\,
            carryout => \b2v_inst20.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19547\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_4\,
            carryout => \b2v_inst20.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19604\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_5\,
            carryout => \b2v_inst20.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20927\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_6\,
            carryout => b2v_inst20_un4_counter_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19541\,
            lcout => \b2v_inst20_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__23545\,
            in1 => \N__22777\,
            in2 => \N__25449\,
            in3 => \N__24620\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_39_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_7_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__19537\,
            in1 => \N__19598\,
            in2 => \N__19526\,
            in3 => \N__22908\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_13_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22642\,
            in1 => \N__24943\,
            in2 => \N__19523\,
            in3 => \N__22778\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_10_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19610\,
            in2 => \_gnd_net_\,
            in3 => \N__22641\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_RNO_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20833\,
            in1 => \N__20818\,
            in2 => \N__21005\,
            in3 => \N__20803\,
            lcout => \b2v_inst20.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_8_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__22776\,
            in1 => \N__23544\,
            in2 => \N__24631\,
            in3 => \N__29966\,
            lcout => \b2v_inst11.un1_dutycycle_53_39_d_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNITSFK3_10_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011111111"
        )
    port map (
            in0 => \N__34252\,
            in1 => \N__25532\,
            in2 => \N__25496\,
            in3 => \N__22646\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNITSFK3Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI9LPN6_10_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001111111111"
        )
    port map (
            in0 => \N__24995\,
            in1 => \N__27650\,
            in2 => \N__19592\,
            in3 => \N__34812\,
            lcout => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10\,
            ltout => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI3ER99_10_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31226\,
            in1 => \N__19576\,
            in2 => \N__19589\,
            in3 => \N__22555\,
            lcout => \b2v_inst11.dutycycleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_10_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__19586\,
            in2 => \N__19580\,
            in3 => \N__31227\,
            lcout => \b2v_inst11.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36604\,
            ce => 'H',
            sr => \N__31043\
        );

    \b2v_inst11.dutycycle_RNIQ9K59_9_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31225\,
            in1 => \N__19675\,
            in2 => \N__19562\,
            in3 => \N__22684\,
            lcout => \b2v_inst11.dutycycleZ0Z_1\,
            ltout => \b2v_inst11.dutycycleZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNITSFK3_9_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__25531\,
            in1 => \N__25492\,
            in2 => \N__19568\,
            in3 => \N__34251\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNITSFK3Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI9LPN6_9_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011111"
        )
    port map (
            in0 => \N__34811\,
            in1 => \N__24994\,
            in2 => \N__19565\,
            in3 => \N__27646\,
            lcout => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9\,
            ltout => \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_9_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__22685\,
            in1 => \N__19676\,
            in2 => \N__19679\,
            in3 => \N__31228\,
            lcout => \b2v_inst11.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36604\,
            ce => 'H',
            sr => \N__31043\
        );

    \b2v_inst11.dutycycle_RNI_4_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24608\,
            in2 => \_gnd_net_\,
            in3 => \N__22774\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_30_a1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_7_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001110"
        )
    port map (
            in0 => \N__23542\,
            in1 => \N__22637\,
            in2 => \N__19664\,
            in3 => \N__22912\,
            lcout => \b2v_inst11.un1_dutycycle_53_44_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_13_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__25138\,
            in1 => \N__25081\,
            in2 => \N__22660\,
            in3 => \N__24916\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_13_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19625\,
            in1 => \N__19650\,
            in2 => \N__19655\,
            in3 => \N__19637\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_6_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25423\,
            in1 => \N__22773\,
            in2 => \N__25142\,
            in3 => \N__29964\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_4_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__22772\,
            in1 => \N__25134\,
            in2 => \N__24627\,
            in3 => \N__25424\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_8_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23541\,
            in2 => \N__25141\,
            in3 => \N__22771\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_8\,
            ltout => \b2v_inst11.dutycycle_RNI_3Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_11_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000100"
        )
    port map (
            in0 => \N__20921\,
            in1 => \N__25215\,
            in2 => \N__19619\,
            in3 => \N__22636\,
            lcout => \b2v_inst11.un1_dutycycle_53_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_11_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111111"
        )
    port map (
            in0 => \N__25060\,
            in1 => \N__22650\,
            in2 => \N__22795\,
            in3 => \N__25197\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010000000"
        )
    port map (
            in0 => \N__22913\,
            in1 => \N__23553\,
            in2 => \N__23438\,
            in3 => \N__24555\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_7\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_5_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22788\,
            in1 => \N__35192\,
            in2 => \N__19706\,
            in3 => \N__29941\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__23434\,
            in1 => \N__30168\,
            in2 => \N__31378\,
            in3 => \N__24557\,
            lcout => \b2v_inst11.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_0_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__24556\,
            in1 => \N__31365\,
            in2 => \_gnd_net_\,
            in3 => \N__30167\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_12_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21035\,
            in1 => \N__23554\,
            in2 => \N__25088\,
            in3 => \N__22789\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_13_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__25061\,
            in1 => \N__19703\,
            in2 => \N__23095\,
            in3 => \N__24917\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21601\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20153\,
            in3 => \N__19682\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19739\,
            in3 => \N__19892\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32048\,
            in2 => \N__19730\,
            in3 => \N__19883\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19880\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__20169\,
            in1 => \N__20170\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21602\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_15_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24713\,
            in3 => \N__19859\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19850\,
            in2 => \N__19817\,
            in3 => \N__19787\,
            lcout => \b2v_inst11.curr_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36652\,
            ce => \N__32184\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21584\,
            in3 => \N__21558\,
            lcout => \b2v_inst11.mult1_un47_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21582\,
            in2 => \N__21563\,
            in3 => \N__21538\,
            lcout => \b2v_inst11.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__21583\,
            in1 => \_gnd_net_\,
            in2 => \N__21542\,
            in3 => \N__21562\,
            lcout => \b2v_inst11.mult1_un40_sum_i_5\,
            ltout => \b2v_inst11.mult1_un40_sum_i_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20186\,
            in3 => \N__20182\,
            lcout => \b2v_inst11.mult1_un47_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21578\,
            lcout => \b2v_inst11.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI4M8F1_10_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20144\,
            in1 => \N__20123\,
            in2 => \_gnd_net_\,
            in3 => \N__20107\,
            lcout => \b2v_inst16.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21109\,
            lcout => \b2v_inst11.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIANKU4_14_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001100"
        )
    port map (
            in0 => \N__25322\,
            in1 => \N__24993\,
            in2 => \N__34286\,
            in3 => \N__23087\,
            lcout => \b2v_inst11.N_155_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20444\,
            lcout => \b2v_inst11.mult1_un117_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__32813\,
            in1 => \N__27464\,
            in2 => \N__30688\,
            in3 => \N__27533\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21836\,
            lcout => \b2v_inst11.un85_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21745\,
            lcout => \b2v_inst11.mult1_un124_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22124\,
            lcout => \b2v_inst11.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20540\,
            lcout => \b2v_inst11.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21139\,
            lcout => \b2v_inst11.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21454\,
            lcout => \b2v_inst11.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21646\,
            lcout => \b2v_inst11.mult1_un131_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21962\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20240\,
            lcout => \b2v_inst11.mult1_un103_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21529\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20318\,
            in2 => \N__20510\,
            in3 => \N__20312\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21757\,
            in2 => \N__21704\,
            in3 => \N__20309\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20471\,
            in2 => \N__21746\,
            in3 => \N__20306\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21744\,
            in2 => \N__20456\,
            in3 => \N__20303\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21641\,
            in1 => \N__20350\,
            in2 => \N__20339\,
            in3 => \N__20300\,
            lcout => \b2v_inst11.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20378\,
            in3 => \N__20297\,
            lcout => \b2v_inst11.mult1_un131_sum_s_8\,
            ltout => \b2v_inst11.mult1_un131_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20294\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21184\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20492\,
            in2 => \N__20395\,
            in3 => \N__20483\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20391\,
            in2 => \N__20480\,
            in3 => \N__20465\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20462\,
            in2 => \N__20440\,
            in3 => \N__20447\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20436\,
            in2 => \N__20414\,
            in3 => \N__20405\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21736\,
            in1 => \N__20402\,
            in2 => \N__20396\,
            in3 => \N__20369\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20366\,
            in3 => \N__20357\,
            lcout => \b2v_inst11.mult1_un124_sum_s_8\,
            ltout => \b2v_inst11.mult1_un124_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20354\,
            in3 => \N__20351\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_1_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__33305\,
            in1 => \N__31369\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.g3_0\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30038\,
            in2 => \N__22090\,
            in3 => \N__20588\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22086\,
            in2 => \N__22010\,
            in3 => \N__20576\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21989\,
            in2 => \N__22120\,
            in3 => \N__20567\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22116\,
            in2 => \N__21974\,
            in3 => \N__20558\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20535\,
            in1 => \N__21923\,
            in2 => \N__22091\,
            in3 => \N__20546\,
            lcout => \b2v_inst11.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22148\,
            in3 => \N__20543\,
            lcout => \b2v_inst11.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21727\,
            lcout => \b2v_inst11.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31379\,
            lcout => \b2v_inst11.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_1_c_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22379\,
            in2 => \N__22358\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => \b2v_inst20.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24239\,
            in2 => \_gnd_net_\,
            in3 => \N__20645\,
            lcout => \b2v_inst20.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_1\,
            carryout => \b2v_inst20.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24128\,
            in2 => \_gnd_net_\,
            in3 => \N__20642\,
            lcout => \b2v_inst20.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_2\,
            carryout => \b2v_inst20.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22283\,
            in2 => \_gnd_net_\,
            in3 => \N__20639\,
            lcout => \b2v_inst20.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_3\,
            carryout => \b2v_inst20.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22310\,
            in2 => \_gnd_net_\,
            in3 => \N__20636\,
            lcout => \b2v_inst20.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_4\,
            carryout => \b2v_inst20.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22400\,
            in2 => \_gnd_net_\,
            in3 => \N__20633\,
            lcout => \b2v_inst20.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_5\,
            carryout => \b2v_inst20.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_7_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22234\,
            in2 => \_gnd_net_\,
            in3 => \N__20630\,
            lcout => \b2v_inst20.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_6\,
            carryout => \b2v_inst20.counter_1_cry_7\,
            clk => \N__36193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_8_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20627\,
            in2 => \_gnd_net_\,
            in3 => \N__20615\,
            lcout => \b2v_inst20.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_7\,
            carryout => \b2v_inst20.counter_1_cry_8\,
            clk => \N__36193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_9_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20612\,
            in2 => \_gnd_net_\,
            in3 => \N__20600\,
            lcout => \b2v_inst20.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \b2v_inst20.counter_1_cry_9\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_10_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20788\,
            in2 => \_gnd_net_\,
            in3 => \N__20774\,
            lcout => \b2v_inst20.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_9\,
            carryout => \b2v_inst20.counter_1_cry_10\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_11_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20771\,
            in2 => \_gnd_net_\,
            in3 => \N__20759\,
            lcout => \b2v_inst20.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_10\,
            carryout => \b2v_inst20.counter_1_cry_11\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_12_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20756\,
            in2 => \_gnd_net_\,
            in3 => \N__20744\,
            lcout => \b2v_inst20.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_11\,
            carryout => \b2v_inst20.counter_1_cry_12\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_13_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20741\,
            in2 => \_gnd_net_\,
            in3 => \N__20729\,
            lcout => \b2v_inst20.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_12\,
            carryout => \b2v_inst20.counter_1_cry_13\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_14_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20725\,
            in2 => \_gnd_net_\,
            in3 => \N__20711\,
            lcout => \b2v_inst20.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_13\,
            carryout => \b2v_inst20.counter_1_cry_14\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_15_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20708\,
            in2 => \_gnd_net_\,
            in3 => \N__20696\,
            lcout => \b2v_inst20.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_14\,
            carryout => \b2v_inst20.counter_1_cry_15\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_16_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20693\,
            in2 => \_gnd_net_\,
            in3 => \N__20681\,
            lcout => \b2v_inst20.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_15\,
            carryout => \b2v_inst20.counter_1_cry_16\,
            clk => \N__36167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_17_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20677\,
            in2 => \_gnd_net_\,
            in3 => \N__20663\,
            lcout => \b2v_inst20.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \b2v_inst20.counter_1_cry_17\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_18_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20660\,
            in2 => \_gnd_net_\,
            in3 => \N__20648\,
            lcout => \b2v_inst20.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_17\,
            carryout => \b2v_inst20.counter_1_cry_18\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_19_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20912\,
            in2 => \_gnd_net_\,
            in3 => \N__20900\,
            lcout => \b2v_inst20.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_18\,
            carryout => \b2v_inst20.counter_1_cry_19\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_20_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20896\,
            in2 => \_gnd_net_\,
            in3 => \N__20882\,
            lcout => \b2v_inst20.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_19\,
            carryout => \b2v_inst20.counter_1_cry_20\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_21_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20879\,
            in2 => \_gnd_net_\,
            in3 => \N__20867\,
            lcout => \b2v_inst20.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_20\,
            carryout => \b2v_inst20.counter_1_cry_21\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_22_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20864\,
            in2 => \_gnd_net_\,
            in3 => \N__20852\,
            lcout => \b2v_inst20.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_21\,
            carryout => \b2v_inst20.counter_1_cry_22\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_23_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20849\,
            in2 => \_gnd_net_\,
            in3 => \N__20837\,
            lcout => \b2v_inst20.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_22\,
            carryout => \b2v_inst20.counter_1_cry_23\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_24_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20834\,
            in2 => \_gnd_net_\,
            in3 => \N__20822\,
            lcout => \b2v_inst20.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_23\,
            carryout => \b2v_inst20.counter_1_cry_24\,
            clk => \N__36322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_25_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20819\,
            in2 => \_gnd_net_\,
            in3 => \N__20807\,
            lcout => \b2v_inst20.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \b2v_inst20.counter_1_cry_25\,
            clk => \N__36339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_26_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20804\,
            in2 => \_gnd_net_\,
            in3 => \N__20792\,
            lcout => \b2v_inst20.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_25\,
            carryout => \b2v_inst20.counter_1_cry_26\,
            clk => \N__36339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_27_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21004\,
            in2 => \_gnd_net_\,
            in3 => \N__20990\,
            lcout => \b2v_inst20.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_26\,
            carryout => \b2v_inst20.counter_1_cry_27\,
            clk => \N__36339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_28_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20975\,
            in3 => \N__20987\,
            lcout => \b2v_inst20.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_27\,
            carryout => \b2v_inst20.counter_1_cry_28\,
            clk => \N__36339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_29_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20963\,
            in3 => \N__20984\,
            lcout => \b2v_inst20.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_28\,
            carryout => \b2v_inst20.counter_1_cry_29\,
            clk => \N__36339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_30_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20951\,
            in3 => \N__20981\,
            lcout => \b2v_inst20.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_29\,
            carryout => \b2v_inst20.counter_1_cry_30\,
            clk => \N__36339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_31_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20978\,
            lcout => \b2v_inst20.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_RNO_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20971\,
            in1 => \N__20959\,
            in2 => \N__20950\,
            in3 => \N__20935\,
            lcout => \b2v_inst20.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_8_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__22760\,
            in1 => \N__25450\,
            in2 => \_gnd_net_\,
            in3 => \N__23531\,
            lcout => \b2v_inst11.un1_dutycycle_53_9_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIO6J59_8_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__31221\,
            in1 => \N__21055\,
            in2 => \N__22814\,
            in3 => \N__23587\,
            lcout => \b2v_inst11.dutycycleZ1Z_5\,
            ltout => \b2v_inst11.dutycycleZ1Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_3_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__22761\,
            in1 => \N__24567\,
            in2 => \N__20915\,
            in3 => \N__23422\,
            lcout => \b2v_inst11.un1_dutycycle_53_3_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_8_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__22813\,
            in1 => \N__21056\,
            in2 => \N__31244\,
            in3 => \N__23588\,
            lcout => \b2v_inst11.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36437\,
            ce => 'H',
            sr => \N__31032\
        );

    \b2v_inst11.dutycycle_RNI_7_3_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__23435\,
            in1 => \N__25451\,
            in2 => \N__22790\,
            in3 => \N__23532\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_7Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_7_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__21047\,
            in1 => \N__22914\,
            in2 => \N__21041\,
            in3 => \N__29969\,
            lcout => \b2v_inst11.dutycycle_RNI_8Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100010101"
        )
    port map (
            in0 => \N__23543\,
            in1 => \N__24568\,
            in2 => \N__22791\,
            in3 => \N__25452\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_26_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_7_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001100"
        )
    port map (
            in0 => \N__25453\,
            in1 => \N__22915\,
            in2 => \N__21038\,
            in3 => \N__29970\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIGFG69_13_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__21025\,
            in1 => \N__33850\,
            in2 => \N__24731\,
            in3 => \N__23017\,
            lcout => \b2v_inst11.dutycycleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_13_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__23018\,
            in1 => \N__21026\,
            in2 => \N__33887\,
            in3 => \N__24727\,
            lcout => \b2v_inst11.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36198\,
            ce => 'H',
            sr => \N__31039\
        );

    \b2v_inst11.dutycycle_4_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__23198\,
            in1 => \N__21016\,
            in2 => \N__22943\,
            in3 => \N__33854\,
            lcout => \b2v_inst11.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36198\,
            ce => 'H',
            sr => \N__31039\
        );

    \b2v_inst11.dutycycle_RNIGQE59_4_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33849\,
            in1 => \N__22939\,
            in2 => \N__21017\,
            in3 => \N__23197\,
            lcout => \b2v_inst11.dutycycleZ0Z_7\,
            ltout => \b2v_inst11.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_4_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21086\,
            in3 => \N__22781\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_7_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111000110"
        )
    port map (
            in0 => \N__21083\,
            in1 => \N__21071\,
            in2 => \N__21077\,
            in3 => \N__22918\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_11_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__25219\,
            in1 => \_gnd_net_\,
            in2 => \N__21074\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_11_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25218\,
            in2 => \_gnd_net_\,
            in3 => \N__23546\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_2_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__23398\,
            in1 => \_gnd_net_\,
            in2 => \N__29971\,
            in3 => \N__33191\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100101101"
        )
    port map (
            in0 => \N__31374\,
            in1 => \N__33707\,
            in2 => \N__21065\,
            in3 => \N__24588\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_2_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21062\,
            in3 => \N__33192\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_7_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001010110100"
        )
    port map (
            in0 => \N__22917\,
            in1 => \N__24595\,
            in2 => \N__23570\,
            in3 => \N__23401\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__23399\,
            in1 => \N__31375\,
            in2 => \N__24621\,
            in3 => \N__29957\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_5_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__21209\,
            in1 => \N__21161\,
            in2 => \N__21059\,
            in3 => \N__35184\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_7_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__23400\,
            in1 => \_gnd_net_\,
            in2 => \N__24622\,
            in3 => \N__22916\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_3_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__31373\,
            in1 => \N__29953\,
            in2 => \_gnd_net_\,
            in3 => \N__23397\,
            lcout => \b2v_inst11.d_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30176\,
            in2 => \N__23423\,
            in3 => \N__31376\,
            lcout => \b2v_inst11.g0_i_a7_1_2\,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21203\,
            in2 => \N__30184\,
            in3 => \N__21197\,
            lcout => \b2v_inst11.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33166\,
            in2 => \N__24491\,
            in3 => \N__21194\,
            lcout => \b2v_inst11.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_1\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21191\,
            in2 => \N__33186\,
            in3 => \N__21164\,
            lcout => \b2v_inst11.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_2\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21160\,
            in2 => \N__21149\,
            in3 => \N__21119\,
            lcout => \b2v_inst11.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_3\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21116\,
            in2 => \N__35198\,
            in3 => \N__21089\,
            lcout => \b2v_inst11.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_4\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35188\,
            in2 => \N__21506\,
            in3 => \N__21473\,
            lcout => \b2v_inst11.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_5\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22661\,
            in2 => \N__21470\,
            in3 => \N__21434\,
            lcout => \b2v_inst11.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_6\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25220\,
            in2 => \N__21431\,
            in3 => \N__21398\,
            lcout => \b2v_inst11.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25087\,
            in2 => \N__21395\,
            in3 => \N__21362\,
            lcout => \b2v_inst11.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_8\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21359\,
            in2 => \N__24950\,
            in3 => \N__21329\,
            lcout => \b2v_inst11.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_9\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21326\,
            in2 => \N__23076\,
            in3 => \N__21287\,
            lcout => \b2v_inst11.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_10\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24699\,
            in2 => \N__21284\,
            in3 => \N__21254\,
            lcout => \b2v_inst11.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_11\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24939\,
            in2 => \N__21251\,
            in3 => \N__21212\,
            lcout => \b2v_inst11.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_12\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23061\,
            in2 => \N__21614\,
            in3 => \N__21587\,
            lcout => \b2v_inst11.mult1_un47_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_13\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23282\,
            in2 => \N__24711\,
            in3 => \N__21566\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_14\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21512\,
            in2 => \N__24703\,
            in3 => \N__21548\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \b2v_inst11.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.CO2_THRU_LUT4_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21545\,
            lcout => \b2v_inst11.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21695\,
            lcout => \b2v_inst11.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o2_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34621\,
            in2 => \_gnd_net_\,
            in3 => \N__34455\,
            lcout => \b2v_inst11.N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21530\,
            lcout => \b2v_inst11.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_14_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23309\,
            in3 => \N__23057\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIL6AH3_6_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21797\,
            in1 => \N__26864\,
            in2 => \_gnd_net_\,
            in3 => \N__22459\,
            lcout => \b2v_inst5.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_6_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36403\,
            ce => \N__26865\,
            sr => \N__27341\
        );

    \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__21791\,
            in1 => \N__21773\,
            in2 => \_gnd_net_\,
            in3 => \N__34932\,
            lcout => \b2v_inst6.N_192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__34620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32873\,
            lcout => \b2v_inst11.N_161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21740\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21694\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21680\,
            in2 => \N__21904\,
            in3 => \N__21671\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_2_c\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21900\,
            in2 => \N__21668\,
            in3 => \N__21659\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_3_c\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21656\,
            in2 => \N__21647\,
            in3 => \N__21650\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_4_c\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21645\,
            in2 => \N__21623\,
            in3 => \N__21914\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_5_c\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21827\,
            in1 => \N__21911\,
            in2 => \N__21905\,
            in3 => \N__21887\,
            lcout => \b2v_inst11.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_6_c\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21884\,
            in3 => \N__21875\,
            lcout => \b2v_inst11.mult1_un138_sum_s_8\,
            ltout => \b2v_inst11.mult1_un138_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21872\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23342\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21869\,
            in2 => \N__22045\,
            in3 => \N__21860\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22041\,
            in2 => \N__21857\,
            in3 => \N__21848\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21845\,
            in2 => \N__21835\,
            in3 => \N__21839\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21831\,
            in2 => \N__21809\,
            in3 => \N__21800\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21950\,
            in1 => \N__22052\,
            in2 => \N__22046\,
            in3 => \N__22028\,
            lcout => \b2v_inst11.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22025\,
            in3 => \N__22016\,
            lcout => \b2v_inst11.mult1_un145_sum_s_8\,
            ltout => \b2v_inst11.mult1_un145_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22013\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33197\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23333\,
            in2 => \N__22165\,
            in3 => \N__22001\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22161\,
            in2 => \N__21998\,
            in3 => \N__21983\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21980\,
            in2 => \N__21958\,
            in3 => \N__21965\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21954\,
            in2 => \N__21932\,
            in3 => \N__21917\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22112\,
            in1 => \N__22172\,
            in2 => \N__22166\,
            in3 => \N__22139\,
            lcout => \b2v_inst11.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22136\,
            in3 => \N__22127\,
            lcout => \b2v_inst11.mult1_un152_sum_s_8\,
            ltout => \b2v_inst11.mult1_un152_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22094\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIB8QH1_0_1_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001001100"
        )
    port map (
            in0 => \N__23897\,
            in1 => \N__24054\,
            in2 => \N__29150\,
            in3 => \N__22061\,
            lcout => \b2v_inst36.un12_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIB8QH1_1_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22060\,
            in1 => \N__29134\,
            in2 => \_gnd_net_\,
            in3 => \N__23895\,
            lcout => \b2v_inst36.un2_count_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26171\,
            in1 => \N__24055\,
            in2 => \N__24038\,
            in3 => \N__28939\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIDPQG1_11_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22067\,
            in2 => \N__22073\,
            in3 => \N__29135\,
            lcout => \b2v_inst36.countZ0Z_11\,
            ltout => \b2v_inst36.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_11_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__24037\,
            in1 => \N__26173\,
            in2 => \N__22070\,
            in3 => \N__28941\,
            lcout => \b2v_inst36.count_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36001\,
            ce => \N__29141\,
            sr => \N__28938\
        );

    \b2v_inst36.count_1_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23896\,
            lcout => \b2v_inst36.count_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36001\,
            ce => \N__29141\,
            sr => \N__28938\
        );

    \b2v_inst36.count_0_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__26172\,
            in1 => \N__22185\,
            in2 => \_gnd_net_\,
            in3 => \N__28940\,
            lcout => \b2v_inst36.count_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36001\,
            ce => \N__29141\,
            sr => \N__28938\
        );

    \b2v_inst36.count_RNI1FG91_0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__22186\,
            in1 => \N__28937\,
            in2 => \_gnd_net_\,
            in3 => \N__26170\,
            lcout => \b2v_inst36.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI6K3V_0_0_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24016\,
            in1 => \N__23950\,
            in2 => \N__22190\,
            in3 => \N__23986\,
            lcout => \b2v_inst36.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIL5VG1_15_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22208\,
            in1 => \N__29147\,
            in2 => \_gnd_net_\,
            in3 => \N__24263\,
            lcout => \b2v_inst36.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_15_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36192\,
            ce => \N__29146\,
            sr => \N__28981\
        );

    \b2v_inst36.count_RNIHVSG1_13_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22202\,
            in1 => \N__29108\,
            in2 => \_gnd_net_\,
            in3 => \N__24001\,
            lcout => \b2v_inst36.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_13_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36192\,
            ce => \N__29146\,
            sr => \N__28981\
        );

    \b2v_inst36.count_RNIJ2UG1_14_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22196\,
            in1 => \N__29109\,
            in2 => \_gnd_net_\,
            in3 => \N__23971\,
            lcout => \b2v_inst36.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_14_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36192\,
            ce => \N__29146\,
            sr => \N__28981\
        );

    \b2v_inst36.count_RNI6K3V_0_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__23936\,
            in1 => \N__29110\,
            in2 => \_gnd_net_\,
            in3 => \N__23924\,
            lcout => \b2v_inst36.count_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_7_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22433\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => \N__26872\,
            sr => \N__27343\
        );

    \b2v_inst5.count_RNID0AN3_11_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22521\,
            in1 => \N__22252\,
            in2 => \_gnd_net_\,
            in3 => \N__26856\,
            lcout => \b2v_inst5.un2_count_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_11_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22522\,
            lcout => \b2v_inst5.count_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => \N__26872\,
            sr => \N__27343\
        );

    \b2v_inst5.count_RNIN9BH3_7_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22259\,
            in1 => \N__26855\,
            in2 => \_gnd_net_\,
            in3 => \N__22432\,
            lcout => \b2v_inst5.countZ0Z_7\,
            ltout => \b2v_inst5.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNID0AN3_0_11_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__22253\,
            in1 => \N__26873\,
            in2 => \N__22244\,
            in3 => \N__22523\,
            lcout => \b2v_inst5.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIF3BN3_12_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__22241\,
            in1 => \N__22504\,
            in2 => \N__27342\,
            in3 => \N__26857\,
            lcout => \b2v_inst5.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_12_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27335\,
            lcout => \b2v_inst5.count_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => \N__26872\,
            sr => \N__27343\
        );

    \b2v_inst5.count_14_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24332\,
            in2 => \_gnd_net_\,
            in3 => \N__27344\,
            lcout => \b2v_inst5.count_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => \N__26872\,
            sr => \N__27343\
        );

    \b2v_inst20.un4_counter_1_c_RNO_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__22235\,
            in1 => \N__22305\,
            in2 => \N__22399\,
            in3 => \N__22371\,
            lcout => \b2v_inst20.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_6_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24190\,
            in1 => \N__22409\,
            in2 => \_gnd_net_\,
            in3 => \N__22395\,
            lcout => \b2v_inst20.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_0_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__22351\,
            in1 => \N__24192\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst20.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__24191\,
            in1 => \_gnd_net_\,
            in2 => \N__22378\,
            in3 => \N__22350\,
            lcout => \b2v_inst20.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_RNO_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22349\,
            in1 => \N__24228\,
            in2 => \N__22282\,
            in3 => \N__24120\,
            lcout => \b2v_inst20.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_5_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__22306\,
            in1 => \_gnd_net_\,
            in2 => \N__24194\,
            in3 => \N__22322\,
            lcout => \b2v_inst20.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_4_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__22278\,
            in1 => \N__22292\,
            in2 => \_gnd_net_\,
            in3 => \N__24193\,
            lcout => \b2v_inst20.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__27463\,
            in1 => \N__27044\,
            in2 => \N__27071\,
            in3 => \N__27532\,
            lcout => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_0_c_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24341\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_0_c_RNIKSVJ1_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27307\,
            in1 => \N__26519\,
            in2 => \_gnd_net_\,
            in3 => \N__22262\,
            lcout => \b2v_inst5.count_rst_13\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_0\,
            carryout => \b2v_inst5.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_1_c_RNILU0K1_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27305\,
            in1 => \N__26498\,
            in2 => \_gnd_net_\,
            in3 => \N__22472\,
            lcout => \b2v_inst5.count_rst_12\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_1\,
            carryout => \b2v_inst5.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_2_c_RNIM02K1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__27309\,
            in1 => \_gnd_net_\,
            in2 => \N__26555\,
            in3 => \N__22469\,
            lcout => \b2v_inst5.count_rst_11\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_2\,
            carryout => \b2v_inst5.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24437\,
            in2 => \_gnd_net_\,
            in3 => \N__22466\,
            lcout => \b2v_inst5.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_3\,
            carryout => \b2v_inst5.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_4_c_RNIO44K1_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27308\,
            in1 => \N__26429\,
            in2 => \_gnd_net_\,
            in3 => \N__22463\,
            lcout => \b2v_inst5.count_rst_9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_4\,
            carryout => \b2v_inst5.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_5_c_RNIP65K1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27304\,
            in1 => \N__26398\,
            in2 => \_gnd_net_\,
            in3 => \N__22445\,
            lcout => \b2v_inst5.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_5\,
            carryout => \b2v_inst5.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_6_c_RNIQ86K1_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27306\,
            in1 => \N__22442\,
            in2 => \_gnd_net_\,
            in3 => \N__22421\,
            lcout => \b2v_inst5.count_rst_7\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_6\,
            carryout => \b2v_inst5.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24472\,
            in2 => \_gnd_net_\,
            in3 => \N__22418\,
            lcout => \b2v_inst5.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27023\,
            in2 => \_gnd_net_\,
            in3 => \N__22415\,
            lcout => \b2v_inst5.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_8\,
            carryout => \b2v_inst5.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26651\,
            in2 => \_gnd_net_\,
            in3 => \N__22412\,
            lcout => \b2v_inst5.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_9\,
            carryout => \b2v_inst5.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27313\,
            in1 => \N__22535\,
            in2 => \_gnd_net_\,
            in3 => \N__22508\,
            lcout => \b2v_inst5.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_10\,
            carryout => \b2v_inst5.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24289\,
            in2 => \_gnd_net_\,
            in3 => \N__22493\,
            lcout => \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_11\,
            carryout => \b2v_inst5.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26535\,
            in2 => \_gnd_net_\,
            in3 => \N__22490\,
            lcout => \b2v_inst5.un2_count_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_12\,
            carryout => \b2v_inst5.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24308\,
            in2 => \_gnd_net_\,
            in3 => \N__22487\,
            lcout => \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_13\,
            carryout => \b2v_inst5.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27314\,
            in1 => \N__26615\,
            in2 => \_gnd_net_\,
            in3 => \N__22484\,
            lcout => \b2v_inst5.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_c_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30175\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31350\,
            in2 => \N__27141\,
            in3 => \N__22481\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27130\,
            in2 => \N__33196\,
            in3 => \N__22478\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27135\,
            in2 => \N__23425\,
            in3 => \N__22475\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_2\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27131\,
            in2 => \N__24596\,
            in3 => \N__22928\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_3\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35183\,
            in2 => \N__27142\,
            in3 => \N__22925\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_4\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29906\,
            in2 => \N__27143\,
            in3 => \N__22922\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27139\,
            in2 => \N__22919\,
            in3 => \N__22817\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9J1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__33842\,
            in1 => \N__27118\,
            in2 => \N__23568\,
            in3 => \N__22799\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9JZ0Z1\,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJ1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__33881\,
            in1 => \N__27121\,
            in2 => \N__22796\,
            in3 => \N__22670\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJZ0Z1\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJ1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__33843\,
            in1 => \N__27119\,
            in2 => \N__22667\,
            in3 => \N__22541\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJZ0Z1\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_9\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUF1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__33882\,
            in1 => \N__27122\,
            in2 => \N__25196\,
            in3 => \N__22538\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUFZ0Z1\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_10\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_11_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_11_c_RNI9KVF1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__33844\,
            in1 => \N__25037\,
            in2 => \N__27140\,
            in3 => \N__23021\,
            lcout => \b2v_inst11.dutycycle_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_11_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_12_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27126\,
            in2 => \N__24935\,
            in3 => \N__23009\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_12_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_13_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27120\,
            in2 => \N__23086\,
            in3 => \N__23006\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_13_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24704\,
            in1 => \N__33411\,
            in2 => \_gnd_net_\,
            in3 => \N__23003\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIANKU4_3_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__34289\,
            in1 => \N__25301\,
            in2 => \N__22994\,
            in3 => \N__23449\,
            lcout => \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0\,
            ltout => \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI61IA9_3_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__34799\,
            in1 => \N__22976\,
            in2 => \N__23000\,
            in3 => \N__22956\,
            lcout => \b2v_inst11.dutycycleZ0Z_3\,
            ltout => \b2v_inst11.dutycycleZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_3_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22997\,
            in3 => \N__25246\,
            lcout => \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI52KD2_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__22985\,
            in1 => \N__33848\,
            in2 => \N__22961\,
            in3 => \N__31193\,
            lcout => \b2v_inst11.dutycycle_e_1_3\,
            ltout => \b2v_inst11.dutycycle_e_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_3_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__22957\,
            in1 => \N__22970\,
            in2 => \N__22964\,
            in3 => \N__34800\,
            lcout => \b2v_inst11.dutycycle_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36099\,
            ce => 'H',
            sr => \N__31038\
        );

    \b2v_inst11.dutycycle_RNITSFK3_4_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__25302\,
            in1 => \N__34290\,
            in2 => \N__25250\,
            in3 => \N__24623\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_40_and_i_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIT35D7_4_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__31192\,
            in1 => \N__34798\,
            in2 => \N__23201\,
            in3 => \N__23450\,
            lcout => \b2v_inst11.dutycycle_RNIT35D7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIKLI69_15_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__23140\,
            in1 => \N__33846\,
            in2 => \N__23165\,
            in3 => \N__23155\,
            lcout => \b2v_inst11.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIT35D7_14_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010100010"
        )
    port map (
            in0 => \N__31194\,
            in1 => \N__34804\,
            in2 => \N__23186\,
            in3 => \N__27643\,
            lcout => \b2v_inst11.dutycycle_en_11\,
            ltout => \b2v_inst11.dutycycle_en_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_14_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__23129\,
            in1 => \N__33847\,
            in2 => \N__23171\,
            in3 => \N__23111\,
            lcout => \b2v_inst11.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36394\,
            ce => 'H',
            sr => \N__31021\
        );

    \b2v_inst11.dutycycle_RNIANKU4_15_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001100"
        )
    port map (
            in0 => \N__25320\,
            in1 => \N__24987\,
            in2 => \N__34285\,
            in3 => \N__24688\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_158_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIT35D7_15_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001100"
        )
    port map (
            in0 => \N__27644\,
            in1 => \N__31195\,
            in2 => \N__23168\,
            in3 => \N__34805\,
            lcout => \b2v_inst11.dutycycle_RNIT35D7Z0Z_15\,
            ltout => \b2v_inst11.dutycycle_RNIT35D7Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_15_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__23156\,
            in1 => \N__33917\,
            in2 => \N__23144\,
            in3 => \N__23141\,
            lcout => \b2v_inst11.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36394\,
            ce => 'H',
            sr => \N__31021\
        );

    \b2v_inst11.dutycycle_RNIIIH69_14_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__23128\,
            in1 => \N__33845\,
            in2 => \N__23120\,
            in3 => \N__23110\,
            lcout => \b2v_inst11.dutycycleZ0Z_12\,
            ltout => \b2v_inst11.dutycycleZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_14_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24689\,
            in2 => \N__23312\,
            in3 => \N__23305\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIM50S4_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__23273\,
            in1 => \N__34807\,
            in2 => \N__23261\,
            in3 => \N__33929\,
            lcout => \b2v_inst11.dutycycle_set_1\,
            ltout => \b2v_inst11.dutycycle_set_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_5_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__23219\,
            in1 => \N__31191\,
            in2 => \N__23264\,
            in3 => \N__34643\,
            lcout => \b2v_inst11.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36315\,
            ce => 'H',
            sr => \N__31020\
        );

    \b2v_inst11.func_state_RNISPKF1_0_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__29638\,
            in1 => \N__33415\,
            in2 => \N__34287\,
            in3 => \N__30276\,
            lcout => \b2v_inst11.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIBGDMD_6_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__23237\,
            in1 => \N__23227\,
            in2 => \N__23606\,
            in3 => \N__31190\,
            lcout => \b2v_inst11.dutycycleZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNISPKF1_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__29639\,
            in1 => \N__33416\,
            in2 => \N__34288\,
            in3 => \N__30277\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_300_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIN71S4_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110011"
        )
    port map (
            in0 => \N__33928\,
            in1 => \N__34806\,
            in2 => \N__23252\,
            in3 => \N__23249\,
            lcout => \b2v_inst11.dutycycle_set_0_0\,
            ltout => \b2v_inst11.dutycycle_set_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_6_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__23228\,
            in1 => \N__31249\,
            in2 => \N__23231\,
            in3 => \N__23605\,
            lcout => \b2v_inst11.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36315\,
            ce => 'H',
            sr => \N__31020\
        );

    \b2v_inst11.dutycycle_RNIFNB2O_5_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__23218\,
            in1 => \N__31189\,
            in2 => \N__23210\,
            in3 => \N__34642\,
            lcout => \b2v_inst11.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5DSV7_6_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111111111"
        )
    port map (
            in0 => \N__23321\,
            in1 => \N__24866\,
            in2 => \N__25259\,
            in3 => \N__34796\,
            lcout => \b2v_inst11.dutycycle_eena_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_6_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33049\,
            lcout => \b2v_inst11.N_200_i\,
            ltout => \b2v_inst11.N_200_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__33886\,
            in1 => \_gnd_net_\,
            in2 => \N__23594\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI9LPN6_8_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__34797\,
            in1 => \N__23456\,
            in2 => \N__23591\,
            in3 => \N__25240\,
            lcout => \b2v_inst11.dutycycle_eena_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNITSFK3_8_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__25239\,
            in1 => \N__25316\,
            in2 => \N__34311\,
            in3 => \N__23569\,
            lcout => \b2v_inst11.un1_clk_100khz_32_and_i_0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33885\,
            in2 => \N__33279\,
            in3 => \N__25238\,
            lcout => \b2v_inst11.un1_clk_100khz_40_and_i_0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23424\,
            in2 => \_gnd_net_\,
            in3 => \N__30154\,
            lcout => \b2v_inst11.mult1_un145_sum\,
            ltout => \b2v_inst11.mult1_un145_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23336\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIGUKJ1_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__34457\,
            in1 => \N__30275\,
            in2 => \N__34312\,
            in3 => \N__33417\,
            lcout => \b2v_inst11.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_7_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__28422\,
            in1 => \N__23615\,
            in2 => \_gnd_net_\,
            in3 => \N__23663\,
            lcout => \b2v_inst11.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_8_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25717\,
            lcout => \b2v_inst11.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36479\,
            ce => \N__28570\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI342J_8_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__30637\,
            in1 => \N__28489\,
            in2 => \N__25721\,
            in3 => \N__23630\,
            lcout => \b2v_inst11.count_clkZ0Z_8\,
            ltout => \b2v_inst11.count_clkZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_2_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__25831\,
            in1 => \N__25868\,
            in2 => \N__23624\,
            in3 => \N__25655\,
            lcout => OPEN,
            ltout => \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_6_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__25765\,
            in1 => \N__28424\,
            in2 => \N__23621\,
            in3 => \N__23662\,
            lcout => \b2v_inst11.count_clk_RNIZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_3_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__25863\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25732\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_2_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__25764\,
            in1 => \N__25653\,
            in2 => \N__23618\,
            in3 => \N__25830\,
            lcout => \b2v_inst11.N_379\,
            ltout => \b2v_inst11.N_379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28214\,
            in1 => \N__28423\,
            in2 => \N__23609\,
            in3 => \N__23645\,
            lcout => \b2v_inst11.count_clk_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_9_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36481\,
            ce => \N__28541\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI573J_9_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__30635\,
            in1 => \N__28542\,
            in2 => \N__23675\,
            in3 => \N__25693\,
            lcout => \b2v_inst11.count_clkZ0Z_9\,
            ltout => \b2v_inst11.count_clkZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_1_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__23723\,
            in1 => \N__25801\,
            in2 => \N__23666\,
            in3 => \N__28215\,
            lcout => \b2v_inst11.N_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_5_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25783\,
            lcout => \b2v_inst11.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36481\,
            ce => \N__28541\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNITQUI_5_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__28539\,
            in1 => \N__23654\,
            in2 => \N__25787\,
            in3 => \N__30636\,
            lcout => \b2v_inst11.count_clkZ0Z_5\,
            ltout => \b2v_inst11.count_clkZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_5_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__25705\,
            in1 => \_gnd_net_\,
            in2 => \N__23648\,
            in3 => \N__23722\,
            lcout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIQA5D_1_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__28540\,
            in1 => \N__23636\,
            in2 => \N__30706\,
            in3 => \N__28190\,
            lcout => \b2v_inst11.count_clkZ0Z_1\,
            ltout => \b2v_inst11.count_clkZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_1_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28110\,
            in2 => \N__23639\,
            in3 => \N__28173\,
            lcout => \b2v_inst11.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36481\,
            ce => \N__28541\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_11_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25882\,
            lcout => \b2v_inst11.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36485\,
            ce => \N__28568\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_14_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25918\,
            lcout => \b2v_inst11.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36485\,
            ce => \N__28568\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVFGI_15_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28571\,
            in1 => \N__30634\,
            in2 => \N__23708\,
            in3 => \N__25897\,
            lcout => \b2v_inst11.count_clkZ0Z_15\,
            ltout => \b2v_inst11.count_clkZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_15_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25930\,
            in1 => \N__28325\,
            in2 => \N__23726\,
            in3 => \N__28177\,
            lcout => \b2v_inst11.N_175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNITCFI_14_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__25919\,
            in1 => \N__23714\,
            in2 => \N__30727\,
            in3 => \N__28569\,
            lcout => \b2v_inst11.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_15_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25898\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36485\,
            ce => \N__28568\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIFESH1_3_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23686\,
            in1 => \N__29117\,
            in2 => \_gnd_net_\,
            in3 => \N__23696\,
            lcout => \b2v_inst36.un2_count_1_axb_3\,
            ltout => \b2v_inst36.un2_count_1_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26142\,
            in1 => \N__23827\,
            in2 => \N__23699\,
            in3 => \N__28916\,
            lcout => \b2v_inst36.count_rst_11\,
            ltout => \b2v_inst36.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIFESH1_0_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__23687\,
            in1 => \N__29118\,
            in2 => \N__23690\,
            in3 => \N__23877\,
            lcout => \b2v_inst36.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_3_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26143\,
            in1 => \N__23828\,
            in2 => \N__23846\,
            in3 => \N__28960\,
            lcout => \b2v_inst36.count_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__29145\,
            sr => \N__28959\
        );

    \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__23860\,
            in1 => \N__28914\,
            in2 => \N__26174\,
            in3 => \N__23878\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIDBRH1_2_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29116\,
            in1 => \_gnd_net_\,
            in2 => \N__23678\,
            in3 => \N__23762\,
            lcout => \b2v_inst36.countZ0Z_2\,
            ltout => \b2v_inst36.countZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_2_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__23861\,
            in1 => \N__28915\,
            in2 => \N__23765\,
            in3 => \N__26145\,
            lcout => \b2v_inst36.count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__29145\,
            sr => \N__28959\
        );

    \b2v_inst36.count_5_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26144\,
            in1 => \N__23786\,
            in2 => \N__23809\,
            in3 => \N__28961\,
            lcout => \b2v_inst36.count_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__29145\,
            sr => \N__28959\
        );

    \b2v_inst36.count_7_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__24082\,
            in1 => \N__28920\,
            in2 => \N__24104\,
            in3 => \N__26153\,
            lcout => \b2v_inst36.count_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36263\,
            ce => \N__29096\,
            sr => \N__28980\
        );

    \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__28918\,
            in1 => \N__24103\,
            in2 => \N__24086\,
            in3 => \N__26147\,
            lcout => \b2v_inst36.count_rst_7\,
            ltout => \b2v_inst36.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNINQ0I1_7_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29095\,
            in1 => \_gnd_net_\,
            in2 => \N__23756\,
            in3 => \N__23743\,
            lcout => \b2v_inst36.un2_count_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__23782\,
            in1 => \N__28917\,
            in2 => \N__23810\,
            in3 => \N__26146\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIJKUH1_5_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29094\,
            in1 => \_gnd_net_\,
            in2 => \N__23753\,
            in3 => \N__23750\,
            lcout => \b2v_inst36.countZ0Z_5\,
            ltout => \b2v_inst36.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNINQ0I1_0_7_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__23744\,
            in1 => \N__23735\,
            in2 => \N__23729\,
            in3 => \N__29097\,
            lcout => \b2v_inst36.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26148\,
            in1 => \N__25999\,
            in2 => \N__25970\,
            in3 => \N__28919\,
            lcout => \b2v_inst36.count_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_0_c_RNO_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23935\,
            in1 => \N__29093\,
            in2 => \_gnd_net_\,
            in3 => \N__23923\,
            lcout => \b2v_inst36.un2_count_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_0_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23912\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_0_c_RNI4JMI_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28945\,
            in1 => \N__23906\,
            in2 => \_gnd_net_\,
            in3 => \N__23882\,
            lcout => \b2v_inst36.count_rst_13\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_0\,
            carryout => \b2v_inst36.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23879\,
            in2 => \_gnd_net_\,
            in3 => \N__23849\,
            lcout => \b2v_inst36.un2_count_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_1\,
            carryout => \b2v_inst36.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23845\,
            in2 => \_gnd_net_\,
            in3 => \N__23816\,
            lcout => \b2v_inst36.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_2\,
            carryout => \b2v_inst36.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28973\,
            in1 => \N__26045\,
            in2 => \_gnd_net_\,
            in3 => \N__23813\,
            lcout => \b2v_inst36.count_rst_10\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_3\,
            carryout => \b2v_inst36.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23802\,
            in2 => \_gnd_net_\,
            in3 => \N__23771\,
            lcout => \b2v_inst36.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_4\,
            carryout => \b2v_inst36.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_5_c_RNILNVH1_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28974\,
            in1 => \N__26066\,
            in2 => \_gnd_net_\,
            in3 => \N__23768\,
            lcout => \b2v_inst36.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_5\,
            carryout => \b2v_inst36.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24099\,
            in2 => \_gnd_net_\,
            in3 => \N__24068\,
            lcout => \b2v_inst36.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_6\,
            carryout => \b2v_inst36.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25969\,
            in3 => \N__24065\,
            lcout => \b2v_inst36.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28964\,
            in1 => \N__29188\,
            in2 => \_gnd_net_\,
            in3 => \N__24062\,
            lcout => \b2v_inst36.count_rst_5\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_8\,
            carryout => \b2v_inst36.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26204\,
            in2 => \_gnd_net_\,
            in3 => \N__24059\,
            lcout => \b2v_inst36.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_9\,
            carryout => \b2v_inst36.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24056\,
            in2 => \_gnd_net_\,
            in3 => \N__24023\,
            lcout => \b2v_inst36.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_10\,
            carryout => \b2v_inst36.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_11_c_RNIFSRG1_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28975\,
            in1 => \N__26336\,
            in2 => \_gnd_net_\,
            in3 => \N__24020\,
            lcout => \b2v_inst36.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_11\,
            carryout => \b2v_inst36.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28963\,
            in1 => \N__24017\,
            in2 => \_gnd_net_\,
            in3 => \N__23990\,
            lcout => \b2v_inst36.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_12\,
            carryout => \b2v_inst36.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28976\,
            in1 => \N__23987\,
            in2 => \_gnd_net_\,
            in3 => \N__23957\,
            lcout => \b2v_inst36.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_13\,
            carryout => \b2v_inst36.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28965\,
            in1 => \N__23954\,
            in2 => \_gnd_net_\,
            in3 => \N__23939\,
            lcout => \b2v_inst36.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24173\,
            in2 => \_gnd_net_\,
            in3 => \N__30509\,
            lcout => \SYNTHESIZED_WIRE_1keep_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_2_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24171\,
            in1 => \N__24251\,
            in2 => \_gnd_net_\,
            in3 => \N__24238\,
            lcout => \b2v_inst20.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_fast_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27045\,
            in2 => \_gnd_net_\,
            in3 => \N__24174\,
            lcout => \SYNTHESIZED_WIRE_1keep_3_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_rep1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__29608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24175\,
            lcout => \SYNTHESIZED_WIRE_1keep_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.G_146_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29607\,
            in2 => \_gnd_net_\,
            in3 => \N__24170\,
            lcout => \G_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI3E27_0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__29294\,
            in1 => \N__29242\,
            in2 => \_gnd_net_\,
            in3 => \N__29342\,
            lcout => OPEN,
            ltout => \b2v_inst36.curr_state_RNI3E27Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_RNIPUMD_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__26015\,
            in1 => \_gnd_net_\,
            in2 => \N__24215\,
            in3 => \N__30510\,
            lcout => dsw_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24172\,
            in1 => \N__24140\,
            in2 => \_gnd_net_\,
            in3 => \N__24124\,
            lcout => \b2v_inst20.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24301\,
            in1 => \N__26940\,
            in2 => \_gnd_net_\,
            in3 => \N__27215\,
            lcout => \b2v_inst5.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36586\,
            ce => \N__26800\,
            sr => \N__27323\
        );

    \b2v_inst5.count_RNIH6CN3_13_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24368\,
            in1 => \N__26798\,
            in2 => \_gnd_net_\,
            in3 => \N__24377\,
            lcout => \b2v_inst5.countZ0Z_13\,
            ltout => \b2v_inst5.countZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_13_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__27324\,
            in1 => \N__26941\,
            in2 => \N__24371\,
            in3 => \N__24389\,
            lcout => \b2v_inst5.count_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36586\,
            ce => \N__26800\,
            sr => \N__27323\
        );

    \b2v_inst5.count_RNIMP4T1_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24359\,
            in1 => \N__24352\,
            in2 => \_gnd_net_\,
            in3 => \N__26796\,
            lcout => \b2v_inst5.count_i_0\,
            ltout => \b2v_inst5.count_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIL9B73_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26939\,
            in2 => \N__24362\,
            in3 => \N__27214\,
            lcout => \b2v_inst5.count_rst_14\,
            ltout => \b2v_inst5.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24353\,
            in2 => \N__24344\,
            in3 => \N__26797\,
            lcout => \b2v_inst5.un2_count_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIJ9DN3_14_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__26799\,
            in1 => \N__24328\,
            in2 => \N__27289\,
            in3 => \N__24317\,
            lcout => \b2v_inst5.countZ0Z_14\,
            ltout => \b2v_inst5.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIMP4T1_0_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__26614\,
            in1 => \N__24302\,
            in2 => \N__24293\,
            in3 => \N__24290\,
            lcout => \b2v_inst5.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIU15T1_0_8_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__24272\,
            in1 => \N__24432\,
            in2 => \N__26848\,
            in3 => \N__24449\,
            lcout => \b2v_inst5.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__27217\,
            in1 => \N__24460\,
            in2 => \N__24476\,
            in3 => \N__26963\,
            lcout => \b2v_inst5.count_rst_6\,
            ltout => \b2v_inst5.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIU15T1_8_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24448\,
            in2 => \N__24479\,
            in3 => \N__26802\,
            lcout => \b2v_inst5.un2_count_1_axb_8\,
            ltout => \b2v_inst5.un2_count_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_8_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__27219\,
            in1 => \N__24461\,
            in2 => \N__24452\,
            in3 => \N__26964\,
            lcout => \b2v_inst5.count_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36447\,
            ce => \N__26821\,
            sr => \N__27303\
        );

    \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26962\,
            in1 => \N__24433\,
            in2 => \N__24416\,
            in3 => \N__27216\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIH08H3_4_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26801\,
            in1 => \_gnd_net_\,
            in2 => \N__24440\,
            in3 => \N__24395\,
            lcout => \b2v_inst5.countZ0Z_4\,
            ltout => \b2v_inst5.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_4_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__24415\,
            in1 => \N__26979\,
            in2 => \N__24398\,
            in3 => \N__27220\,
            lcout => \b2v_inst5.count_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36447\,
            ce => \N__26821\,
            sr => \N__27303\
        );

    \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__27218\,
            in1 => \N__24388\,
            in2 => \N__26981\,
            in3 => \N__26536\,
            lcout => \b2v_inst5.count_rst_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_12_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__24812\,
            in1 => \N__24788\,
            in2 => \N__31248\,
            in3 => \N__24799\,
            lcout => \b2v_inst11.dutycycleZ1Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36636\,
            ce => 'H',
            sr => \N__31037\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_12_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__25112\,
            in1 => \N__33866\,
            in2 => \N__25079\,
            in3 => \N__24827\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_396_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIANKU4_12_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25321\,
            in2 => \N__24818\,
            in3 => \N__34182\,
            lcout => \b2v_inst11.N_234_N\,
            ltout => \b2v_inst11.N_234_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICO933_12_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100111111"
        )
    port map (
            in0 => \N__25056\,
            in1 => \N__34738\,
            in2 => \N__24815\,
            in3 => \N__33867\,
            lcout => \b2v_inst11.dutycycle_eena_9\,
            ltout => \b2v_inst11.dutycycle_eena_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIHFVH5_12_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__24803\,
            in1 => \N__24787\,
            in2 => \N__24779\,
            in3 => \N__31151\,
            lcout => \b2v_inst11.dutycycleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_11_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__31153\,
            in1 => \N__24767\,
            in2 => \N__24761\,
            in3 => \N__24740\,
            lcout => \b2v_inst11.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36636\,
            ce => 'H',
            sr => \N__31037\
        );

    \b2v_inst11.dutycycle_RNICO933_11_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101011111"
        )
    port map (
            in0 => \N__34739\,
            in1 => \N__33937\,
            in2 => \N__24776\,
            in3 => \N__25111\,
            lcout => \b2v_inst11.dutycycle_eena_7\,
            ltout => \b2v_inst11.dutycycle_eena_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIFCUH5_11_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31152\,
            in1 => \N__24754\,
            in2 => \N__24743\,
            in3 => \N__24739\,
            lcout => \b2v_inst11.dutycycleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIT35D7_13_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010100010"
        )
    port map (
            in0 => \N__31196\,
            in1 => \N__34743\,
            in2 => \N__24875\,
            in3 => \N__27636\,
            lcout => \b2v_inst11.dutycycle_RNIT35D7Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_11_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25036\,
            in1 => \N__25178\,
            in2 => \_gnd_net_\,
            in3 => \N__24676\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100110000"
        )
    port map (
            in0 => \N__33187\,
            in1 => \N__24632\,
            in2 => \N__31377\,
            in3 => \N__35175\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_11_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25177\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_11\,
            ltout => \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24853\,
            in2 => \N__25091\,
            in3 => \N__25035\,
            lcout => \b2v_inst11.N_365\,
            ltout => \b2v_inst11.N_365_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__33165\,
            in1 => \_gnd_net_\,
            in2 => \N__25001\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_366\,
            ltout => \b2v_inst11.N_366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33467\,
            in2 => \N__24998\,
            in3 => \N__33406\,
            lcout => \b2v_inst11.un1_func_state25_6_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIANKU4_13_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101010"
        )
    port map (
            in0 => \N__24986\,
            in1 => \N__25312\,
            in2 => \N__34300\,
            in3 => \N__24951\,
            lcout => \b2v_inst11.N_153_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNILF063_7_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110101010"
        )
    port map (
            in0 => \N__27622\,
            in1 => \N__25479\,
            in2 => \N__25460\,
            in3 => \N__25549\,
            lcout => \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_6_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__33891\,
            in1 => \N__33281\,
            in2 => \_gnd_net_\,
            in3 => \N__29926\,
            lcout => \b2v_inst11.g2_i_a6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__27662\,
            in1 => \N__24854\,
            in2 => \N__33074\,
            in3 => \N__33174\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDUQ02_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001101"
        )
    port map (
            in0 => \N__34623\,
            in1 => \N__27389\,
            in2 => \N__32911\,
            in3 => \N__33280\,
            lcout => \b2v_inst11.func_state_RNIDUQ02Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNIDUQ02Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNILF063_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25325\,
            in3 => \N__25512\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI8H551_7_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__27661\,
            in2 => \N__25553\,
            in3 => \N__25459\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5ELP4_7_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34221\,
            in2 => \N__25271\,
            in3 => \N__25268\,
            lcout => \b2v_inst11.un1_clk_100khz_36_and_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32897\,
            in1 => \N__34602\,
            in2 => \N__34456\,
            in3 => \N__30895\,
            lcout => \b2v_inst11.func_state_RNI8H551Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNILBJP_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__27459\,
            in1 => \N__27528\,
            in2 => \N__29637\,
            in3 => \N__25565\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI9MT83_6_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__25559\,
            in1 => \N__27590\,
            in2 => \N__25262\,
            in3 => \N__34219\,
            lcout => \b2v_inst11.g2_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_6_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27621\,
            lcout => \b2v_inst11.func_state_RNI_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__29891\,
            in1 => \N__30126\,
            in2 => \N__31364\,
            in3 => \N__35135\,
            lcout => \b2v_inst11.N_395\,
            ltout => \b2v_inst11.N_395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_5_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25223\,
            in3 => \N__27580\,
            lcout => \b2v_inst11.dutycycle_RNI_6Z0Z_5\,
            ltout => \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI3NQD_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34016\,
            in1 => \N__32823\,
            in2 => \N__25568\,
            in3 => \N__35062\,
            lcout => \b2v_inst11.g0_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIA70J1_6_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__29886\,
            in1 => \N__34624\,
            in2 => \N__35095\,
            in3 => \N__25538\,
            lcout => \b2v_inst11.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_0_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__25521\,
            in1 => \N__33258\,
            in2 => \_gnd_net_\,
            in3 => \N__25454\,
            lcout => \b2v_inst11.un1_clk_100khz_36_and_i_o3_0_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI8H551_6_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011000100"
        )
    port map (
            in0 => \N__33259\,
            in1 => \N__32874\,
            in2 => \N__34622\,
            in3 => \N__34452\,
            lcout => \b2v_inst11.g0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNILF063_0_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__25522\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25483\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_eena_5_d_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIANKU4_7_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011101110111"
        )
    port map (
            in0 => \N__25455\,
            in1 => \N__33933\,
            in2 => \N__25361\,
            in3 => \N__34277\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_eena_5_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI2IQ6C_7_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011000100"
        )
    port map (
            in0 => \N__34814\,
            in1 => \N__31240\,
            in2 => \N__25358\,
            in3 => \N__25355\,
            lcout => \b2v_inst11.dutycycle_RNI2IQ6CZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI4SIH2_1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__27645\,
            in1 => \N__32875\,
            in2 => \N__33938\,
            in3 => \N__34929\,
            lcout => \b2v_inst11.count_clk_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI34G9_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34453\,
            in1 => \N__29786\,
            in2 => \N__35599\,
            in3 => \N__30820\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_1_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__33260\,
            in1 => \N__30286\,
            in2 => \N__25622\,
            in3 => \N__35031\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__33501\,
            in1 => \N__34040\,
            in2 => \_gnd_net_\,
            in3 => \N__27803\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIICTM5_0_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__25619\,
            in1 => \N__32214\,
            in2 => \N__25610\,
            in3 => \N__28007\,
            lcout => \b2v_inst11.count_clk_en\,
            ltout => \b2v_inst11.count_clk_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIP95D_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__25607\,
            in1 => \N__28025\,
            in2 => \N__25595\,
            in3 => \N__30604\,
            lcout => \b2v_inst11.count_clkZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__25592\,
            in1 => \N__34066\,
            in2 => \N__27809\,
            in3 => \N__33633\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_o_N_329_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__35595\,
            in1 => \N__31427\,
            in2 => \N__25580\,
            in3 => \N__33419\,
            lcout => \b2v_inst11.un1_func_state25_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_1_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35025\,
            in2 => \_gnd_net_\,
            in3 => \N__35594\,
            lcout => \b2v_inst11.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIDQ4A1_7_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__27844\,
            in1 => \_gnd_net_\,
            in2 => \N__33513\,
            in3 => \N__34041\,
            lcout => \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7\,
            ltout => \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_2_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__30914\,
            in1 => \N__25577\,
            in2 => \N__25571\,
            in3 => \N__35026\,
            lcout => \b2v_inst11.un1_func_state25_6_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNINHRI_2_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__25679\,
            in1 => \N__28487\,
            in2 => \N__25637\,
            in3 => \N__30612\,
            lcout => \b2v_inst11.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_2_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25633\,
            lcout => \b2v_inst11.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36656\,
            ce => \N__28583\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIPKSI_3_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__25847\,
            in1 => \N__28485\,
            in2 => \N__30638\,
            in3 => \N__25673\,
            lcout => \b2v_inst11.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25846\,
            lcout => \b2v_inst11.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36656\,
            ce => \N__28583\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIRNTI_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__25667\,
            in1 => \N__28488\,
            in2 => \N__25817\,
            in3 => \N__30613\,
            lcout => \b2v_inst11.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_4_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25813\,
            lcout => \b2v_inst11.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36656\,
            ce => \N__28583\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVTVI_6_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__25661\,
            in1 => \N__28486\,
            in2 => \N__25751\,
            in3 => \N__30611\,
            lcout => \b2v_inst11.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_6_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25747\,
            lcout => \b2v_inst11.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36656\,
            ce => \N__28583\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28169\,
            in2 => \N__28219\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28127\,
            in1 => \N__25654\,
            in2 => \_gnd_net_\,
            in3 => \N__25625\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_1\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28105\,
            in1 => \N__25864\,
            in2 => \_gnd_net_\,
            in3 => \N__25838\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_2\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28128\,
            in1 => \_gnd_net_\,
            in2 => \N__25835\,
            in3 => \N__25805\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_3\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28103\,
            in1 => \N__25802\,
            in2 => \_gnd_net_\,
            in3 => \N__25772\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_4\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28129\,
            in1 => \_gnd_net_\,
            in2 => \N__25769\,
            in3 => \N__25739\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_5\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28104\,
            in1 => \N__28413\,
            in2 => \_gnd_net_\,
            in3 => \N__25736\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_6\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28126\,
            in1 => \N__25733\,
            in2 => \_gnd_net_\,
            in3 => \N__25709\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28097\,
            in1 => \N__25706\,
            in2 => \_gnd_net_\,
            in3 => \N__25685\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28108\,
            in1 => \N__28337\,
            in2 => \_gnd_net_\,
            in3 => \N__25682\,
            lcout => \b2v_inst11.count_clk_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28098\,
            in1 => \N__28351\,
            in2 => \_gnd_net_\,
            in3 => \N__25940\,
            lcout => \b2v_inst11.count_clk_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_10\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28107\,
            in1 => \N__28298\,
            in2 => \_gnd_net_\,
            in3 => \N__25937\,
            lcout => \b2v_inst11.count_clk_1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_11\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28099\,
            in1 => \N__28358\,
            in2 => \_gnd_net_\,
            in3 => \N__25934\,
            lcout => \b2v_inst11.count_clk_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_12\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28106\,
            in1 => \N__25931\,
            in2 => \_gnd_net_\,
            in3 => \N__25910\,
            lcout => \b2v_inst11.count_clk_1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_13\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__25907\,
            in1 => \N__28109\,
            in2 => \_gnd_net_\,
            in3 => \N__25901\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIN3CI_11_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__25889\,
            in1 => \N__25883\,
            in2 => \N__28582\,
            in3 => \N__30574\,
            lcout => \b2v_inst11.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m4_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000100000"
        )
    port map (
            in0 => \N__29247\,
            in1 => \N__29318\,
            in2 => \N__29293\,
            in3 => \N__26133\,
            lcout => OPEN,
            ltout => \b2v_inst36.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNIT62Q_0_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26036\,
            in2 => \N__25871\,
            in3 => \N__30558\,
            lcout => \b2v_inst36.curr_stateZ0Z_0\,
            ltout => \b2v_inst36.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m6_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001010"
        )
    port map (
            in0 => \N__29248\,
            in1 => \N__26132\,
            in2 => \N__26039\,
            in3 => \N__29326\,
            lcout => \b2v_inst36.curr_state_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_0_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101100000001000"
        )
    port map (
            in0 => \N__29284\,
            in1 => \N__29245\,
            in2 => \N__29334\,
            in3 => \N__26152\,
            lcout => \b2v_inst36.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36234\,
            ce => \N__32174\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_1_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101110"
        )
    port map (
            in0 => \N__29246\,
            in1 => \N__29325\,
            in2 => \N__26169\,
            in3 => \N__29285\,
            lcout => \b2v_inst36.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36234\,
            ce => \N__32174\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNIU72Q_1_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26030\,
            in1 => \N__26024\,
            in2 => \_gnd_net_\,
            in3 => \N__30557\,
            lcout => \b2v_inst36.curr_stateZ0Z_1\,
            ltout => \b2v_inst36.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNIRQCA_0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__30559\,
            in1 => \N__29249\,
            in2 => \N__26018\,
            in3 => \N__29282\,
            lcout => \b2v_inst36.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__29283\,
            in1 => \_gnd_net_\,
            in2 => \N__29333\,
            in3 => \N__29244\,
            lcout => \b2v_inst36.DSW_PWROK_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36234\,
            ce => \N__32174\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_8_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26154\,
            in1 => \N__25962\,
            in2 => \N__26003\,
            in3 => \N__28935\,
            lcout => \b2v_inst36.count_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36450\,
            ce => \N__29148\,
            sr => \N__28982\
        );

    \b2v_inst36.count_RNIPT1I1_8_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29106\,
            in1 => \N__25982\,
            in2 => \_gnd_net_\,
            in3 => \N__25976\,
            lcout => \b2v_inst36.countZ0Z_8\,
            ltout => \b2v_inst36.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI4VQN1_0_10_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__29149\,
            in1 => \N__26075\,
            in2 => \N__25943\,
            in3 => \N__26213\,
            lcout => OPEN,
            ltout => \b2v_inst36.un12_clk_100khz_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNILGID6_1_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26255\,
            in1 => \N__26249\,
            in2 => \N__26243\,
            in3 => \N__26240\,
            lcout => OPEN,
            ltout => \b2v_inst36.un12_clk_100khz_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI0RKG9_6_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26228\,
            in1 => \N__26342\,
            in2 => \N__26219\,
            in3 => \N__26303\,
            lcout => \b2v_inst36.N_1_i\,
            ltout => \b2v_inst36.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__28936\,
            in1 => \N__26200\,
            in2 => \N__26216\,
            in3 => \N__26189\,
            lcout => \b2v_inst36.count_rst_4\,
            ltout => \b2v_inst36.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI4VQN1_10_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26074\,
            in2 => \N__26207\,
            in3 => \N__29107\,
            lcout => \b2v_inst36.un2_count_1_axb_10\,
            ltout => \b2v_inst36.un2_count_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_10_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__28934\,
            in1 => \N__26188\,
            in2 => \N__26177\,
            in3 => \N__26155\,
            lcout => \b2v_inst36.count_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36450\,
            ce => \N__29148\,
            sr => \N__28982\
        );

    \b2v_inst36.count_4_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26060\,
            lcout => \b2v_inst36.count_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36244\,
            ce => \N__29132\,
            sr => \N__28962\
        );

    \b2v_inst36.count_RNICQ3V_6_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26350\,
            in1 => \N__29120\,
            in2 => \_gnd_net_\,
            in3 => \N__26367\,
            lcout => \b2v_inst36.un2_count_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_6_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26368\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36244\,
            ce => \N__29132\,
            sr => \N__28962\
        );

    \b2v_inst36.count_RNIHHTH1_4_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26059\,
            in1 => \N__29119\,
            in2 => \_gnd_net_\,
            in3 => \N__26051\,
            lcout => \b2v_inst36.countZ0Z_4\,
            ltout => \b2v_inst36.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNICQ3V_0_6_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__29122\,
            in1 => \N__26369\,
            in2 => \N__26354\,
            in3 => \N__26351\,
            lcout => \b2v_inst36.un12_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIPRQ41_12_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26330\,
            in1 => \N__29121\,
            in2 => \_gnd_net_\,
            in3 => \N__26316\,
            lcout => \b2v_inst36.un2_count_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_12_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26317\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36244\,
            ce => \N__29132\,
            sr => \N__28962\
        );

    \b2v_inst36.count_RNIPRQ41_0_12_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010001"
        )
    port map (
            in0 => \N__26329\,
            in1 => \N__29189\,
            in2 => \N__26321\,
            in3 => \N__29133\,
            lcout => \b2v_inst36.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_3_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26575\,
            lcout => \b2v_inst5.count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36356\,
            ce => \N__26863\,
            sr => \N__27302\
        );

    \b2v_inst5.count_RNIBN4H3_1_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26282\,
            in1 => \N__26297\,
            in2 => \_gnd_net_\,
            in3 => \N__26825\,
            lcout => \b2v_inst5.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_1_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36356\,
            ce => \N__26863\,
            sr => \N__27302\
        );

    \b2v_inst5.count_RNIDQ5H3_2_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26276\,
            in1 => \N__26261\,
            in2 => \_gnd_net_\,
            in3 => \N__26826\,
            lcout => \b2v_inst5.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_2_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26275\,
            lcout => \b2v_inst5.count_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36356\,
            ce => \N__26863\,
            sr => \N__27302\
        );

    \b2v_inst5.count_RNIFT6H3_3_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26576\,
            in1 => \N__26561\,
            in2 => \_gnd_net_\,
            in3 => \N__26827\,
            lcout => \b2v_inst5.countZ0Z_3\,
            ltout => \b2v_inst5.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI_1_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__26540\,
            in1 => \N__26515\,
            in2 => \N__26501\,
            in3 => \N__26494\,
            lcout => \b2v_inst5.un12_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIJ39H3_5_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26903\,
            in1 => \N__26882\,
            in2 => \_gnd_net_\,
            in3 => \N__26828\,
            lcout => \b2v_inst5.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI7BCA2_0_10_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__26633\,
            in1 => \N__26815\,
            in2 => \N__26455\,
            in3 => \N__27015\,
            lcout => OPEN,
            ltout => \b2v_inst5.un12_clk_100khz_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI870S9_8_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26480\,
            in1 => \N__26471\,
            in2 => \N__26462\,
            in3 => \N__26375\,
            lcout => \b2v_inst5.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI7BCA2_10_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26632\,
            in1 => \_gnd_net_\,
            in2 => \N__26456\,
            in3 => \N__26813\,
            lcout => \b2v_inst5.un2_count_1_axb_10\,
            ltout => \b2v_inst5.un2_count_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_10_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__26666\,
            in1 => \N__26975\,
            in2 => \N__26459\,
            in3 => \N__27330\,
            lcout => \b2v_inst5.count_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36350\,
            ce => \N__26820\,
            sr => \N__27329\
        );

    \b2v_inst5.count_RNI3QEK5_11_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__26441\,
            in1 => \N__26425\,
            in2 => \N__26411\,
            in3 => \N__26402\,
            lcout => \b2v_inst5.un12_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIRFDH3_9_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26814\,
            in1 => \_gnd_net_\,
            in2 => \N__26675\,
            in3 => \N__26909\,
            lcout => \b2v_inst5.countZ0Z_9\,
            ltout => \b2v_inst5.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_9_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__26974\,
            in1 => \N__27293\,
            in2 => \N__26678\,
            in3 => \N__26999\,
            lcout => \b2v_inst5.count_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36350\,
            ce => \N__26820\,
            sr => \N__27329\
        );

    \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__26665\,
            in1 => \N__26973\,
            in2 => \N__27325\,
            in3 => \N__26647\,
            lcout => \b2v_inst5.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIKEUB2_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32248\,
            in2 => \N__32237\,
            in3 => \N__30391\,
            lcout => \b2v_inst5.curr_stateZ0Z_1\,
            ltout => \b2v_inst5.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26624\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.curr_state_RNIZ0Z_1\,
            ltout => \b2v_inst5.curr_state_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIRH7S1_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__32986\,
            in1 => \N__27357\,
            in2 => \N__26621\,
            in3 => \N__31124\,
            lcout => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\,
            ltout => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNILCEN3_15_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26600\,
            in1 => \_gnd_net_\,
            in2 => \N__26618\,
            in3 => \N__26588\,
            lcout => \b2v_inst5.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_15_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26599\,
            lcout => \b2v_inst5.count_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36360\,
            ce => \N__26819\,
            sr => \N__27331\
        );

    \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26582\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26938\,
            lcout => \N_413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__27019\,
            in1 => \N__26998\,
            in2 => \N__26980\,
            in3 => \N__27213\,
            lcout => \b2v_inst5.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_5_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26902\,
            lcout => \b2v_inst5.count_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36360\,
            ce => \N__26819\,
            sr => \N__27331\
        );

    \b2v_inst5.curr_state_RNI65HI_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26696\,
            in2 => \N__30602\,
            in3 => \N__26717\,
            lcout => \b2v_inst5.curr_stateZ0Z_0\,
            ltout => \b2v_inst5.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m6_i_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__32988\,
            in1 => \N__27382\,
            in2 => \N__26720\,
            in3 => \N__26707\,
            lcout => \b2v_inst5.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27381\,
            in1 => \N__32987\,
            in2 => \_gnd_net_\,
            in3 => \N__26690\,
            lcout => \RSMRSTn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36448\,
            ce => \N__32176\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__27358\,
            in1 => \N__27513\,
            in2 => \_gnd_net_\,
            in3 => \N__26706\,
            lcout => \b2v_inst5.m4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI65HI_0_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26689\,
            lcout => \b2v_inst5.N_2898_i\,
            ltout => \b2v_inst5.N_2898_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27512\,
            in2 => \N__26711\,
            in3 => \N__26708\,
            lcout => \b2v_inst5.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36448\,
            ce => \N__32176\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNID8DP1_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32990\,
            in1 => \N__27373\,
            in2 => \_gnd_net_\,
            in3 => \N__26688\,
            lcout => \curr_state_RNID8DP1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIVF6A1_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32989\,
            in1 => \N__27383\,
            in2 => \N__27362\,
            in3 => \N__30420\,
            lcout => \b2v_inst5.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_8_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33385\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_172_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI5DLR_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__34615\,
            in1 => \N__32910\,
            in2 => \_gnd_net_\,
            in3 => \N__35096\,
            lcout => \b2v_inst11.un1_clk_100khz_2_i_o3_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111011111"
        )
    port map (
            in0 => \N__34619\,
            in1 => \N__29623\,
            in2 => \N__27445\,
            in3 => \N__27495\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_6_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33384\,
            in2 => \_gnd_net_\,
            in3 => \N__33293\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111111"
        )
    port map (
            in0 => \N__28246\,
            in1 => \N__33898\,
            in2 => \N__27056\,
            in3 => \N__34052\,
            lcout => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_RNI8DFE_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27046\,
            in1 => \_gnd_net_\,
            in2 => \N__27514\,
            in3 => \N__27432\,
            lcout => rsmrstn,
            ltout => \rsmrstn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__34405\,
            in1 => \N__30309\,
            in2 => \N__27053\,
            in3 => \N__29624\,
            lcout => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__27499\,
            in1 => \N__29570\,
            in2 => \N__27050\,
            in3 => \N__27433\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__32907\,
            in1 => \N__34614\,
            in2 => \_gnd_net_\,
            in3 => \N__34181\,
            lcout => \b2v_inst11.N_168\,
            ltout => \b2v_inst11.N_168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__30515\,
            in1 => \N__32908\,
            in2 => \N__27536\,
            in3 => \N__34625\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.VCCST_EN_i_0_o3_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101111111"
        )
    port map (
            in0 => \N__32906\,
            in1 => \N__30514\,
            in2 => \N__27527\,
            in3 => \N__27458\,
            lcout => \VCCST_EN_i_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIDQ4A1_6_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111111"
        )
    port map (
            in0 => \N__33477\,
            in1 => \N__27573\,
            in2 => \N__27982\,
            in3 => \N__33079\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_clk_RNIDQ4A1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIQK9K2_6_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33407\,
            in2 => \N__27407\,
            in3 => \N__27404\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIH3DN3_6_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__34884\,
            in1 => \_gnd_net_\,
            in2 => \N__27398\,
            in3 => \N__34432\,
            lcout => \b2v_inst11.N_186_i\,
            ltout => \b2v_inst11.N_186_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIN1E71_2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__33098\,
            in1 => \N__32909\,
            in2 => \N__27395\,
            in3 => \N__34883\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_115_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAEUL3_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31211\,
            in2 => \N__27392\,
            in3 => \N__34737\,
            lcout => \b2v_inst11.dutycycle_RNIAEUL3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_0_1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__34601\,
            in1 => \N__32905\,
            in2 => \N__34454\,
            in3 => \N__35094\,
            lcout => \b2v_inst11.N_381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_6_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29797\,
            in1 => \N__33304\,
            in2 => \N__27785\,
            in3 => \N__29942\,
            lcout => \b2v_inst11.g0_i_a7_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIUCAD1_0_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27740\,
            lcout => \b2v_inst16.N_268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__34014\,
            in1 => \N__30893\,
            in2 => \N__27974\,
            in3 => \N__27668\,
            lcout => \b2v_inst11.N_159\,
            ltout => \b2v_inst11.N_159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_4_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27653\,
            in3 => \N__27574\,
            lcout => \b2v_inst11.N_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI2MQD_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34600\,
            in1 => \N__27579\,
            in2 => \N__27975\,
            in3 => \N__30894\,
            lcout => \b2v_inst11.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_ss0_i_0_a2_2_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__32904\,
            in1 => \N__34599\,
            in2 => \_gnd_net_\,
            in3 => \N__34220\,
            lcout => \b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30778\,
            in1 => \N__34015\,
            in2 => \N__35108\,
            in3 => \N__35600\,
            lcout => \b2v_inst11.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__33716\,
            in1 => \N__31312\,
            in2 => \N__30144\,
            in3 => \N__29890\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_0\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30777\,
            in1 => \N__27584\,
            in2 => \N__27539\,
            in3 => \N__30896\,
            lcout => \b2v_inst11.N_406\,
            ltout => \b2v_inst11.N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVT4P1_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34748\,
            in2 => \N__27872\,
            in3 => \N__35084\,
            lcout => \b2v_inst11.func_state_1_m2_ns_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__27869\,
            in1 => \N__28016\,
            in2 => \N__33632\,
            in3 => \N__28284\,
            lcout => \b2v_inst11.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_en_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32824\,
            in2 => \N__32224\,
            in3 => \N__34894\,
            lcout => \b2v_inst11.func_state_enZ0\,
            ltout => \b2v_inst11.func_state_enZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDHTPG_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__27868\,
            in1 => \N__33618\,
            in2 => \N__27860\,
            in3 => \N__28015\,
            lcout => \b2v_inst11.func_state\,
            ltout => \b2v_inst11.func_state_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27857\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_2946_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI5DLR_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__30290\,
            in1 => \N__35030\,
            in2 => \N__27854\,
            in3 => \N__30883\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINIV94_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27807\,
            in1 => \N__27823\,
            in2 => \N__27833\,
            in3 => \N__27830\,
            lcout => \b2v_inst11.func_state_RNINIV94_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF1Q43_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011101110111"
        )
    port map (
            in0 => \N__27824\,
            in1 => \N__27808\,
            in2 => \N__30307\,
            in3 => \N__30884\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m2_ns_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINCPR4_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__27928\,
            in1 => \N__30841\,
            in2 => \N__27788\,
            in3 => \N__35586\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m2_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIPBBTD_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110001011"
        )
    port map (
            in0 => \N__30761\,
            in1 => \N__27884\,
            in2 => \N__28019\,
            in3 => \N__27927\,
            lcout => \b2v_inst11.func_state_1_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNID7Q51_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000100"
        )
    port map (
            in0 => \N__30882\,
            in1 => \N__34085\,
            in2 => \N__35072\,
            in3 => \N__35584\,
            lcout => \b2v_inst11.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__34433\,
            in1 => \N__34201\,
            in2 => \N__30306\,
            in3 => \N__30623\,
            lcout => \b2v_inst11.N_382\,
            ltout => \b2v_inst11.N_382_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI794G3_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__28001\,
            in1 => \N__35585\,
            in2 => \N__27992\,
            in3 => \N__34048\,
            lcout => \b2v_inst11.func_state_1_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIHJNV7_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__27989\,
            in1 => \N__31239\,
            in2 => \N__27983\,
            in3 => \N__27944\,
            lcout => \b2v_inst11.dutycycle_RNIHJNV7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI98MHC_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001111"
        )
    port map (
            in0 => \N__30757\,
            in1 => \N__27932\,
            in2 => \N__27914\,
            in3 => \N__27883\,
            lcout => \b2v_inst11.func_state_1_m2_1\,
            ltout => \b2v_inst11.func_state_1_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIUE8EF_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__28258\,
            in1 => \N__33617\,
            in2 => \N__27905\,
            in3 => \N__28285\,
            lcout => \b2v_inst11.func_stateZ0Z_0\,
            ltout => \b2v_inst11.func_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI57FD1_0_1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30308\,
            in1 => \N__30603\,
            in2 => \N__27902\,
            in3 => \N__34200\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIHVOG4_1_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__28229\,
            in1 => \N__27899\,
            in2 => \N__27887\,
            in3 => \N__34747\,
            lcout => \b2v_inst11.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__28286\,
            in1 => \N__28268\,
            in2 => \N__28262\,
            in3 => \N__33622\,
            lcout => \b2v_inst11.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__33418\,
            in1 => \N__28247\,
            in2 => \_gnd_net_\,
            in3 => \N__35083\,
            lcout => \b2v_inst11.func_state_1_m2s2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28090\,
            in1 => \N__28223\,
            in2 => \_gnd_net_\,
            in3 => \N__28155\,
            lcout => \b2v_inst11.count_clk_RNIZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28089\,
            lcout => \b2v_inst11.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36657\,
            ce => \N__28572\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI8F1AB_2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35681\,
            in1 => \N__35886\,
            in2 => \_gnd_net_\,
            in3 => \N__35699\,
            lcout => \b2v_inst11.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIAI2AB_3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35887\,
            in1 => \N__36728\,
            in2 => \_gnd_net_\,
            in3 => \N__36746\,
            lcout => \b2v_inst11.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNICA5EB_13_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35711\,
            in1 => \N__35890\,
            in2 => \_gnd_net_\,
            in3 => \N__35726\,
            lcout => \b2v_inst11.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNICL3AB_4_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35888\,
            in1 => \N__36701\,
            in2 => \_gnd_net_\,
            in3 => \N__36719\,
            lcout => \b2v_inst11.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIED6EB_14_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31439\,
            in1 => \N__35891\,
            in2 => \_gnd_net_\,
            in3 => \N__31454\,
            lcout => \b2v_inst11.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIEO4AB_5_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35889\,
            in1 => \N__36674\,
            in2 => \_gnd_net_\,
            in3 => \N__36692\,
            lcout => \b2v_inst11.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_10_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28369\,
            lcout => \b2v_inst11.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36552\,
            ce => \N__28538\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_12_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28315\,
            lcout => \b2v_inst11.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36552\,
            ce => \N__28538\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI111J_7_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__28385\,
            in1 => \N__28554\,
            in2 => \N__28397\,
            in3 => \N__30680\,
            lcout => \b2v_inst11.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_7_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28393\,
            lcout => \b2v_inst11.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36541\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIEN0E_10_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__28556\,
            in1 => \N__28379\,
            in2 => \N__28373\,
            in3 => \N__30681\,
            lcout => \b2v_inst11.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIR9EI_13_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__28598\,
            in1 => \N__28589\,
            in2 => \N__30725\,
            in3 => \N__28558\,
            lcout => \b2v_inst11.count_clkZ0Z_13\,
            ltout => \b2v_inst11.count_clkZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_10_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28297\,
            in1 => \N__28352\,
            in2 => \N__28340\,
            in3 => \N__28336\,
            lcout => \b2v_inst11.un2_count_clk_17_0_o2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIP6DI_12_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__28316\,
            in1 => \N__28304\,
            in2 => \N__30724\,
            in3 => \N__28557\,
            lcout => \b2v_inst11.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_13_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28597\,
            lcout => \b2v_inst11.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36541\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32102\,
            in2 => \N__32687\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_1_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_RNID98I1_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32616\,
            in1 => \N__31574\,
            in2 => \_gnd_net_\,
            in3 => \N__28445\,
            lcout => \b2v_inst6.count_rst_12\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_1\,
            carryout => \b2v_inst6.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31615\,
            in3 => \N__28442\,
            lcout => \b2v_inst6.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_2\,
            carryout => \b2v_inst6.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31495\,
            in3 => \N__28439\,
            lcout => \b2v_inst6.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_3\,
            carryout => \b2v_inst6.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32015\,
            in2 => \_gnd_net_\,
            in3 => \N__28436\,
            lcout => \b2v_inst6.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_4\,
            carryout => \b2v_inst6.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28628\,
            in2 => \_gnd_net_\,
            in3 => \N__28433\,
            lcout => \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_5\,
            carryout => \b2v_inst6.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28682\,
            in2 => \_gnd_net_\,
            in3 => \N__28430\,
            lcout => \b2v_inst6.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_6\,
            carryout => \b2v_inst6.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32455\,
            in2 => \_gnd_net_\,
            in3 => \N__28427\,
            lcout => \b2v_inst6.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_7\,
            carryout => \b2v_inst6.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29425\,
            in2 => \_gnd_net_\,
            in3 => \N__28619\,
            lcout => \b2v_inst6.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_9_c_RNILPGI1_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32617\,
            in1 => \N__28775\,
            in2 => \_gnd_net_\,
            in3 => \N__28616\,
            lcout => \b2v_inst6.count_rst_4\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_9\,
            carryout => \b2v_inst6.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31847\,
            in2 => \_gnd_net_\,
            in3 => \N__28613\,
            lcout => \b2v_inst6.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_10\,
            carryout => \b2v_inst6.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_11_c_RNIU1QP1_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32618\,
            in1 => \N__31754\,
            in2 => \_gnd_net_\,
            in3 => \N__28610\,
            lcout => \b2v_inst6.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_11\,
            carryout => \b2v_inst6.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_12_c_RNIV3RP1_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32620\,
            in1 => \N__31682\,
            in2 => \_gnd_net_\,
            in3 => \N__28607\,
            lcout => \b2v_inst6.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_12\,
            carryout => \b2v_inst6.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_13_c_RNI06SP1_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32619\,
            in1 => \N__31787\,
            in2 => \_gnd_net_\,
            in3 => \N__28604\,
            lcout => \b2v_inst6.un2_count_1_cry_13_c_RNI06SPZ0Z1\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_13\,
            carryout => \b2v_inst6.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_14_c_RNI18TP1_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32621\,
            in1 => \N__28691\,
            in2 => \_gnd_net_\,
            in3 => \N__28601\,
            lcout => \b2v_inst6.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_10_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28794\,
            lcout => \b2v_inst6.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36510\,
            ce => \N__32422\,
            sr => \N__32651\
        );

    \b2v_inst6.count_15_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28700\,
            lcout => \b2v_inst6.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36556\,
            ce => \N__32429\,
            sr => \N__32607\
        );

    \b2v_inst6.count_13_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31712\,
            lcout => \b2v_inst6.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36556\,
            ce => \N__32429\,
            sr => \N__32607\
        );

    \b2v_inst6.count_RNIT5A54_15_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32361\,
            in1 => \N__28706\,
            in2 => \_gnd_net_\,
            in3 => \N__28699\,
            lcout => \b2v_inst6.countZ0Z_15\,
            ltout => \b2v_inst6.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIPV754_0_13_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__31696\,
            in1 => \N__32362\,
            in2 => \N__28685\,
            in3 => \N__31711\,
            lcout => \b2v_inst6.count_1_i_a3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_7_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__28681\,
            in1 => \N__31942\,
            in2 => \N__28667\,
            in3 => \N__32615\,
            lcout => \b2v_inst6.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36556\,
            ce => \N__32429\,
            sr => \N__32607\
        );

    \b2v_inst6.count_RNIV0AS3_7_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28642\,
            in1 => \N__32360\,
            in2 => \_gnd_net_\,
            in3 => \N__28649\,
            lcout => \b2v_inst6.un2_count_1_axb_7\,
            ltout => \b2v_inst6.un2_count_1_axb_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_6_c_RNIIJDI1_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__28663\,
            in1 => \N__31941\,
            in2 => \N__28652\,
            in3 => \N__32614\,
            lcout => \b2v_inst6.count_rst_7\,
            ltout => \b2v_inst6.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIV0AS3_0_7_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__28643\,
            in1 => \N__32363\,
            in2 => \N__28634\,
            in3 => \N__32014\,
            lcout => \b2v_inst6.count_1_i_a3_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIALQ32_1_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__29729\,
            in1 => \N__32547\,
            in2 => \_gnd_net_\,
            in3 => \N__31209\,
            lcout => \b2v_inst6.count_en\,
            ltout => \b2v_inst6.count_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNITT8S3_6_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__32548\,
            in1 => \N__31655\,
            in2 => \N__28631\,
            in3 => \N__31672\,
            lcout => \b2v_inst6.countZ0Z_6\,
            ltout => \b2v_inst6.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNICITT3_0_10_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__32367\,
            in1 => \N__28796\,
            in2 => \N__29348\,
            in3 => \N__28808\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_1_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI3F438_12_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000110000"
        )
    port map (
            in0 => \N__31748\,
            in1 => \N__31730\,
            in2 => \N__29345\,
            in3 => \N__32368\,
            lcout => \b2v_inst6.count_1_i_a3_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNINSDS_0_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__29341\,
            in1 => \N__29292\,
            in2 => \N__29243\,
            in3 => \N__31210\,
            lcout => \b2v_inst36.curr_state_RNINSDSZ0Z_0\,
            ltout => \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIR03I1_9_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29168\,
            in2 => \N__29192\,
            in3 => \N__29156\,
            lcout => \b2v_inst36.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_9_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36402\,
            ce => \N__29126\,
            sr => \N__28972\
        );

    \b2v_inst6.count_RNICITT3_10_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28807\,
            in1 => \N__28795\,
            in2 => \_gnd_net_\,
            in3 => \N__32366\,
            lcout => \b2v_inst6.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un8_rsmrst_pwrgd_4_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28766\,
            in1 => \N__28751\,
            in2 => \N__28739\,
            in3 => \N__28718\,
            lcout => \SYNTHESIZED_WIRE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_8_c_RNIKNFI1_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__32542\,
            in1 => \N__29407\,
            in2 => \N__29426\,
            in3 => \N__31954\,
            lcout => \b2v_inst6.count_rst_5\,
            ltout => \b2v_inst6.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI37CS3_9_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32365\,
            in1 => \_gnd_net_\,
            in2 => \N__28709\,
            in3 => \N__32467\,
            lcout => \b2v_inst6.un2_count_1_axb_9\,
            ltout => \b2v_inst6.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_9_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__32649\,
            in1 => \N__29408\,
            in2 => \N__29396\,
            in3 => \N__31955\,
            lcout => \b2v_inst6.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36568\,
            ce => \N__32428\,
            sr => \N__32648\
        );

    \b2v_inst6.un2_count_1_cry_7_c_RNIJLEI1_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__32451\,
            in1 => \N__31952\,
            in2 => \N__29390\,
            in3 => \N__32541\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI14BS3_8_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__29372\,
            in1 => \_gnd_net_\,
            in2 => \N__29393\,
            in3 => \N__32364\,
            lcout => \b2v_inst6.countZ0Z_8\,
            ltout => \b2v_inst6.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_8_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__29389\,
            in1 => \N__31953\,
            in2 => \N__29375\,
            in3 => \N__32543\,
            lcout => \b2v_inst6.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36568\,
            ce => \N__32428\,
            sr => \N__32648\
        );

    \b2v_inst6.curr_state_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29354\,
            lcout => \b2v_inst6.curr_state_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36635\,
            ce => \N__32183\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__31951\,
            in1 => \N__29514\,
            in2 => \N__29704\,
            in3 => \N__29537\,
            lcout => \b2v_inst6.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36635\,
            ce => \N__32183\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m4_0_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__29515\,
            in1 => \N__29535\,
            in2 => \N__29705\,
            in3 => \N__31949\,
            lcout => OPEN,
            ltout => \b2v_inst6.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI5DHS1_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29363\,
            in2 => \N__29357\,
            in3 => \N__30597\,
            lcout => \b2v_inst6.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m6_i_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__29536\,
            in1 => \N__31950\,
            in2 => \_gnd_net_\,
            in3 => \N__29725\,
            lcout => \b2v_inst6.N_42\,
            ltout => \b2v_inst6.N_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI8KCH_1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29546\,
            in2 => \N__29540\,
            in3 => \N__30595\,
            lcout => \b2v_inst6.curr_stateZ0Z_1\,
            ltout => \b2v_inst6.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29522\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.N_3053_i\,
            ltout => \b2v_inst6.N_3053_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIM6FE1_1_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29516\,
            in1 => \N__29756\,
            in2 => \N__29519\,
            in3 => \N__30596\,
            lcout => \b2v_inst6.curr_state_RNIM6FE1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29451\,
            lcout => \b2v_inst6.N_3034_i\,
            ltout => \b2v_inst6.N_3034_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIUP4B1_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29436\,
            in2 => \N__29501\,
            in3 => \N__29754\,
            lcout => \b2v_inst6.N_276_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIUP4B1_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__29755\,
            in1 => \_gnd_net_\,
            in2 => \N__29441\,
            in3 => \N__29452\,
            lcout => \b2v_inst6.curr_state_RNIUP4B1Z0Z_0\,
            ltout => \b2v_inst6.curr_state_RNIUP4B1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU8MF3_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__29680\,
            in1 => \N__29713\,
            in2 => \N__29498\,
            in3 => \N__32215\,
            lcout => OPEN,
            ltout => \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29495\,
            in3 => \N__34927\,
            lcout => \N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__29453\,
            in1 => \N__29440\,
            in2 => \_gnd_net_\,
            in3 => \N__29753\,
            lcout => \N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__29714\,
            in1 => \N__29697\,
            in2 => \N__32225\,
            in3 => \N__29681\,
            lcout => \b2v_inst6.delayed_vccin_vccinaux_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34061\,
            in2 => \_gnd_net_\,
            in3 => \N__35109\,
            lcout => \b2v_inst11.N_172\,
            ltout => \b2v_inst11.N_172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_3_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001010"
        )
    port map (
            in0 => \N__33078\,
            in1 => \N__29672\,
            in2 => \N__29657\,
            in3 => \N__33311\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIKAJP_6_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__29654\,
            in1 => \N__33377\,
            in2 => \N__29642\,
            in3 => \N__34919\,
            lcout => \b2v_inst11.g0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINGLA1_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__35110\,
            in1 => \N__30047\,
            in2 => \N__30326\,
            in3 => \N__29636\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI4KE12_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__29585\,
            in1 => \N__34495\,
            in2 => \N__29573\,
            in3 => \N__35111\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32896\,
            in2 => \_gnd_net_\,
            in3 => \N__34494\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_0_o3_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__29561\,
            in1 => \N__31332\,
            in2 => \N__33314\,
            in3 => \N__30143\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.N_224_i_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__34421\,
            in1 => \N__34241\,
            in2 => \N__30325\,
            in3 => \N__30598\,
            lcout => \b2v_inst11.N_224_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI34G9_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34422\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34064\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNII5M67_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__29980\,
            in1 => \N__30007\,
            in2 => \N__30020\,
            in3 => \N__29995\,
            lcout => \b2v_inst11.dutycycleZ0Z_2\,
            ltout => \b2v_inst11.dutycycleZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30041\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_2_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__30019\,
            in1 => \N__30008\,
            in2 => \N__29984\,
            in3 => \N__29996\,
            lcout => \b2v_inst11.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36207\,
            ce => 'H',
            sr => \N__30984\
        );

    \b2v_inst11.dutycycle_RNI_0_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29962\,
            in1 => \N__29809\,
            in2 => \N__30166\,
            in3 => \N__31310\,
            lcout => \b2v_inst11.N_293_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31311\,
            in1 => \N__29963\,
            in2 => \N__29813\,
            in3 => \N__30142\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_2_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34059\,
            in2 => \_gnd_net_\,
            in3 => \N__35091\,
            lcout => \b2v_inst11.func_state_RNI_2Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIN1E71_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110001"
        )
    port map (
            in0 => \N__32895\,
            in1 => \N__34931\,
            in2 => \N__29771\,
            in3 => \N__29768\,
            lcout => \b2v_inst11.N_119_f0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010010001"
        )
    port map (
            in0 => \N__35583\,
            in1 => \N__34060\,
            in2 => \N__30785\,
            in3 => \N__35093\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_ss0_i_0_o3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIHVOG4_0_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111101"
        )
    port map (
            in0 => \N__34810\,
            in1 => \N__30230\,
            in2 => \N__30764\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI57FD1_1_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__34250\,
            in1 => \N__35092\,
            in2 => \N__30705\,
            in3 => \N__30324\,
            lcout => \b2v_inst11.N_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIN52J1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110001"
        )
    port map (
            in0 => \N__35105\,
            in1 => \N__30224\,
            in2 => \N__33515\,
            in3 => \N__30898\,
            lcout => \b2v_inst11.dutycycle_1_0_1\,
            ltout => \b2v_inst11.dutycycle_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIB6O76_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__31236\,
            in1 => \N__31051\,
            in2 => \N__30209\,
            in3 => \N__31256\,
            lcout => \b2v_inst11.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011111000"
        )
    port map (
            in0 => \N__30206\,
            in1 => \N__31238\,
            in2 => \N__30200\,
            in3 => \N__30056\,
            lcout => \b2v_inst11.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36416\,
            ce => 'H',
            sr => \N__31036\
        );

    \b2v_inst11.dutycycle_RNIAA6Q3_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111101"
        )
    port map (
            in0 => \N__34808\,
            in1 => \N__30115\,
            in2 => \N__34938\,
            in3 => \N__31387\,
            lcout => \b2v_inst11.dutycycle_eena\,
            ltout => \b2v_inst11.dutycycle_eena_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI0QQU5_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__30196\,
            in1 => \N__31235\,
            in2 => \N__30188\,
            in3 => \N__30055\,
            lcout => \b2v_inst11.dutycycleZ0Z_0\,
            ltout => \b2v_inst11.dutycycleZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__30897\,
            in1 => \N__33509\,
            in2 => \N__30059\,
            in3 => \N__35104\,
            lcout => \b2v_inst11.dutycycle_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAA6Q3_1_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100111011"
        )
    port map (
            in0 => \N__34926\,
            in1 => \N__34809\,
            in2 => \N__31391\,
            in3 => \N__31309\,
            lcout => \b2v_inst11.dutycycle_eena_0\,
            ltout => \b2v_inst11.dutycycle_eena_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__31237\,
            in1 => \N__31061\,
            in2 => \N__31055\,
            in3 => \N__31052\,
            lcout => \b2v_inst11.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36416\,
            ce => 'H',
            sr => \N__31036\
        );

    \b2v_inst11.count_off_RNIL5413_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35326\,
            in2 => \_gnd_net_\,
            in3 => \N__35271\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_off_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI8BS7B_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35231\,
            in2 => \N__30917\,
            in3 => \N__35929\,
            lcout => \b2v_inst11.count_offZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30848\,
            in1 => \N__31420\,
            in2 => \_gnd_net_\,
            in3 => \N__30827\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_330_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30902\,
            lcout => \b2v_inst11.func_state_RNI_0Z0Z_0\,
            ltout => \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8BVM1_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30842\,
            in1 => \N__30826\,
            in2 => \N__30803\,
            in3 => \N__35577\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIL5413_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__35107\,
            in1 => \N__35587\,
            in2 => \N__30800\,
            in3 => \N__30797\,
            lcout => \b2v_inst11.N_125\,
            ltout => \b2v_inst11.N_125_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIL5413_1_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35362\,
            in2 => \N__31430\,
            in3 => \N__35325\,
            lcout => \b2v_inst11.count_off_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__34493\,
            in1 => \N__32894\,
            in2 => \N__34445\,
            in3 => \N__34301\,
            lcout => \b2v_inst11.N_382_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35327\,
            in2 => \N__35363\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_RNIJ7933_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35272\,
            in1 => \N__35626\,
            in2 => \_gnd_net_\,
            in3 => \N__31409\,
            lcout => \b2v_inst11.count_off_1_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_1\,
            carryout => \b2v_inst11.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_2_c_RNIK9A33_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35276\,
            in1 => \N__35416\,
            in2 => \_gnd_net_\,
            in3 => \N__31406\,
            lcout => \b2v_inst11.count_off_1_3\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_2\,
            carryout => \b2v_inst11.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_3_c_RNILBB33_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35273\,
            in1 => \N__35392\,
            in2 => \_gnd_net_\,
            in3 => \N__31403\,
            lcout => \b2v_inst11.count_off_1_4\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_3\,
            carryout => \b2v_inst11.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_4_c_RNIMDC33_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35277\,
            in1 => \N__35653\,
            in2 => \_gnd_net_\,
            in3 => \N__31400\,
            lcout => \b2v_inst11.count_off_1_5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_4\,
            carryout => \b2v_inst11.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_5_c_RNINFD33_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35274\,
            in1 => \N__35671\,
            in2 => \_gnd_net_\,
            in3 => \N__31397\,
            lcout => \b2v_inst11.count_off_1_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_5\,
            carryout => \b2v_inst11.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_6_c_RNIOHE33_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35278\,
            in1 => \N__35458\,
            in2 => \_gnd_net_\,
            in3 => \N__31394\,
            lcout => \b2v_inst11.count_off_1_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_6\,
            carryout => \b2v_inst11.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_7_c_RNIPJF33_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35275\,
            in1 => \N__35437\,
            in2 => \_gnd_net_\,
            in3 => \N__31478\,
            lcout => \b2v_inst11.count_off_1_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_7\,
            carryout => \b2v_inst11.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_8_c_RNIQLG33_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35297\,
            in1 => \N__35210\,
            in2 => \_gnd_net_\,
            in3 => \N__31475\,
            lcout => \b2v_inst11.count_off_1_9\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_9_c_RNIRNH33_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__35301\,
            in1 => \_gnd_net_\,
            in2 => \N__35813\,
            in3 => \N__31472\,
            lcout => \b2v_inst11.count_off_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_9\,
            carryout => \b2v_inst11.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_10_c_RNI35P63_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35298\,
            in1 => \N__35782\,
            in2 => \_gnd_net_\,
            in3 => \N__31469\,
            lcout => \b2v_inst11.count_off_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_10\,
            carryout => \b2v_inst11.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_11_c_RNI47Q63_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35303\,
            in1 => \N__35756\,
            in2 => \_gnd_net_\,
            in3 => \N__31466\,
            lcout => \b2v_inst11.count_off_1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_11\,
            carryout => \b2v_inst11.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_12_c_RNI59R63_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35299\,
            in1 => \N__35506\,
            in2 => \_gnd_net_\,
            in3 => \N__31463\,
            lcout => \b2v_inst11.count_off_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_12\,
            carryout => \b2v_inst11.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_13_c_RNI6BS63_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35302\,
            in1 => \N__35482\,
            in2 => \_gnd_net_\,
            in3 => \N__31460\,
            lcout => \b2v_inst11.count_off_1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_13\,
            carryout => \b2v_inst11.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DT63_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35300\,
            in1 => \N__35524\,
            in2 => \_gnd_net_\,
            in3 => \N__31457\,
            lcout => \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DTZ0Z63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_14_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31453\,
            lcout => \b2v_inst11.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36618\,
            ce => \N__35941\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIGG7EB_15_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31568\,
            in1 => \N__31559\,
            in2 => \_gnd_net_\,
            in3 => \N__35937\,
            lcout => \b2v_inst11.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_15_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31567\,
            lcout => \b2v_inst11.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36489\,
            ce => \N__35942\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIGR5AB_6_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31541\,
            in1 => \N__31552\,
            in2 => \_gnd_net_\,
            in3 => \N__35934\,
            lcout => \b2v_inst11.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_6_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31553\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36489\,
            ce => \N__35942\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIIU6AB_7_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31523\,
            in1 => \N__31534\,
            in2 => \_gnd_net_\,
            in3 => \N__35935\,
            lcout => \b2v_inst11.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_7_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36489\,
            ce => \N__35942\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIK18AB_8_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31505\,
            in1 => \N__31516\,
            in2 => \_gnd_net_\,
            in3 => \N__35936\,
            lcout => \b2v_inst11.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_8_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31517\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36489\,
            ce => \N__35942\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_3_c_RNIFDAI1_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__31945\,
            in1 => \N__31645\,
            in2 => \N__31496\,
            in3 => \N__32623\,
            lcout => \b2v_inst6.count_rst_10\,
            ltout => \b2v_inst6.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIPN6S3_4_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31627\,
            in2 => \N__31499\,
            in3 => \N__32397\,
            lcout => \b2v_inst6.un2_count_1_axb_4\,
            ltout => \b2v_inst6.un2_count_1_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_4_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__31947\,
            in1 => \N__31646\,
            in2 => \N__31637\,
            in3 => \N__32626\,
            lcout => \b2v_inst6.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36349\,
            ce => \N__32432\,
            sr => \N__32635\
        );

    \b2v_inst6.count_RNIPN6S3_0_4_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__31611\,
            in1 => \N__31634\,
            in2 => \N__32431\,
            in3 => \N__31628\,
            lcout => \b2v_inst6.count_1_i_a3_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_2_c_RNIEB9I1_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__31944\,
            in1 => \N__31591\,
            in2 => \N__31616\,
            in3 => \N__32622\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNINK5S3_3_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31580\,
            in2 => \N__31619\,
            in3 => \N__32396\,
            lcout => \b2v_inst6.countZ0Z_3\,
            ltout => \b2v_inst6.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_3_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__31946\,
            in1 => \N__31592\,
            in2 => \N__31583\,
            in3 => \N__32625\,
            lcout => \b2v_inst6.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36349\,
            ce => \N__32432\,
            sr => \N__32635\
        );

    \b2v_inst6.count_11_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__32624\,
            in1 => \N__31855\,
            in2 => \N__31973\,
            in3 => \N__31948\,
            lcout => \b2v_inst6.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36349\,
            ce => \N__32432\,
            sr => \N__32635\
        );

    \b2v_inst6.count_14_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31796\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36530\,
            ce => \N__32430\,
            sr => \N__32650\
        );

    \b2v_inst6.count_RNILH4S3_2_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31764\,
            in1 => \N__31780\,
            in2 => \_gnd_net_\,
            in3 => \N__32373\,
            lcout => \b2v_inst6.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_2_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31766\,
            lcout => \b2v_inst6.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36530\,
            ce => \N__32430\,
            sr => \N__32650\
        );

    \b2v_inst6.count_RNIR2954_14_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31802\,
            in1 => \N__31795\,
            in2 => \_gnd_net_\,
            in3 => \N__32376\,
            lcout => \b2v_inst6.countZ0Z_14\,
            ltout => \b2v_inst6.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNILH4S3_0_2_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__32377\,
            in1 => \N__31781\,
            in2 => \N__31769\,
            in3 => \N__31765\,
            lcout => \b2v_inst6.count_1_i_a3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNINS654_12_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31723\,
            in1 => \N__31743\,
            in2 => \_gnd_net_\,
            in3 => \N__32374\,
            lcout => \b2v_inst6.un2_count_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_12_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31744\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36530\,
            ce => \N__32430\,
            sr => \N__32650\
        );

    \b2v_inst6.count_RNIPV754_13_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31710\,
            in1 => \N__31697\,
            in2 => \_gnd_net_\,
            in3 => \N__32375\,
            lcout => \b2v_inst6.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_6_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32611\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31676\,
            lcout => \b2v_inst6.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36367\,
            ce => \N__32427\,
            sr => \N__32613\
        );

    \b2v_inst6.count_RNI_0_0_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32711\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32076\,
            lcout => \b2v_inst6.N_394\,
            ltout => \b2v_inst6.N_394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_4_c_RNIGFBI1_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__32609\,
            in1 => \N__31993\,
            in2 => \N__31649\,
            in3 => \N__32013\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIRQ7S3_5_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31979\,
            in2 => \N__32018\,
            in3 => \N__32358\,
            lcout => \b2v_inst6.countZ0Z_5\,
            ltout => \b2v_inst6.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_5_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__32612\,
            in1 => \N__31994\,
            in2 => \N__31982\,
            in3 => \N__31923\,
            lcout => \b2v_inst6.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36367\,
            ce => \N__32427\,
            sr => \N__32613\
        );

    \b2v_inst6.un2_count_1_cry_10_c_RNITVOP1_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31966\,
            in1 => \N__31943\,
            in2 => \N__31856\,
            in3 => \N__32610\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNILP554_11_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32359\,
            in1 => \_gnd_net_\,
            in2 => \N__31877\,
            in3 => \N__31874\,
            lcout => \b2v_inst6.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIM6FE1_0_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__32710\,
            in1 => \N__32077\,
            in2 => \_gnd_net_\,
            in3 => \N__32608\,
            lcout => \b2v_inst6.count_RNIM6FE1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNISCBO3_0_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32699\,
            in1 => \N__31865\,
            in2 => \_gnd_net_\,
            in3 => \N__32331\,
            lcout => \b2v_inst6.countZ0Z_0\,
            ltout => \b2v_inst6.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIM6FE1_1_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32680\,
            in2 => \N__31859\,
            in3 => \N__32582\,
            lcout => \b2v_inst6.count_rst_13\,
            ltout => \b2v_inst6.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNITDBO3_0_1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000100010"
        )
    port map (
            in0 => \N__31854\,
            in1 => \N__32662\,
            in2 => \N__31826\,
            in3 => \N__32330\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_1_i_a3_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIOD8DF_1_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31823\,
            in1 => \N__31814\,
            in2 => \N__31805\,
            in3 => \N__32264\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_1_i_a3_12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI9EPHV_2_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32735\,
            in1 => \N__32729\,
            in2 => \N__32720\,
            in3 => \N__32717\,
            lcout => \b2v_inst6.N_389\,
            ltout => \b2v_inst6.N_389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_0_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32078\,
            in2 => \N__32702\,
            in3 => \N__32583\,
            lcout => \b2v_inst6.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36480\,
            ce => \N__32423\,
            sr => \N__32641\
        );

    \b2v_inst6.count_RNITDBO3_1_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32663\,
            in1 => \N__32693\,
            in2 => \_gnd_net_\,
            in3 => \N__32332\,
            lcout => \b2v_inst6.un2_count_1_axb_1\,
            ltout => \b2v_inst6.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_1_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32100\,
            in2 => \N__32666\,
            in3 => \N__32584\,
            lcout => \b2v_inst6.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36480\,
            ce => \N__32423\,
            sr => \N__32641\
        );

    \b2v_inst6.count_RNI37CS3_0_9_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__32474\,
            in1 => \N__32468\,
            in2 => \N__32456\,
            in3 => \N__32372\,
            lcout => \b2v_inst6.count_1_i_a3_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_1_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32255\,
            lcout => \b2v_inst5.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36598\,
            ce => \N__32178\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_0_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32101\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.N_3036_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst31.un6_output_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34928\,
            in1 => \N__33011\,
            in2 => \N__33005\,
            in3 => \N__32972\,
            lcout => vccinaux_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33730\,
            in1 => \N__33312\,
            in2 => \_gnd_net_\,
            in3 => \N__32927\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI7FEU3_0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33920\,
            in1 => \N__32750\,
            in2 => \N__32918\,
            in3 => \N__34062\,
            lcout => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_rn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GPIO_FPGA_SoC_4_RNI8H551_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__34388\,
            in1 => \N__32915\,
            in2 => \_gnd_net_\,
            in3 => \N__34604\,
            lcout => \G_6_i_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_2_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001111"
        )
    port map (
            in0 => \N__33150\,
            in1 => \N__32762\,
            in2 => \N__33731\,
            in3 => \N__34063\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_172_m1_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQK9K2_2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011100000"
        )
    port map (
            in0 => \N__32761\,
            in1 => \N__33500\,
            in2 => \N__32753\,
            in3 => \N__33921\,
            lcout => \b2v_inst11.un1_dutycycle_172_m1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_5_1_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__33378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33313\,
            lcout => \b2v_inst11.N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.g0_0_0_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34395\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34603\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_0_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI0GIO3_6_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__34813\,
            in1 => \N__32744\,
            in2 => \N__32738\,
            in3 => \N__34284\,
            lcout => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQK9K2_3_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000101110"
        )
    port map (
            in0 => \N__34065\,
            in1 => \N__33206\,
            in2 => \N__33514\,
            in3 => \N__33918\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQK9K2_0_5_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__33205\,
            in1 => \N__33146\,
            in2 => \N__33533\,
            in3 => \N__35200\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_4690_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIK9J85_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__33527\,
            in1 => \N__33437\,
            in2 => \N__33530\,
            in3 => \N__33019\,
            lcout => \b2v_inst11.N_6063_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_7_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33380\,
            in2 => \_gnd_net_\,
            in3 => \N__33307\,
            lcout => \b2v_inst11.N_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQK9K2_5_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__33521\,
            in1 => \N__33674\,
            in2 => \N__35204\,
            in3 => \N__33508\,
            lcout => \b2v_inst11.un1_dutycycle_172_m0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111110"
        )
    port map (
            in0 => \N__33431\,
            in1 => \N__33379\,
            in2 => \N__33023\,
            in3 => \N__33306\,
            lcout => \b2v_inst11.N_3099_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010011001"
        )
    port map (
            in0 => \N__35089\,
            in1 => \N__33170\,
            in2 => \_gnd_net_\,
            in3 => \N__34056\,
            lcout => \b2v_inst11.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_3_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35090\,
            in1 => \N__33086\,
            in2 => \N__33080\,
            in3 => \N__34058\,
            lcout => \b2v_inst11.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_5_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010001"
        )
    port map (
            in0 => \N__34057\,
            in1 => \N__35199\,
            in2 => \_gnd_net_\,
            in3 => \N__35088\,
            lcout => OPEN,
            ltout => \N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GPIO_FPGA_SoC_4_RNI498D2_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__34961\,
            in1 => \N__34249\,
            in2 => \N__34949\,
            in3 => \N__34930\,
            lcout => OPEN,
            ltout => \b2v_inst11_un1_clk_100khz_52_and_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINTLA9_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__34826\,
            in1 => \N__34078\,
            in2 => \N__34817\,
            in3 => \N__34795\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIBNRBI_5_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34661\,
            in1 => \_gnd_net_\,
            in2 => \N__34652\,
            in3 => \N__34649\,
            lcout => \b2v_inst11.dutycycle_eena_14_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_4_i_a2_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__34555\,
            in1 => \N__34396\,
            in2 => \_gnd_net_\,
            in3 => \N__34248\,
            lcout => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__34067\,
            in1 => \N__33919\,
            in2 => \_gnd_net_\,
            in3 => \N__33726\,
            lcout => \b2v_inst11.g0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33665\,
            in2 => \_gnd_net_\,
            in3 => \N__33639\,
            lcout => \b2v_inst16.N_208_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI9CS7B_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35339\,
            in1 => \N__33539\,
            in2 => \_gnd_net_\,
            in3 => \N__35930\,
            lcout => \b2v_inst11.count_offZ0Z_1\,
            ltout => \b2v_inst11.count_offZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__35672\,
            in1 => \N__35654\,
            in2 => \N__35630\,
            in3 => \N__35627\,
            lcout => OPEN,
            ltout => \b2v_inst11.un34_clk_100khz_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_0_1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35468\,
            in1 => \N__35369\,
            in2 => \N__35603\,
            in3 => \N__35819\,
            lcout => \b2v_inst11.count_off_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_15_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35528\,
            in1 => \N__35513\,
            in2 => \N__35489\,
            in3 => \N__35332\,
            lcout => \b2v_inst11.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_3_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35462\,
            in1 => \N__35441\,
            in2 => \N__35420\,
            in3 => \N__35393\,
            lcout => \b2v_inst11.un34_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_1_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__35295\,
            in1 => \_gnd_net_\,
            in2 => \N__35333\,
            in3 => \N__35358\,
            lcout => \b2v_inst11.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36579\,
            ce => \N__35939\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35328\,
            in2 => \_gnd_net_\,
            in3 => \N__35296\,
            lcout => \b2v_inst11.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36579\,
            ce => \N__35939\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_9_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35219\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36603\,
            ce => \N__35940\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIM49AB_9_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35225\,
            in1 => \N__35218\,
            in2 => \_gnd_net_\,
            in3 => \N__35896\,
            lcout => \b2v_inst11.count_offZ0Z_9\,
            ltout => \b2v_inst11.count_offZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_9_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35783\,
            in1 => \N__35812\,
            in2 => \N__35822\,
            in3 => \N__35755\,
            lcout => \b2v_inst11.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIVLRAB_10_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35789\,
            in1 => \N__35797\,
            in2 => \_gnd_net_\,
            in3 => \N__35897\,
            lcout => \b2v_inst11.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_10_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36603\,
            ce => \N__35940\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI843EB_11_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35762\,
            in1 => \N__35770\,
            in2 => \_gnd_net_\,
            in3 => \N__35898\,
            lcout => \b2v_inst11.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_11_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36603\,
            ce => \N__35940\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIA74EB_12_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35744\,
            in1 => \N__35732\,
            in2 => \_gnd_net_\,
            in3 => \N__35895\,
            lcout => \b2v_inst11.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_12_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35743\,
            lcout => \b2v_inst11.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36665\,
            ce => \N__35938\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_13_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35725\,
            lcout => \b2v_inst11.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36665\,
            ce => \N__35938\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_2_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35695\,
            lcout => \b2v_inst11.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36665\,
            ce => \N__35938\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36665\,
            ce => \N__35938\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_4_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36715\,
            lcout => \b2v_inst11.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36665\,
            ce => \N__35938\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36688\,
            lcout => \b2v_inst11.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36665\,
            ce => \N__35938\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
