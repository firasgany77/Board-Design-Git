// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 24 2022 21:31:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    input SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    input VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    input VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__37287;
    wire N__37286;
    wire N__37285;
    wire N__37278;
    wire N__37277;
    wire N__37276;
    wire N__37269;
    wire N__37268;
    wire N__37267;
    wire N__37260;
    wire N__37259;
    wire N__37258;
    wire N__37251;
    wire N__37250;
    wire N__37249;
    wire N__37242;
    wire N__37241;
    wire N__37240;
    wire N__37233;
    wire N__37232;
    wire N__37231;
    wire N__37224;
    wire N__37223;
    wire N__37222;
    wire N__37215;
    wire N__37214;
    wire N__37213;
    wire N__37206;
    wire N__37205;
    wire N__37204;
    wire N__37197;
    wire N__37196;
    wire N__37195;
    wire N__37188;
    wire N__37187;
    wire N__37186;
    wire N__37179;
    wire N__37178;
    wire N__37177;
    wire N__37170;
    wire N__37169;
    wire N__37168;
    wire N__37161;
    wire N__37160;
    wire N__37159;
    wire N__37152;
    wire N__37151;
    wire N__37150;
    wire N__37143;
    wire N__37142;
    wire N__37141;
    wire N__37134;
    wire N__37133;
    wire N__37132;
    wire N__37125;
    wire N__37124;
    wire N__37123;
    wire N__37116;
    wire N__37115;
    wire N__37114;
    wire N__37107;
    wire N__37106;
    wire N__37105;
    wire N__37098;
    wire N__37097;
    wire N__37096;
    wire N__37089;
    wire N__37088;
    wire N__37087;
    wire N__37080;
    wire N__37079;
    wire N__37078;
    wire N__37071;
    wire N__37070;
    wire N__37069;
    wire N__37062;
    wire N__37061;
    wire N__37060;
    wire N__37053;
    wire N__37052;
    wire N__37051;
    wire N__37044;
    wire N__37043;
    wire N__37042;
    wire N__37035;
    wire N__37034;
    wire N__37033;
    wire N__37026;
    wire N__37025;
    wire N__37024;
    wire N__37017;
    wire N__37016;
    wire N__37015;
    wire N__37008;
    wire N__37007;
    wire N__37006;
    wire N__36999;
    wire N__36998;
    wire N__36997;
    wire N__36990;
    wire N__36989;
    wire N__36988;
    wire N__36981;
    wire N__36980;
    wire N__36979;
    wire N__36972;
    wire N__36971;
    wire N__36970;
    wire N__36963;
    wire N__36962;
    wire N__36961;
    wire N__36954;
    wire N__36953;
    wire N__36952;
    wire N__36945;
    wire N__36944;
    wire N__36943;
    wire N__36936;
    wire N__36935;
    wire N__36934;
    wire N__36927;
    wire N__36926;
    wire N__36925;
    wire N__36918;
    wire N__36917;
    wire N__36916;
    wire N__36909;
    wire N__36908;
    wire N__36907;
    wire N__36900;
    wire N__36899;
    wire N__36898;
    wire N__36891;
    wire N__36890;
    wire N__36889;
    wire N__36882;
    wire N__36881;
    wire N__36880;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36864;
    wire N__36863;
    wire N__36862;
    wire N__36855;
    wire N__36854;
    wire N__36853;
    wire N__36846;
    wire N__36845;
    wire N__36844;
    wire N__36837;
    wire N__36836;
    wire N__36835;
    wire N__36828;
    wire N__36827;
    wire N__36826;
    wire N__36819;
    wire N__36818;
    wire N__36817;
    wire N__36810;
    wire N__36809;
    wire N__36808;
    wire N__36801;
    wire N__36800;
    wire N__36799;
    wire N__36792;
    wire N__36791;
    wire N__36790;
    wire N__36783;
    wire N__36782;
    wire N__36781;
    wire N__36774;
    wire N__36773;
    wire N__36772;
    wire N__36765;
    wire N__36764;
    wire N__36763;
    wire N__36746;
    wire N__36743;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36661;
    wire N__36658;
    wire N__36657;
    wire N__36656;
    wire N__36653;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36643;
    wire N__36640;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36628;
    wire N__36623;
    wire N__36620;
    wire N__36619;
    wire N__36618;
    wire N__36615;
    wire N__36608;
    wire N__36605;
    wire N__36604;
    wire N__36603;
    wire N__36602;
    wire N__36599;
    wire N__36598;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36586;
    wire N__36583;
    wire N__36582;
    wire N__36581;
    wire N__36580;
    wire N__36579;
    wire N__36576;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36568;
    wire N__36565;
    wire N__36560;
    wire N__36557;
    wire N__36556;
    wire N__36553;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36542;
    wire N__36541;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36531;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36514;
    wire N__36511;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36503;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36491;
    wire N__36490;
    wire N__36489;
    wire N__36486;
    wire N__36485;
    wire N__36482;
    wire N__36481;
    wire N__36480;
    wire N__36479;
    wire N__36474;
    wire N__36471;
    wire N__36470;
    wire N__36469;
    wire N__36468;
    wire N__36465;
    wire N__36454;
    wire N__36451;
    wire N__36450;
    wire N__36449;
    wire N__36448;
    wire N__36447;
    wire N__36442;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36436;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36422;
    wire N__36421;
    wire N__36420;
    wire N__36417;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36403;
    wire N__36402;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36394;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36372;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36360;
    wire N__36357;
    wire N__36356;
    wire N__36351;
    wire N__36350;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36339;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36315;
    wire N__36314;
    wire N__36309;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36267;
    wire N__36264;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36213;
    wire N__36210;
    wire N__36209;
    wire N__36208;
    wire N__36207;
    wire N__36202;
    wire N__36199;
    wire N__36198;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36173;
    wire N__36168;
    wire N__36167;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36139;
    wire N__36136;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36103;
    wire N__36100;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36054;
    wire N__36047;
    wire N__36040;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36011;
    wire N__36002;
    wire N__36001;
    wire N__35994;
    wire N__35989;
    wire N__35986;
    wire N__35979;
    wire N__35974;
    wire N__35971;
    wire N__35962;
    wire N__35959;
    wire N__35942;
    wire N__35941;
    wire N__35940;
    wire N__35939;
    wire N__35938;
    wire N__35937;
    wire N__35936;
    wire N__35935;
    wire N__35934;
    wire N__35931;
    wire N__35930;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35896;
    wire N__35895;
    wire N__35892;
    wire N__35891;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35875;
    wire N__35868;
    wire N__35859;
    wire N__35856;
    wire N__35843;
    wire N__35834;
    wire N__35831;
    wire N__35822;
    wire N__35819;
    wire N__35816;
    wire N__35813;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35798;
    wire N__35797;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35771;
    wire N__35770;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35756;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35744;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35654;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35630;
    wire N__35627;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35603;
    wire N__35600;
    wire N__35599;
    wire N__35596;
    wire N__35595;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35585;
    wire N__35584;
    wire N__35583;
    wire N__35578;
    wire N__35577;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35542;
    wire N__35537;
    wire N__35528;
    wire N__35525;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35441;
    wire N__35438;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35420;
    wire N__35417;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35393;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35362;
    wire N__35359;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35344;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35332;
    wire N__35329;
    wire N__35328;
    wire N__35327;
    wire N__35326;
    wire N__35325;
    wire N__35318;
    wire N__35315;
    wire N__35310;
    wire N__35303;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35299;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35295;
    wire N__35288;
    wire N__35279;
    wire N__35278;
    wire N__35277;
    wire N__35276;
    wire N__35275;
    wire N__35274;
    wire N__35273;
    wire N__35272;
    wire N__35271;
    wire N__35266;
    wire N__35261;
    wire N__35254;
    wire N__35245;
    wire N__35242;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35219;
    wire N__35218;
    wire N__35213;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35200;
    wire N__35199;
    wire N__35198;
    wire N__35193;
    wire N__35192;
    wire N__35189;
    wire N__35188;
    wire N__35185;
    wire N__35184;
    wire N__35183;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35175;
    wire N__35172;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35139;
    wire N__35136;
    wire N__35135;
    wire N__35128;
    wire N__35121;
    wire N__35118;
    wire N__35111;
    wire N__35110;
    wire N__35109;
    wire N__35108;
    wire N__35107;
    wire N__35106;
    wire N__35105;
    wire N__35104;
    wire N__35097;
    wire N__35096;
    wire N__35095;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35091;
    wire N__35090;
    wire N__35089;
    wire N__35088;
    wire N__35085;
    wire N__35084;
    wire N__35083;
    wire N__35078;
    wire N__35073;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35062;
    wire N__35059;
    wire N__35052;
    wire N__35045;
    wire N__35040;
    wire N__35037;
    wire N__35032;
    wire N__35031;
    wire N__35030;
    wire N__35027;
    wire N__35026;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35014;
    wire N__35007;
    wire N__35004;
    wire N__34999;
    wire N__34996;
    wire N__34991;
    wire N__34986;
    wire N__34983;
    wire N__34976;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34938;
    wire N__34933;
    wire N__34932;
    wire N__34931;
    wire N__34930;
    wire N__34929;
    wire N__34928;
    wire N__34927;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34884;
    wire N__34883;
    wire N__34878;
    wire N__34875;
    wire N__34870;
    wire N__34865;
    wire N__34862;
    wire N__34857;
    wire N__34854;
    wire N__34849;
    wire N__34846;
    wire N__34837;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34811;
    wire N__34810;
    wire N__34809;
    wire N__34808;
    wire N__34807;
    wire N__34806;
    wire N__34805;
    wire N__34804;
    wire N__34801;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34792;
    wire N__34787;
    wire N__34784;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34757;
    wire N__34752;
    wire N__34749;
    wire N__34748;
    wire N__34747;
    wire N__34744;
    wire N__34743;
    wire N__34740;
    wire N__34739;
    wire N__34738;
    wire N__34737;
    wire N__34732;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34699;
    wire N__34694;
    wire N__34691;
    wire N__34686;
    wire N__34683;
    wire N__34678;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34642;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34624;
    wire N__34623;
    wire N__34622;
    wire N__34621;
    wire N__34620;
    wire N__34619;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34604;
    wire N__34603;
    wire N__34602;
    wire N__34601;
    wire N__34600;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34556;
    wire N__34555;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34539;
    wire N__34536;
    wire N__34531;
    wire N__34526;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34508;
    wire N__34503;
    wire N__34496;
    wire N__34495;
    wire N__34494;
    wire N__34493;
    wire N__34488;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34469;
    wire N__34462;
    wire N__34457;
    wire N__34456;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34434;
    wire N__34433;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34422;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34405;
    wire N__34400;
    wire N__34397;
    wire N__34396;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34355;
    wire N__34352;
    wire N__34343;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34312;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34301;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34290;
    wire N__34289;
    wire N__34288;
    wire N__34287;
    wire N__34286;
    wire N__34285;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34277;
    wire N__34270;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34252;
    wire N__34251;
    wire N__34250;
    wire N__34249;
    wire N__34248;
    wire N__34245;
    wire N__34242;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34230;
    wire N__34225;
    wire N__34222;
    wire N__34221;
    wire N__34220;
    wire N__34219;
    wire N__34216;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34201;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34186;
    wire N__34183;
    wire N__34182;
    wire N__34181;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34117;
    wire N__34110;
    wire N__34107;
    wire N__34102;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34067;
    wire N__34066;
    wire N__34065;
    wire N__34064;
    wire N__34063;
    wire N__34062;
    wire N__34061;
    wire N__34060;
    wire N__34059;
    wire N__34058;
    wire N__34057;
    wire N__34056;
    wire N__34053;
    wire N__34052;
    wire N__34049;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34041;
    wire N__34040;
    wire N__34035;
    wire N__34032;
    wire N__34027;
    wire N__34020;
    wire N__34017;
    wire N__34016;
    wire N__34015;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34000;
    wire N__33995;
    wire N__33990;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33938;
    wire N__33937;
    wire N__33934;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33921;
    wire N__33920;
    wire N__33919;
    wire N__33918;
    wire N__33917;
    wire N__33914;
    wire N__33909;
    wire N__33904;
    wire N__33899;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33891;
    wire N__33888;
    wire N__33887;
    wire N__33886;
    wire N__33885;
    wire N__33884;
    wire N__33883;
    wire N__33882;
    wire N__33881;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33867;
    wire N__33866;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33854;
    wire N__33851;
    wire N__33850;
    wire N__33849;
    wire N__33848;
    wire N__33847;
    wire N__33846;
    wire N__33845;
    wire N__33844;
    wire N__33843;
    wire N__33842;
    wire N__33837;
    wire N__33832;
    wire N__33827;
    wire N__33824;
    wire N__33819;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33796;
    wire N__33793;
    wire N__33786;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33764;
    wire N__33759;
    wire N__33754;
    wire N__33745;
    wire N__33740;
    wire N__33731;
    wire N__33730;
    wire N__33727;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33716;
    wire N__33711;
    wire N__33708;
    wire N__33707;
    wire N__33704;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33639;
    wire N__33634;
    wire N__33633;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33622;
    wire N__33619;
    wire N__33618;
    wire N__33617;
    wire N__33614;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33583;
    wire N__33578;
    wire N__33577;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33514;
    wire N__33513;
    wire N__33510;
    wire N__33509;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33501;
    wire N__33500;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33451;
    wire N__33448;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33418;
    wire N__33417;
    wire N__33416;
    wire N__33415;
    wire N__33412;
    wire N__33411;
    wire N__33408;
    wire N__33407;
    wire N__33406;
    wire N__33403;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33385;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33378;
    wire N__33377;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33361;
    wire N__33356;
    wire N__33353;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33330;
    wire N__33327;
    wire N__33314;
    wire N__33313;
    wire N__33312;
    wire N__33311;
    wire N__33308;
    wire N__33307;
    wire N__33306;
    wire N__33305;
    wire N__33304;
    wire N__33299;
    wire N__33294;
    wire N__33293;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33281;
    wire N__33280;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33258;
    wire N__33253;
    wire N__33250;
    wire N__33243;
    wire N__33240;
    wire N__33235;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33206;
    wire N__33205;
    wire N__33200;
    wire N__33197;
    wire N__33196;
    wire N__33193;
    wire N__33192;
    wire N__33191;
    wire N__33188;
    wire N__33187;
    wire N__33186;
    wire N__33183;
    wire N__33178;
    wire N__33175;
    wire N__33174;
    wire N__33171;
    wire N__33170;
    wire N__33167;
    wire N__33166;
    wire N__33165;
    wire N__33162;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33150;
    wire N__33147;
    wire N__33146;
    wire N__33141;
    wire N__33138;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33114;
    wire N__33111;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33079;
    wire N__33078;
    wire N__33075;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33050;
    wire N__33049;
    wire N__33046;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33028;
    wire N__33023;
    wire N__33020;
    wire N__33019;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32989;
    wire N__32988;
    wire N__32987;
    wire N__32986;
    wire N__32983;
    wire N__32976;
    wire N__32973;
    wire N__32972;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32911;
    wire N__32910;
    wire N__32909;
    wire N__32908;
    wire N__32907;
    wire N__32906;
    wire N__32905;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32881;
    wire N__32876;
    wire N__32875;
    wire N__32874;
    wire N__32873;
    wire N__32870;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32847;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32828;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32813;
    wire N__32808;
    wire N__32803;
    wire N__32800;
    wire N__32797;
    wire N__32792;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32770;
    wire N__32765;
    wire N__32762;
    wire N__32761;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32710;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32671;
    wire N__32666;
    wire N__32663;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32641;
    wire N__32636;
    wire N__32635;
    wire N__32630;
    wire N__32627;
    wire N__32626;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32622;
    wire N__32621;
    wire N__32620;
    wire N__32619;
    wire N__32618;
    wire N__32617;
    wire N__32616;
    wire N__32615;
    wire N__32614;
    wire N__32613;
    wire N__32612;
    wire N__32611;
    wire N__32610;
    wire N__32609;
    wire N__32608;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32596;
    wire N__32585;
    wire N__32584;
    wire N__32583;
    wire N__32582;
    wire N__32577;
    wire N__32570;
    wire N__32567;
    wire N__32562;
    wire N__32549;
    wire N__32548;
    wire N__32547;
    wire N__32544;
    wire N__32543;
    wire N__32542;
    wire N__32541;
    wire N__32536;
    wire N__32531;
    wire N__32524;
    wire N__32517;
    wire N__32512;
    wire N__32507;
    wire N__32504;
    wire N__32497;
    wire N__32490;
    wire N__32483;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32456;
    wire N__32455;
    wire N__32452;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32432;
    wire N__32431;
    wire N__32430;
    wire N__32429;
    wire N__32428;
    wire N__32427;
    wire N__32424;
    wire N__32423;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32397;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32383;
    wire N__32378;
    wire N__32377;
    wire N__32376;
    wire N__32375;
    wire N__32374;
    wire N__32373;
    wire N__32372;
    wire N__32369;
    wire N__32368;
    wire N__32367;
    wire N__32366;
    wire N__32365;
    wire N__32364;
    wire N__32363;
    wire N__32362;
    wire N__32361;
    wire N__32360;
    wire N__32359;
    wire N__32358;
    wire N__32353;
    wire N__32344;
    wire N__32333;
    wire N__32332;
    wire N__32331;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32317;
    wire N__32312;
    wire N__32303;
    wire N__32298;
    wire N__32295;
    wire N__32290;
    wire N__32283;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32224;
    wire N__32223;
    wire N__32222;
    wire N__32221;
    wire N__32220;
    wire N__32219;
    wire N__32216;
    wire N__32215;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32184;
    wire N__32183;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32175;
    wire N__32174;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32101;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32078;
    wire N__32077;
    wire N__32076;
    wire N__32073;
    wire N__32068;
    wire N__32063;
    wire N__32060;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32052;
    wire N__32049;
    wire N__32048;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32029;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32014;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31994;
    wire N__31993;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31955;
    wire N__31954;
    wire N__31953;
    wire N__31952;
    wire N__31951;
    wire N__31950;
    wire N__31949;
    wire N__31948;
    wire N__31947;
    wire N__31946;
    wire N__31945;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31936;
    wire N__31931;
    wire N__31924;
    wire N__31923;
    wire N__31912;
    wire N__31909;
    wire N__31904;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31884;
    wire N__31877;
    wire N__31874;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31855;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31835;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31795;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31781;
    wire N__31780;
    wire N__31777;
    wire N__31774;
    wire N__31769;
    wire N__31766;
    wire N__31765;
    wire N__31764;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31745;
    wire N__31744;
    wire N__31743;
    wire N__31740;
    wire N__31735;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31712;
    wire N__31711;
    wire N__31710;
    wire N__31705;
    wire N__31702;
    wire N__31697;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31645;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31627;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31615;
    wire N__31612;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31592;
    wire N__31591;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31567;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31552;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31534;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31516;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31387;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31377;
    wire N__31376;
    wire N__31375;
    wire N__31374;
    wire N__31373;
    wire N__31370;
    wire N__31369;
    wire N__31366;
    wire N__31365;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31351;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31332;
    wire N__31327;
    wire N__31324;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31312;
    wire N__31311;
    wire N__31310;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31298;
    wire N__31291;
    wire N__31288;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31272;
    wire N__31267;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31249;
    wire N__31248;
    wire N__31245;
    wire N__31244;
    wire N__31241;
    wire N__31240;
    wire N__31239;
    wire N__31238;
    wire N__31237;
    wire N__31236;
    wire N__31235;
    wire N__31232;
    wire N__31229;
    wire N__31228;
    wire N__31227;
    wire N__31226;
    wire N__31225;
    wire N__31222;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31211;
    wire N__31210;
    wire N__31209;
    wire N__31200;
    wire N__31197;
    wire N__31196;
    wire N__31195;
    wire N__31194;
    wire N__31193;
    wire N__31192;
    wire N__31191;
    wire N__31190;
    wire N__31189;
    wire N__31186;
    wire N__31177;
    wire N__31172;
    wire N__31165;
    wire N__31162;
    wire N__31157;
    wire N__31154;
    wire N__31153;
    wire N__31152;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31140;
    wire N__31135;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31119;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31101;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31070;
    wire N__31061;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31051;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31039;
    wire N__31038;
    wire N__31037;
    wire N__31036;
    wire N__31033;
    wire N__31032;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31021;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30985;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30952;
    wire N__30947;
    wire N__30944;
    wire N__30939;
    wire N__30936;
    wire N__30931;
    wire N__30928;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30898;
    wire N__30897;
    wire N__30896;
    wire N__30895;
    wire N__30894;
    wire N__30893;
    wire N__30890;
    wire N__30885;
    wire N__30884;
    wire N__30883;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30871;
    wire N__30866;
    wire N__30859;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30827;
    wire N__30826;
    wire N__30821;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30811;
    wire N__30808;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30778;
    wire N__30777;
    wire N__30774;
    wire N__30769;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30734;
    wire N__30733;
    wire N__30732;
    wire N__30731;
    wire N__30730;
    wire N__30729;
    wire N__30728;
    wire N__30727;
    wire N__30726;
    wire N__30725;
    wire N__30724;
    wire N__30719;
    wire N__30714;
    wire N__30707;
    wire N__30706;
    wire N__30705;
    wire N__30702;
    wire N__30701;
    wire N__30700;
    wire N__30699;
    wire N__30698;
    wire N__30695;
    wire N__30694;
    wire N__30693;
    wire N__30692;
    wire N__30691;
    wire N__30690;
    wire N__30689;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30681;
    wire N__30680;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30653;
    wire N__30644;
    wire N__30639;
    wire N__30638;
    wire N__30637;
    wire N__30636;
    wire N__30635;
    wire N__30634;
    wire N__30633;
    wire N__30632;
    wire N__30631;
    wire N__30628;
    wire N__30627;
    wire N__30624;
    wire N__30623;
    wire N__30614;
    wire N__30613;
    wire N__30612;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30604;
    wire N__30603;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30597;
    wire N__30596;
    wire N__30595;
    wire N__30592;
    wire N__30583;
    wire N__30580;
    wire N__30579;
    wire N__30578;
    wire N__30577;
    wire N__30576;
    wire N__30575;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30563;
    wire N__30560;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30552;
    wire N__30549;
    wire N__30544;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30527;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30515;
    wire N__30514;
    wire N__30511;
    wire N__30510;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30496;
    wire N__30489;
    wire N__30482;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30464;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30429;
    wire N__30424;
    wire N__30421;
    wire N__30420;
    wire N__30415;
    wire N__30410;
    wire N__30407;
    wire N__30402;
    wire N__30399;
    wire N__30392;
    wire N__30391;
    wire N__30388;
    wire N__30379;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30361;
    wire N__30358;
    wire N__30351;
    wire N__30348;
    wire N__30337;
    wire N__30326;
    wire N__30325;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30310;
    wire N__30309;
    wire N__30308;
    wire N__30307;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30290;
    wire N__30287;
    wire N__30286;
    wire N__30283;
    wire N__30278;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30272;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30251;
    wire N__30248;
    wire N__30241;
    wire N__30230;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30196;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30184;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30176;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30168;
    wire N__30167;
    wire N__30166;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30144;
    wire N__30143;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30126;
    wire N__30119;
    wire N__30116;
    wire N__30115;
    wire N__30112;
    wire N__30107;
    wire N__30102;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30078;
    wire N__30073;
    wire N__30068;
    wire N__30059;
    wire N__30056;
    wire N__30055;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30019;
    wire N__30016;
    wire N__30011;
    wire N__30008;
    wire N__30007;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29995;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29980;
    wire N__29975;
    wire N__29972;
    wire N__29971;
    wire N__29970;
    wire N__29969;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29963;
    wire N__29962;
    wire N__29961;
    wire N__29958;
    wire N__29957;
    wire N__29954;
    wire N__29953;
    wire N__29948;
    wire N__29943;
    wire N__29942;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29927;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29912;
    wire N__29907;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29892;
    wire N__29891;
    wire N__29890;
    wire N__29887;
    wire N__29886;
    wire N__29883;
    wire N__29878;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29826;
    wire N__29813;
    wire N__29810;
    wire N__29809;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29755;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29743;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29714;
    wire N__29713;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29681;
    wire N__29680;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29638;
    wire N__29637;
    wire N__29636;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29624;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29609;
    wire N__29608;
    wire N__29607;
    wire N__29602;
    wire N__29597;
    wire N__29592;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29536;
    wire N__29535;
    wire N__29530;
    wire N__29527;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29515;
    wire N__29514;
    wire N__29511;
    wire N__29506;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29491;
    wire N__29490;
    wire N__29489;
    wire N__29488;
    wire N__29487;
    wire N__29484;
    wire N__29477;
    wire N__29472;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29451;
    wire N__29444;
    wire N__29441;
    wire N__29440;
    wire N__29437;
    wire N__29436;
    wire N__29429;
    wire N__29426;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29408;
    wire N__29407;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29389;
    wire N__29386;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29334;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29301;
    wire N__29294;
    wire N__29293;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29285;
    wire N__29284;
    wire N__29283;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29264;
    wire N__29261;
    wire N__29252;
    wire N__29249;
    wire N__29248;
    wire N__29247;
    wire N__29246;
    wire N__29245;
    wire N__29244;
    wire N__29243;
    wire N__29242;
    wire N__29239;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29206;
    wire N__29203;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29168;
    wire N__29167;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29149;
    wire N__29148;
    wire N__29147;
    wire N__29146;
    wire N__29145;
    wire N__29142;
    wire N__29141;
    wire N__29136;
    wire N__29135;
    wire N__29134;
    wire N__29133;
    wire N__29132;
    wire N__29127;
    wire N__29126;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29120;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29111;
    wire N__29110;
    wire N__29109;
    wire N__29108;
    wire N__29107;
    wire N__29106;
    wire N__29103;
    wire N__29098;
    wire N__29097;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29093;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29070;
    wire N__29063;
    wire N__29060;
    wire N__29053;
    wire N__29048;
    wire N__29043;
    wire N__29032;
    wire N__29029;
    wire N__29024;
    wire N__29021;
    wire N__29016;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28994;
    wire N__28991;
    wire N__28982;
    wire N__28981;
    wire N__28980;
    wire N__28977;
    wire N__28976;
    wire N__28975;
    wire N__28974;
    wire N__28973;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28965;
    wire N__28964;
    wire N__28963;
    wire N__28962;
    wire N__28961;
    wire N__28960;
    wire N__28959;
    wire N__28956;
    wire N__28951;
    wire N__28946;
    wire N__28945;
    wire N__28942;
    wire N__28941;
    wire N__28940;
    wire N__28939;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28918;
    wire N__28917;
    wire N__28916;
    wire N__28915;
    wire N__28914;
    wire N__28911;
    wire N__28904;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28883;
    wire N__28878;
    wire N__28871;
    wire N__28866;
    wire N__28863;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28845;
    wire N__28834;
    wire N__28827;
    wire N__28808;
    wire N__28807;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28795;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28780;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28699;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28667;
    wire N__28664;
    wire N__28663;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28642;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28597;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28572;
    wire N__28571;
    wire N__28570;
    wire N__28569;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28558;
    wire N__28557;
    wire N__28556;
    wire N__28555;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28543;
    wire N__28542;
    wire N__28541;
    wire N__28540;
    wire N__28539;
    wire N__28538;
    wire N__28531;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28501;
    wire N__28498;
    wire N__28493;
    wire N__28490;
    wire N__28489;
    wire N__28488;
    wire N__28487;
    wire N__28486;
    wire N__28485;
    wire N__28480;
    wire N__28475;
    wire N__28468;
    wire N__28465;
    wire N__28456;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28423;
    wire N__28422;
    wire N__28419;
    wire N__28414;
    wire N__28413;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28340;
    wire N__28337;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28286;
    wire N__28285;
    wire N__28284;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28247;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28219;
    wire N__28216;
    wire N__28215;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28177;
    wire N__28174;
    wire N__28173;
    wire N__28170;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28156;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28144;
    wire N__28139;
    wire N__28130;
    wire N__28129;
    wire N__28128;
    wire N__28127;
    wire N__28126;
    wire N__28123;
    wire N__28114;
    wire N__28111;
    wire N__28110;
    wire N__28109;
    wire N__28108;
    wire N__28107;
    wire N__28106;
    wire N__28105;
    wire N__28104;
    wire N__28103;
    wire N__28100;
    wire N__28099;
    wire N__28098;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28090;
    wire N__28089;
    wire N__28080;
    wire N__28073;
    wire N__28070;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28052;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28015;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27975;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27951;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27928;
    wire N__27927;
    wire N__27924;
    wire N__27919;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27872;
    wire N__27869;
    wire N__27868;
    wire N__27863;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27823;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27808;
    wire N__27807;
    wire N__27804;
    wire N__27803;
    wire N__27798;
    wire N__27793;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27740;
    wire N__27737;
    wire N__27736;
    wire N__27735;
    wire N__27734;
    wire N__27731;
    wire N__27726;
    wire N__27723;
    wire N__27722;
    wire N__27721;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27709;
    wire N__27704;
    wire N__27699;
    wire N__27694;
    wire N__27689;
    wire N__27688;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27661;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27646;
    wire N__27645;
    wire N__27644;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27636;
    wire N__27633;
    wire N__27628;
    wire N__27623;
    wire N__27622;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27580;
    wire N__27579;
    wire N__27576;
    wire N__27575;
    wire N__27574;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27532;
    wire N__27529;
    wire N__27528;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27515;
    wire N__27514;
    wire N__27513;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27499;
    wire N__27496;
    wire N__27495;
    wire N__27490;
    wire N__27487;
    wire N__27480;
    wire N__27473;
    wire N__27464;
    wire N__27463;
    wire N__27460;
    wire N__27459;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27437;
    wire N__27434;
    wire N__27433;
    wire N__27432;
    wire N__27429;
    wire N__27424;
    wire N__27421;
    wire N__27414;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27382;
    wire N__27381;
    wire N__27374;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27362;
    wire N__27359;
    wire N__27358;
    wire N__27357;
    wire N__27352;
    wire N__27349;
    wire N__27344;
    wire N__27343;
    wire N__27342;
    wire N__27341;
    wire N__27336;
    wire N__27335;
    wire N__27332;
    wire N__27331;
    wire N__27330;
    wire N__27329;
    wire N__27326;
    wire N__27325;
    wire N__27324;
    wire N__27323;
    wire N__27320;
    wire N__27315;
    wire N__27314;
    wire N__27313;
    wire N__27310;
    wire N__27309;
    wire N__27308;
    wire N__27307;
    wire N__27306;
    wire N__27305;
    wire N__27304;
    wire N__27303;
    wire N__27302;
    wire N__27297;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27289;
    wire N__27284;
    wire N__27279;
    wire N__27274;
    wire N__27271;
    wire N__27262;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27240;
    wire N__27237;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27221;
    wire N__27220;
    wire N__27219;
    wire N__27218;
    wire N__27217;
    wire N__27216;
    wire N__27215;
    wire N__27214;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27185;
    wire N__27174;
    wire N__27169;
    wire N__27166;
    wire N__27143;
    wire N__27142;
    wire N__27141;
    wire N__27140;
    wire N__27139;
    wire N__27136;
    wire N__27135;
    wire N__27132;
    wire N__27131;
    wire N__27130;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27122;
    wire N__27121;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27111;
    wire N__27102;
    wire N__27093;
    wire N__27086;
    wire N__27081;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27046;
    wire N__27045;
    wire N__27044;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27023;
    wire N__27020;
    wire N__27019;
    wire N__27016;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__26999;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26984;
    wire N__26981;
    wire N__26980;
    wire N__26979;
    wire N__26976;
    wire N__26975;
    wire N__26974;
    wire N__26973;
    wire N__26970;
    wire N__26965;
    wire N__26964;
    wire N__26963;
    wire N__26962;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26942;
    wire N__26941;
    wire N__26940;
    wire N__26939;
    wire N__26938;
    wire N__26935;
    wire N__26928;
    wire N__26921;
    wire N__26918;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26865;
    wire N__26864;
    wire N__26863;
    wire N__26858;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26828;
    wire N__26827;
    wire N__26826;
    wire N__26825;
    wire N__26822;
    wire N__26821;
    wire N__26820;
    wire N__26819;
    wire N__26816;
    wire N__26815;
    wire N__26814;
    wire N__26813;
    wire N__26808;
    wire N__26803;
    wire N__26802;
    wire N__26801;
    wire N__26800;
    wire N__26799;
    wire N__26798;
    wire N__26797;
    wire N__26796;
    wire N__26787;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26755;
    wire N__26744;
    wire N__26741;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26707;
    wire N__26706;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26689;
    wire N__26688;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26665;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26633;
    wire N__26632;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26600;
    wire N__26599;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26575;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26519;
    wire N__26516;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26368;
    wire N__26367;
    wire N__26364;
    wire N__26359;
    wire N__26354;
    wire N__26351;
    wire N__26350;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26317;
    wire N__26316;
    wire N__26313;
    wire N__26308;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26296;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26275;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26189;
    wire N__26188;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26173;
    wire N__26172;
    wire N__26171;
    wire N__26170;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26156;
    wire N__26155;
    wire N__26154;
    wire N__26153;
    wire N__26152;
    wire N__26149;
    wire N__26148;
    wire N__26147;
    wire N__26146;
    wire N__26145;
    wire N__26144;
    wire N__26143;
    wire N__26142;
    wire N__26139;
    wire N__26134;
    wire N__26133;
    wire N__26132;
    wire N__26127;
    wire N__26124;
    wire N__26119;
    wire N__26112;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26092;
    wire N__26075;
    wire N__26074;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26059;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25948;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25919;
    wire N__25918;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25897;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25864;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25847;
    wire N__25846;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25831;
    wire N__25830;
    wire N__25827;
    wire N__25822;
    wire N__25817;
    wire N__25814;
    wire N__25813;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25787;
    wire N__25784;
    wire N__25783;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25765;
    wire N__25764;
    wire N__25761;
    wire N__25756;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25721;
    wire N__25718;
    wire N__25717;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25694;
    wire N__25693;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25654;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25637;
    wire N__25634;
    wire N__25633;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25549;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25531;
    wire N__25526;
    wire N__25523;
    wire N__25522;
    wire N__25521;
    wire N__25518;
    wire N__25513;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25496;
    wire N__25493;
    wire N__25492;
    wire N__25487;
    wire N__25484;
    wire N__25483;
    wire N__25480;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25460;
    wire N__25459;
    wire N__25456;
    wire N__25455;
    wire N__25454;
    wire N__25453;
    wire N__25452;
    wire N__25451;
    wire N__25450;
    wire N__25449;
    wire N__25444;
    wire N__25439;
    wire N__25430;
    wire N__25427;
    wire N__25426;
    wire N__25425;
    wire N__25424;
    wire N__25423;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25415;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25403;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25384;
    wire N__25381;
    wire N__25368;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25321;
    wire N__25320;
    wire N__25317;
    wire N__25316;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25302;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25290;
    wire N__25287;
    wire N__25282;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25246;
    wire N__25241;
    wire N__25240;
    wire N__25239;
    wire N__25238;
    wire N__25235;
    wire N__25228;
    wire N__25223;
    wire N__25220;
    wire N__25219;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25215;
    wire N__25212;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25197;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25182;
    wire N__25179;
    wire N__25178;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25161;
    wire N__25156;
    wire N__25153;
    wire N__25142;
    wire N__25141;
    wire N__25140;
    wire N__25139;
    wire N__25138;
    wire N__25135;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25116;
    wire N__25113;
    wire N__25112;
    wire N__25111;
    wire N__25104;
    wire N__25099;
    wire N__25096;
    wire N__25091;
    wire N__25088;
    wire N__25087;
    wire N__25086;
    wire N__25085;
    wire N__25082;
    wire N__25081;
    wire N__25080;
    wire N__25079;
    wire N__25076;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25061;
    wire N__25060;
    wire N__25057;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25043;
    wire N__25038;
    wire N__25037;
    wire N__25036;
    wire N__25035;
    wire N__25030;
    wire N__25027;
    wire N__25020;
    wire N__25017;
    wire N__25012;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24994;
    wire N__24993;
    wire N__24988;
    wire N__24987;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24969;
    wire N__24964;
    wire N__24961;
    wire N__24956;
    wire N__24955;
    wire N__24952;
    wire N__24951;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24943;
    wire N__24940;
    wire N__24939;
    wire N__24936;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24918;
    wire N__24917;
    wire N__24916;
    wire N__24913;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24788;
    wire N__24787;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24743;
    wire N__24740;
    wire N__24739;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24727;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24712;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24704;
    wire N__24703;
    wire N__24700;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24689;
    wire N__24688;
    wire N__24685;
    wire N__24680;
    wire N__24677;
    wire N__24676;
    wire N__24671;
    wire N__24666;
    wire N__24663;
    wire N__24658;
    wire N__24655;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24631;
    wire N__24630;
    wire N__24629;
    wire N__24628;
    wire N__24627;
    wire N__24624;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24609;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24598;
    wire N__24597;
    wire N__24596;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24588;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24572;
    wire N__24569;
    wire N__24568;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24557;
    wire N__24556;
    wire N__24555;
    wire N__24552;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24530;
    wire N__24525;
    wire N__24518;
    wire N__24511;
    wire N__24508;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24461;
    wire N__24460;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24448;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24433;
    wire N__24432;
    wire N__24429;
    wire N__24424;
    wire N__24421;
    wire N__24416;
    wire N__24415;
    wire N__24412;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24352;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24301;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24262;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24228;
    wire N__24223;
    wire N__24220;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24193;
    wire N__24192;
    wire N__24191;
    wire N__24190;
    wire N__24187;
    wire N__24176;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24153;
    wire N__24150;
    wire N__24145;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24124;
    wire N__24121;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24104;
    wire N__24103;
    wire N__24100;
    wire N__24099;
    wire N__24094;
    wire N__24091;
    wire N__24086;
    wire N__24083;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24055;
    wire N__24054;
    wire N__24051;
    wire N__24046;
    wire N__24043;
    wire N__24038;
    wire N__24037;
    wire N__24034;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24002;
    wire N__24001;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23972;
    wire N__23971;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23939;
    wire N__23936;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23924;
    wire N__23923;
    wire N__23920;
    wire N__23917;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23896;
    wire N__23895;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23874;
    wire N__23869;
    wire N__23866;
    wire N__23861;
    wire N__23860;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23828;
    wire N__23827;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23786;
    wire N__23783;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23743;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23722;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23686;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23662;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23605;
    wire N__23602;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23587;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23572;
    wire N__23571;
    wire N__23570;
    wire N__23569;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23563;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23546;
    wire N__23545;
    wire N__23544;
    wire N__23543;
    wire N__23542;
    wire N__23541;
    wire N__23538;
    wire N__23533;
    wire N__23532;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23506;
    wire N__23503;
    wire N__23498;
    wire N__23493;
    wire N__23488;
    wire N__23485;
    wire N__23480;
    wire N__23475;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23449;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23437;
    wire N__23436;
    wire N__23435;
    wire N__23434;
    wire N__23431;
    wire N__23426;
    wire N__23425;
    wire N__23424;
    wire N__23423;
    wire N__23422;
    wire N__23419;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23401;
    wire N__23400;
    wire N__23399;
    wire N__23398;
    wire N__23397;
    wire N__23394;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23355;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23227;
    wire N__23222;
    wire N__23219;
    wire N__23218;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23197;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23155;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23140;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23128;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23110;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23092;
    wire N__23091;
    wire N__23088;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23065;
    wire N__23062;
    wire N__23061;
    wire N__23058;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23040;
    wire N__23037;
    wire N__23032;
    wire N__23021;
    wire N__23018;
    wire N__23017;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22957;
    wire N__22956;
    wire N__22953;
    wire N__22948;
    wire N__22943;
    wire N__22940;
    wire N__22939;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22918;
    wire N__22917;
    wire N__22916;
    wire N__22915;
    wire N__22914;
    wire N__22913;
    wire N__22912;
    wire N__22909;
    wire N__22908;
    wire N__22905;
    wire N__22900;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22878;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22866;
    wire N__22861;
    wire N__22858;
    wire N__22853;
    wire N__22850;
    wire N__22841;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22813;
    wire N__22810;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22795;
    wire N__22792;
    wire N__22791;
    wire N__22790;
    wire N__22789;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22781;
    wire N__22780;
    wire N__22779;
    wire N__22778;
    wire N__22777;
    wire N__22776;
    wire N__22775;
    wire N__22774;
    wire N__22773;
    wire N__22772;
    wire N__22771;
    wire N__22770;
    wire N__22769;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22761;
    wire N__22760;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22742;
    wire N__22735;
    wire N__22732;
    wire N__22723;
    wire N__22716;
    wire N__22707;
    wire N__22702;
    wire N__22685;
    wire N__22684;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22666;
    wire N__22665;
    wire N__22662;
    wire N__22661;
    wire N__22660;
    wire N__22659;
    wire N__22658;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22650;
    wire N__22647;
    wire N__22646;
    wire N__22643;
    wire N__22642;
    wire N__22641;
    wire N__22638;
    wire N__22637;
    wire N__22636;
    wire N__22635;
    wire N__22632;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22603;
    wire N__22596;
    wire N__22591;
    wire N__22588;
    wire N__22583;
    wire N__22578;
    wire N__22575;
    wire N__22556;
    wire N__22555;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22522;
    wire N__22521;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22504;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22459;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22432;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22399;
    wire N__22396;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22384;
    wire N__22379;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22371;
    wire N__22368;
    wire N__22363;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22351;
    wire N__22350;
    wire N__22349;
    wire N__22346;
    wire N__22339;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22306;
    wire N__22305;
    wire N__22302;
    wire N__22297;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22282;
    wire N__22279;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22267;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22186;
    wire N__22185;
    wire N__22182;
    wire N__22177;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22165;
    wire N__22162;
    wire N__22161;
    wire N__22158;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22120;
    wire N__22117;
    wire N__22116;
    wire N__22113;
    wire N__22112;
    wire N__22109;
    wire N__22104;
    wire N__22101;
    wire N__22094;
    wire N__22091;
    wire N__22090;
    wire N__22087;
    wire N__22086;
    wire N__22083;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22060;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22045;
    wire N__22042;
    wire N__22041;
    wire N__22038;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21958;
    wire N__21955;
    wire N__21954;
    wire N__21951;
    wire N__21950;
    wire N__21947;
    wire N__21942;
    wire N__21939;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21904;
    wire N__21901;
    wire N__21900;
    wire N__21897;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21835;
    wire N__21832;
    wire N__21831;
    wire N__21828;
    wire N__21827;
    wire N__21824;
    wire N__21819;
    wire N__21816;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21746;
    wire N__21745;
    wire N__21744;
    wire N__21741;
    wire N__21740;
    wire N__21737;
    wire N__21736;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21716;
    wire N__21713;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21646;
    wire N__21645;
    wire N__21642;
    wire N__21641;
    wire N__21638;
    wire N__21633;
    wire N__21630;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21583;
    wire N__21582;
    wire N__21579;
    wire N__21578;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21562;
    wire N__21559;
    wire N__21558;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21538;
    wire N__21533;
    wire N__21530;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21055;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21025;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21013;
    wire N__21008;
    wire N__21005;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20971;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20959;
    wire N__20954;
    wire N__20951;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20939;
    wire N__20936;
    wire N__20935;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20900;
    wire N__20897;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20882;
    wire N__20879;
    wire N__20878;
    wire N__20875;
    wire N__20872;
    wire N__20867;
    wire N__20864;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20852;
    wire N__20849;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20837;
    wire N__20834;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20822;
    wire N__20819;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20792;
    wire N__20789;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20774;
    wire N__20771;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20759;
    wire N__20756;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20744;
    wire N__20741;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20729;
    wire N__20726;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20711;
    wire N__20708;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20696;
    wire N__20693;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20681;
    wire N__20678;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20663;
    wire N__20660;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20615;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20539;
    wire N__20536;
    wire N__20535;
    wire N__20532;
    wire N__20531;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20517;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20440;
    wire N__20437;
    wire N__20436;
    wire N__20433;
    wire N__20432;
    wire N__20429;
    wire N__20424;
    wire N__20421;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20395;
    wire N__20392;
    wire N__20391;
    wire N__20388;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20245;
    wire N__20242;
    wire N__20241;
    wire N__20240;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20171;
    wire N__20170;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20107;
    wire N__20106;
    wire N__20105;
    wire N__20104;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20096;
    wire N__20095;
    wire N__20094;
    wire N__20093;
    wire N__20090;
    wire N__20089;
    wire N__20088;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20080;
    wire N__20079;
    wire N__20078;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20045;
    wire N__20040;
    wire N__20039;
    wire N__20038;
    wire N__20037;
    wire N__20036;
    wire N__20033;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20008;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19965;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19846;
    wire N__19845;
    wire N__19842;
    wire N__19841;
    wire N__19840;
    wire N__19835;
    wire N__19832;
    wire N__19827;
    wire N__19824;
    wire N__19817;
    wire N__19816;
    wire N__19813;
    wire N__19812;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19787;
    wire N__19784;
    wire N__19783;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19767;
    wire N__19764;
    wire N__19759;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19696;
    wire N__19695;
    wire N__19692;
    wire N__19687;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19651;
    wire N__19650;
    wire N__19645;
    wire N__19642;
    wire N__19637;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19576;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19483;
    wire N__19482;
    wire N__19481;
    wire N__19476;
    wire N__19471;
    wire N__19466;
    wire N__19463;
    wire N__19462;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19447;
    wire N__19446;
    wire N__19445;
    wire N__19442;
    wire N__19441;
    wire N__19440;
    wire N__19439;
    wire N__19438;
    wire N__19437;
    wire N__19434;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19418;
    wire N__19413;
    wire N__19408;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19349;
    wire N__19348;
    wire N__19345;
    wire N__19344;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19312;
    wire N__19311;
    wire N__19310;
    wire N__19305;
    wire N__19300;
    wire N__19295;
    wire N__19294;
    wire N__19291;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19274;
    wire N__19273;
    wire N__19272;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19258;
    wire N__19255;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19243;
    wire N__19240;
    wire N__19239;
    wire N__19236;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19173;
    wire N__19170;
    wire N__19169;
    wire N__19166;
    wire N__19161;
    wire N__19158;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19132;
    wire N__19129;
    wire N__19128;
    wire N__19125;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19051;
    wire N__19048;
    wire N__19047;
    wire N__19044;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18970;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18934;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18847;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18814;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18787;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18748;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18703;
    wire N__18700;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18682;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18634;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18616;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18543;
    wire N__18538;
    wire N__18535;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18508;
    wire N__18505;
    wire N__18504;
    wire N__18501;
    wire N__18500;
    wire N__18497;
    wire N__18492;
    wire N__18489;
    wire N__18482;
    wire N__18479;
    wire N__18478;
    wire N__18475;
    wire N__18474;
    wire N__18473;
    wire N__18472;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18455;
    wire N__18452;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18358;
    wire N__18355;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18319;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18309;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18286;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18244;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18232;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18157;
    wire N__18154;
    wire N__18153;
    wire N__18150;
    wire N__18149;
    wire N__18146;
    wire N__18141;
    wire N__18138;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18004;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17959;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17924;
    wire N__17923;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17905;
    wire N__17904;
    wire N__17903;
    wire N__17900;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17892;
    wire N__17889;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17863;
    wire N__17860;
    wire N__17857;
    wire N__17852;
    wire N__17849;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17821;
    wire N__17818;
    wire N__17815;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17786;
    wire N__17785;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17743;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17731;
    wire N__17730;
    wire N__17729;
    wire N__17728;
    wire N__17727;
    wire N__17726;
    wire N__17725;
    wire N__17724;
    wire N__17723;
    wire N__17722;
    wire N__17721;
    wire N__17718;
    wire N__17717;
    wire N__17716;
    wire N__17715;
    wire N__17714;
    wire N__17713;
    wire N__17712;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17708;
    wire N__17705;
    wire N__17704;
    wire N__17701;
    wire N__17700;
    wire N__17699;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17683;
    wire N__17682;
    wire N__17675;
    wire N__17662;
    wire N__17653;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17628;
    wire N__17625;
    wire N__17620;
    wire N__17615;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17579;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17575;
    wire N__17572;
    wire N__17571;
    wire N__17570;
    wire N__17569;
    wire N__17568;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17564;
    wire N__17561;
    wire N__17550;
    wire N__17547;
    wire N__17544;
    wire N__17543;
    wire N__17542;
    wire N__17541;
    wire N__17532;
    wire N__17529;
    wire N__17524;
    wire N__17519;
    wire N__17516;
    wire N__17511;
    wire N__17508;
    wire N__17503;
    wire N__17500;
    wire N__17489;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17438;
    wire N__17437;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17405;
    wire N__17402;
    wire N__17401;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17383;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17293;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17281;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17263;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17245;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17230;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17209;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17191;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17152;
    wire N__17151;
    wire N__17150;
    wire N__17149;
    wire N__17148;
    wire N__17147;
    wire N__17146;
    wire N__17145;
    wire N__17144;
    wire N__17143;
    wire N__17142;
    wire N__17141;
    wire N__17140;
    wire N__17139;
    wire N__17132;
    wire N__17123;
    wire N__17114;
    wire N__17113;
    wire N__17110;
    wire N__17109;
    wire N__17102;
    wire N__17095;
    wire N__17088;
    wire N__17085;
    wire N__17082;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17062;
    wire N__17057;
    wire N__17054;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17014;
    wire N__17013;
    wire N__17010;
    wire N__17009;
    wire N__17006;
    wire N__17001;
    wire N__16998;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16972;
    wire N__16969;
    wire N__16968;
    wire N__16965;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16939;
    wire N__16938;
    wire N__16935;
    wire N__16934;
    wire N__16931;
    wire N__16926;
    wire N__16923;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16909;
    wire N__16906;
    wire N__16905;
    wire N__16902;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16867;
    wire N__16864;
    wire N__16863;
    wire N__16860;
    wire N__16853;
    wire N__16850;
    wire N__16849;
    wire N__16848;
    wire N__16845;
    wire N__16844;
    wire N__16841;
    wire N__16836;
    wire N__16833;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16801;
    wire N__16798;
    wire N__16797;
    wire N__16794;
    wire N__16787;
    wire N__16784;
    wire N__16783;
    wire N__16780;
    wire N__16779;
    wire N__16778;
    wire N__16777;
    wire N__16772;
    wire N__16769;
    wire N__16764;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16738;
    wire N__16735;
    wire N__16734;
    wire N__16731;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16654;
    wire N__16649;
    wire N__16646;
    wire N__16645;
    wire N__16644;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16621;
    wire N__16620;
    wire N__16617;
    wire N__16612;
    wire N__16607;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16595;
    wire N__16592;
    wire N__16591;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16579;
    wire N__16574;
    wire N__16573;
    wire N__16572;
    wire N__16571;
    wire N__16570;
    wire N__16569;
    wire N__16568;
    wire N__16567;
    wire N__16566;
    wire N__16565;
    wire N__16564;
    wire N__16563;
    wire N__16562;
    wire N__16561;
    wire N__16560;
    wire N__16559;
    wire N__16558;
    wire N__16557;
    wire N__16556;
    wire N__16555;
    wire N__16554;
    wire N__16553;
    wire N__16552;
    wire N__16551;
    wire N__16550;
    wire N__16549;
    wire N__16540;
    wire N__16529;
    wire N__16524;
    wire N__16515;
    wire N__16502;
    wire N__16491;
    wire N__16490;
    wire N__16489;
    wire N__16488;
    wire N__16487;
    wire N__16486;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16387;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16375;
    wire N__16374;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16270;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16238;
    wire N__16237;
    wire N__16236;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16216;
    wire N__16215;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16201;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16180;
    wire N__16175;
    wire N__16172;
    wire N__16171;
    wire N__16170;
    wire N__16167;
    wire N__16160;
    wire N__16157;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16114;
    wire N__16111;
    wire N__16110;
    wire N__16107;
    wire N__16106;
    wire N__16105;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16088;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16060;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15980;
    wire N__15977;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15965;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15911;
    wire N__15910;
    wire N__15909;
    wire N__15906;
    wire N__15901;
    wire N__15898;
    wire N__15893;
    wire N__15892;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15854;
    wire N__15851;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15832;
    wire N__15829;
    wire N__15826;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15808;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15790;
    wire N__15785;
    wire N__15784;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15769;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15756;
    wire N__15749;
    wire N__15748;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15722;
    wire N__15721;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15709;
    wire N__15708;
    wire N__15705;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15680;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15661;
    wire N__15658;
    wire N__15657;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15645;
    wire N__15642;
    wire N__15635;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15617;
    wire N__15614;
    wire N__15613;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15598;
    wire N__15593;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15506;
    wire N__15503;
    wire N__15502;
    wire N__15501;
    wire N__15500;
    wire N__15499;
    wire N__15494;
    wire N__15491;
    wire N__15486;
    wire N__15479;
    wire N__15478;
    wire N__15477;
    wire N__15474;
    wire N__15469;
    wire N__15466;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15451;
    wire N__15448;
    wire N__15447;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15397;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15379;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15364;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15349;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15334;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15301;
    wire N__15298;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15205;
    wire N__15202;
    wire N__15201;
    wire N__15198;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15093;
    wire N__15090;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15010;
    wire N__15009;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14975;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14960;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire VCCG0;
    wire GNDG0;
    wire \b2v_inst16.count_rst_12_cascade_ ;
    wire \b2v_inst16.count_rst_13_cascade_ ;
    wire \b2v_inst16.count_rst_14_cascade_ ;
    wire \b2v_inst16.countZ0Z_9_cascade_ ;
    wire \b2v_inst16.count_4_9 ;
    wire \b2v_inst16.count_rst_6_cascade_ ;
    wire \b2v_inst16.countZ0Z_1_cascade_ ;
    wire \b2v_inst16.count_4_1 ;
    wire \b2v_inst16.count_4_11 ;
    wire \b2v_inst16.count_rst_0_cascade_ ;
    wire \b2v_inst16.countZ0Z_11_cascade_ ;
    wire \b2v_inst16.count_4_8 ;
    wire \b2v_inst16.count_4_6 ;
    wire \b2v_inst16.count_4_15 ;
    wire \b2v_inst200.un25_clk_100khz_1_cascade_ ;
    wire \b2v_inst200.countZ0Z_16 ;
    wire \b2v_inst200.un25_clk_100khz_0 ;
    wire \b2v_inst200.count_RNIZ0Z_1 ;
    wire \b2v_inst200.count_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst200.un2_count_1_axb_1_cascade_ ;
    wire \b2v_inst200.count_3_1 ;
    wire \b2v_inst200.count_3_2 ;
    wire \b2v_inst200.count_3_4 ;
    wire \b2v_inst200.un2_count_1_axb_1 ;
    wire bfn_1_6_0_;
    wire \b2v_inst200.countZ0Z_2 ;
    wire \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_1 ;
    wire \b2v_inst200.un2_count_1_cry_2 ;
    wire \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_3 ;
    wire \b2v_inst200.un2_count_1_cry_4 ;
    wire \b2v_inst200.un2_count_1_cry_5_cZ0 ;
    wire \b2v_inst200.un2_count_1_cry_6 ;
    wire \b2v_inst200.un2_count_1_cry_7 ;
    wire \b2v_inst200.un2_count_1_cry_8 ;
    wire bfn_1_7_0_;
    wire \b2v_inst200.un2_count_1_cry_9 ;
    wire \b2v_inst200.un2_count_1_cry_10 ;
    wire \b2v_inst200.un2_count_1_cry_11 ;
    wire \b2v_inst200.un2_count_1_cry_12 ;
    wire \b2v_inst200.un2_count_1_cry_13 ;
    wire \b2v_inst200.un2_count_1_cry_14 ;
    wire \b2v_inst200.un2_count_1_axb_16 ;
    wire \b2v_inst200.count_1_16 ;
    wire \b2v_inst200.un2_count_1_cry_15 ;
    wire \b2v_inst200.un2_count_1_cry_16 ;
    wire bfn_1_8_0_;
    wire bfn_1_9_0_;
    wire \b2v_inst11.mult1_un68_sum_cry_2 ;
    wire \b2v_inst11.mult1_un68_sum_cry_3 ;
    wire \b2v_inst11.mult1_un68_sum_cry_4 ;
    wire \b2v_inst11.mult1_un68_sum_cry_5 ;
    wire \b2v_inst11.mult1_un68_sum_cry_6 ;
    wire \b2v_inst11.mult1_un68_sum_cry_7 ;
    wire \b2v_inst11.mult1_un68_sum_s_8_cascade_ ;
    wire bfn_1_10_0_;
    wire \b2v_inst11.mult1_un75_sum_cry_2 ;
    wire \b2v_inst11.mult1_un68_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_3 ;
    wire \b2v_inst11.mult1_un68_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_4 ;
    wire \b2v_inst11.mult1_un68_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_5 ;
    wire \b2v_inst11.mult1_un68_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un68_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6 ;
    wire \b2v_inst11.mult1_un75_sum_axb_8 ;
    wire \b2v_inst11.mult1_un75_sum_cry_7 ;
    wire \b2v_inst11.mult1_un75_sum_s_8_cascade_ ;
    wire bfn_1_11_0_;
    wire \b2v_inst11.mult1_un89_sum_cry_2 ;
    wire \b2v_inst11.mult1_un89_sum_cry_3 ;
    wire \b2v_inst11.mult1_un89_sum_cry_4 ;
    wire \b2v_inst11.mult1_un89_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6 ;
    wire \b2v_inst11.mult1_un89_sum_cry_7 ;
    wire \b2v_inst11.mult1_un89_sum_s_8_cascade_ ;
    wire bfn_1_12_0_;
    wire \b2v_inst11.mult1_un96_sum_cry_2 ;
    wire \b2v_inst11.mult1_un89_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_3 ;
    wire \b2v_inst11.mult1_un89_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_4 ;
    wire \b2v_inst11.mult1_un89_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un89_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_6 ;
    wire \b2v_inst11.mult1_un96_sum_axb_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_7 ;
    wire \b2v_inst11.mult1_un96_sum_s_8_cascade_ ;
    wire \b2v_inst11.count_0_8 ;
    wire \b2v_inst11.count_0_9 ;
    wire \b2v_inst11.count_0_10 ;
    wire \b2v_inst11.count_0_11 ;
    wire \b2v_inst11.count_1_1_cascade_ ;
    wire \b2v_inst11.countZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_0_1 ;
    wire \b2v_inst11.count_0_2 ;
    wire \b2v_inst11.count_0_12 ;
    wire bfn_1_15_0_;
    wire \b2v_inst11.count_1_2 ;
    wire \b2v_inst11.un1_count_cry_1_cZ0 ;
    wire \b2v_inst11.un1_count_cry_2 ;
    wire \b2v_inst11.un1_count_cry_3 ;
    wire \b2v_inst11.un1_count_cry_4 ;
    wire \b2v_inst11.un1_count_cry_5 ;
    wire \b2v_inst11.un1_count_cry_6 ;
    wire \b2v_inst11.count_1_8 ;
    wire \b2v_inst11.un1_count_cry_7 ;
    wire \b2v_inst11.un1_count_cry_8 ;
    wire \b2v_inst11.count_1_9 ;
    wire bfn_1_16_0_;
    wire \b2v_inst11.count_1_10 ;
    wire \b2v_inst11.un1_count_cry_9 ;
    wire \b2v_inst11.count_1_11 ;
    wire \b2v_inst11.un1_count_cry_10 ;
    wire \b2v_inst11.count_1_12 ;
    wire \b2v_inst11.un1_count_cry_11 ;
    wire \b2v_inst11.un1_count_cry_12 ;
    wire \b2v_inst11.un1_count_cry_13 ;
    wire \b2v_inst11.un1_count_cry_14 ;
    wire \b2v_inst16.count_rst_9_cascade_ ;
    wire \b2v_inst16.countZ0Z_4_cascade_ ;
    wire \b2v_inst16.count_4_4 ;
    wire \b2v_inst16.count_rst_10_cascade_ ;
    wire \b2v_inst16.countZ0Z_5_cascade_ ;
    wire \b2v_inst16.count_4_5 ;
    wire \b2v_inst16.count_4_7 ;
    wire \b2v_inst16.countZ0Z_2_cascade_ ;
    wire \b2v_inst16.count_4_i_a3_8_0 ;
    wire \b2v_inst16.count_4_i_a3_9_0_cascade_ ;
    wire \b2v_inst16.count_4_i_a3_7_0 ;
    wire \b2v_inst16.count_rst_5 ;
    wire \b2v_inst16.countZ0Z_0_cascade_ ;
    wire \b2v_inst16.N_414 ;
    wire \b2v_inst16.count_4_0 ;
    wire \b2v_inst16.count_4_2 ;
    wire \b2v_inst16.countZ0Z_0 ;
    wire \b2v_inst16.countZ0Z_1 ;
    wire bfn_2_3_0_;
    wire \b2v_inst16.un4_count_1_axb_2 ;
    wire \b2v_inst16.un4_count_1_cry_1_c_RNIAGMEZ0 ;
    wire \b2v_inst16.un4_count_1_cry_1 ;
    wire \b2v_inst16.un4_count_1_cry_2 ;
    wire \b2v_inst16.countZ0Z_4 ;
    wire \b2v_inst16.un4_count_1_cry_3_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_3 ;
    wire \b2v_inst16.countZ0Z_5 ;
    wire \b2v_inst16.un4_count_1_cry_4_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_4 ;
    wire \b2v_inst16.countZ0Z_6 ;
    wire \b2v_inst16.count_rst_11 ;
    wire \b2v_inst16.un4_count_1_cry_5 ;
    wire \b2v_inst16.countZ0Z_7 ;
    wire \b2v_inst16.un4_count_1_cry_6_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_6 ;
    wire \b2v_inst16.countZ0Z_8 ;
    wire \b2v_inst16.un4_count_1_cry_7_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_7 ;
    wire \b2v_inst16.un4_count_1_cry_8 ;
    wire \b2v_inst16.countZ0Z_9 ;
    wire \b2v_inst16.un4_count_1_cry_8_THRU_CO ;
    wire bfn_2_4_0_;
    wire \b2v_inst16.un4_count_1_cry_9 ;
    wire \b2v_inst16.countZ0Z_11 ;
    wire \b2v_inst16.un4_count_1_cry_10_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_10 ;
    wire \b2v_inst16.un4_count_1_cry_11 ;
    wire \b2v_inst16.un4_count_1_cry_12 ;
    wire \b2v_inst16.un4_count_1_cry_13 ;
    wire \b2v_inst16.countZ0Z_15 ;
    wire \b2v_inst16.un4_count_1_cry_14 ;
    wire \b2v_inst16.count_rst_4 ;
    wire \b2v_inst200.count_3_14 ;
    wire \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ;
    wire \b2v_inst200.count_3_6 ;
    wire \b2v_inst200.count_1_6 ;
    wire \b2v_inst200.count_3_7 ;
    wire \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ;
    wire \b2v_inst200.count_0_17 ;
    wire \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ;
    wire \b2v_inst200.countZ0Z_17 ;
    wire \b2v_inst200.count_1_10 ;
    wire \b2v_inst200.count_3_10 ;
    wire \b2v_inst200.count_1_0 ;
    wire \b2v_inst200.countZ0Z_10 ;
    wire \b2v_inst200.count_1_8 ;
    wire \b2v_inst200.count_3_8 ;
    wire \b2v_inst200.un2_count_1_axb_8 ;
    wire \b2v_inst200.un2_count_1_axb_15 ;
    wire \b2v_inst200.count_3_15 ;
    wire \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71 ;
    wire \b2v_inst200.countZ0Z_6 ;
    wire \b2v_inst200.un25_clk_100khz_7 ;
    wire \b2v_inst200.un25_clk_100khz_13 ;
    wire \b2v_inst200.un25_clk_100khz_6_cascade_ ;
    wire \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_ ;
    wire \b2v_inst200.countZ0Z_0 ;
    wire \b2v_inst200.count_3_0 ;
    wire \b2v_inst200.un2_count_1_axb_9 ;
    wire \b2v_inst200.count_3_12 ;
    wire \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ;
    wire \b2v_inst200.countZ0Z_12 ;
    wire \b2v_inst200.count_3_9 ;
    wire \b2v_inst200.countZ0Z_12_cascade_ ;
    wire \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ;
    wire \b2v_inst200.un2_count_1_axb_5 ;
    wire \b2v_inst200.count_3_11 ;
    wire \b2v_inst200.count_1_11 ;
    wire \b2v_inst200.countZ0Z_11 ;
    wire \b2v_inst200.un2_count_1_axb_3 ;
    wire \b2v_inst200.countZ0Z_14 ;
    wire \b2v_inst200.un25_clk_100khz_4 ;
    wire \b2v_inst200.un25_clk_100khz_5_cascade_ ;
    wire \b2v_inst200.un25_clk_100khz_14 ;
    wire \b2v_inst200.count_3_3 ;
    wire \b2v_inst200.countZ0Z_4 ;
    wire \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ;
    wire \b2v_inst200.un25_clk_100khz_2 ;
    wire \b2v_inst200.count_3_13 ;
    wire \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ;
    wire \b2v_inst200.un2_count_1_axb_13 ;
    wire \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ;
    wire \b2v_inst200.count_3_5 ;
    wire \b2v_inst200.countZ0Z_7 ;
    wire \b2v_inst200.count_en_g ;
    wire \b2v_inst200.un25_clk_100khz_3 ;
    wire bfn_2_9_0_;
    wire \b2v_inst11.mult1_un61_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_2 ;
    wire \b2v_inst11.mult1_un61_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_3 ;
    wire \b2v_inst11.mult1_un61_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_4 ;
    wire \b2v_inst11.mult1_un61_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_5 ;
    wire \b2v_inst11.mult1_un68_sum_axb_8 ;
    wire \b2v_inst11.mult1_un61_sum_cry_6 ;
    wire \b2v_inst11.mult1_un61_sum_cry_7 ;
    wire \b2v_inst11.mult1_un61_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un61_sum_i_0_8 ;
    wire bfn_2_10_0_;
    wire \b2v_inst11.mult1_un82_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_2 ;
    wire \b2v_inst11.mult1_un75_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_3 ;
    wire \b2v_inst11.mult1_un75_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_4 ;
    wire \b2v_inst11.mult1_un75_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_5 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un75_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un89_sum_axb_8 ;
    wire \b2v_inst11.mult1_un82_sum_cry_6 ;
    wire \b2v_inst11.mult1_un82_sum_axb_8 ;
    wire \b2v_inst11.mult1_un82_sum_cry_7 ;
    wire \b2v_inst11.mult1_un54_sum_i_8 ;
    wire \b2v_inst11.mult1_un75_sum_s_8 ;
    wire \b2v_inst11.mult1_un68_sum_i ;
    wire \b2v_inst11.mult1_un82_sum_i ;
    wire \b2v_inst11.mult1_un89_sum_i ;
    wire \b2v_inst11.mult1_un82_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un82_sum_s_8 ;
    wire bfn_2_12_0_;
    wire \b2v_inst11.mult1_un103_sum_cry_2 ;
    wire \b2v_inst11.mult1_un96_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_3 ;
    wire \b2v_inst11.mult1_un96_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_4 ;
    wire \b2v_inst11.mult1_un96_sum_s_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_5 ;
    wire \b2v_inst11.mult1_un96_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un96_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un103_sum_cry_6 ;
    wire \b2v_inst11.mult1_un103_sum_axb_8 ;
    wire \b2v_inst11.mult1_un103_sum_cry_7 ;
    wire \b2v_inst11.mult1_un89_sum_s_8 ;
    wire pwrbtn_led;
    wire \b2v_inst11.curr_state_3_0_cascade_ ;
    wire \b2v_inst11.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_0_sqmuxa_i ;
    wire \b2v_inst11.count_0_sqmuxa_i_cascade_ ;
    wire \b2v_inst11.count_1_0_cascade_ ;
    wire \b2v_inst11.count_0_0 ;
    wire \b2v_inst11.pwm_outZ0 ;
    wire \b2v_inst11.g0_i_o3_0 ;
    wire \b2v_inst11.count_1_3 ;
    wire \b2v_inst11.count_0_3 ;
    wire \b2v_inst11.count_1_13 ;
    wire \b2v_inst11.count_0_13 ;
    wire \b2v_inst11.count_1_4 ;
    wire \b2v_inst11.count_0_4 ;
    wire \b2v_inst11.count_1_5 ;
    wire \b2v_inst11.count_0_5 ;
    wire \b2v_inst11.pwm_out_1_sqmuxa ;
    wire \b2v_inst11.un79_clk_100khzlt6_cascade_ ;
    wire \b2v_inst11.un79_clk_100khzlto15_5_cascade_ ;
    wire \b2v_inst11.un79_clk_100khzlto15_7_cascade_ ;
    wire \b2v_inst11.un79_clk_100khzlto15_3 ;
    wire \b2v_inst11.count_RNIZ0Z_8_cascade_ ;
    wire \b2v_inst11.N_8 ;
    wire \b2v_inst11.count_1_14 ;
    wire \b2v_inst11.count_0_14 ;
    wire \b2v_inst11.count_1_6 ;
    wire \b2v_inst11.count_0_6 ;
    wire \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ;
    wire \b2v_inst11.count_0_15 ;
    wire \b2v_inst11.count_1_7 ;
    wire \b2v_inst11.count_0_7 ;
    wire \b2v_inst200.count_enZ0 ;
    wire pch_pwrok;
    wire vpp_en;
    wire \b2v_inst16.delayed_vddq_pwrgd_eZ0Z_0 ;
    wire \b2v_inst16.delayed_vddq_pwrgd_en ;
    wire \b2v_inst16.N_26 ;
    wire \b2v_inst16.N_416 ;
    wire \b2v_inst16.un4_count_1_cry_2_THRU_CO ;
    wire \b2v_inst16.N_26_cascade_ ;
    wire \b2v_inst16.count_4_i_a3_10_0 ;
    wire \b2v_inst16.countZ0Z_14 ;
    wire \b2v_inst16.count_rst_3 ;
    wire \b2v_inst16.count_4_14 ;
    wire \b2v_inst16.countZ0Z_12 ;
    wire \b2v_inst16.count_rst_1 ;
    wire \b2v_inst16.count_4_12 ;
    wire \b2v_inst16.countZ0Z_13 ;
    wire \b2v_inst16.count_rst_2 ;
    wire \b2v_inst16.count_4_13 ;
    wire \b2v_inst16.N_3079_i ;
    wire \b2v_inst16.count_4_3 ;
    wire \b2v_inst16.count_rst_8 ;
    wire \b2v_inst16.countZ0Z_3 ;
    wire \b2v_inst11.dutycycleZ1Z_7 ;
    wire \b2v_inst11.dutycycleZ1Z_3_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_7_1_cascade_ ;
    wire \b2v_inst16.curr_state_2_1 ;
    wire \b2v_inst16.curr_state_7_0_1 ;
    wire \b2v_inst11.un1_dutycycle_53_44_0_2_cascade_ ;
    wire \b2v_inst11.un2_count_clk_17_0_a2_1_4 ;
    wire \b2v_inst11.N_355_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_55_1_tz ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_11_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_50_a0_1 ;
    wire \b2v_inst11.un1_dutycycle_53_50_a0_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_6_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_12_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_4_1 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_12 ;
    wire \b2v_inst11.un1_dutycycle_53_4_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_6_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_9Z0Z_7 ;
    wire \b2v_inst11.un1_dutycycle_53_46_0_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_11_1_0 ;
    wire bfn_4_9_0_;
    wire \b2v_inst11.mult1_un54_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_2 ;
    wire \b2v_inst11.mult1_un54_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_3 ;
    wire \b2v_inst11.mult1_un54_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_4 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_5 ;
    wire \b2v_inst11.mult1_un61_sum_axb_8 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6 ;
    wire \b2v_inst11.mult1_un54_sum_cry_7 ;
    wire \b2v_inst11.mult1_un54_sum_s_8 ;
    wire \b2v_inst11.mult1_un47_sum_l_fx_3 ;
    wire vpp_ok;
    wire vddq_en;
    wire \b2v_inst11.mult1_un54_sum_i ;
    wire \b2v_inst11.mult1_un61_sum_s_8 ;
    wire \b2v_inst11.mult1_un61_sum_i ;
    wire \b2v_inst11.mult1_un75_sum_i ;
    wire \b2v_inst11.mult1_un68_sum_s_8 ;
    wire \b2v_inst11.countZ0Z_0 ;
    wire \b2v_inst11.N_5980_i ;
    wire bfn_4_11_0_;
    wire \b2v_inst11.countZ0Z_1 ;
    wire \b2v_inst11.N_5981_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_0 ;
    wire \b2v_inst11.countZ0Z_2 ;
    wire \b2v_inst11.N_5982_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_1 ;
    wire \b2v_inst11.countZ0Z_3 ;
    wire \b2v_inst11.N_5983_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_2 ;
    wire \b2v_inst11.countZ0Z_4 ;
    wire \b2v_inst11.N_5984_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_3 ;
    wire \b2v_inst11.countZ0Z_5 ;
    wire \b2v_inst11.N_5985_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_4 ;
    wire \b2v_inst11.countZ0Z_6 ;
    wire \b2v_inst11.N_5986_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_5 ;
    wire \b2v_inst11.countZ0Z_7 ;
    wire \b2v_inst11.N_5987_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_6 ;
    wire \b2v_inst11.un85_clk_100khz_cry_7 ;
    wire \b2v_inst11.countZ0Z_8 ;
    wire \b2v_inst11.N_5988_i ;
    wire bfn_4_12_0_;
    wire \b2v_inst11.countZ0Z_9 ;
    wire \b2v_inst11.N_5989_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_8 ;
    wire \b2v_inst11.mult1_un96_sum_i_8 ;
    wire \b2v_inst11.countZ0Z_10 ;
    wire \b2v_inst11.N_5990_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_9 ;
    wire \b2v_inst11.mult1_un89_sum_i_8 ;
    wire \b2v_inst11.countZ0Z_11 ;
    wire \b2v_inst11.N_5991_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_10 ;
    wire \b2v_inst11.countZ0Z_12 ;
    wire \b2v_inst11.mult1_un82_sum_i_8 ;
    wire \b2v_inst11.N_5992_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_11 ;
    wire \b2v_inst11.mult1_un75_sum_i_8 ;
    wire \b2v_inst11.countZ0Z_13 ;
    wire \b2v_inst11.N_5993_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_12 ;
    wire \b2v_inst11.mult1_un68_sum_i_8 ;
    wire \b2v_inst11.countZ0Z_14 ;
    wire \b2v_inst11.N_5994_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_13 ;
    wire \b2v_inst11.countZ0Z_15 ;
    wire \b2v_inst11.mult1_un61_sum_i_8 ;
    wire \b2v_inst11.N_5995_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_14 ;
    wire \b2v_inst11.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_4_13_0_;
    wire \b2v_inst11.mult1_un110_sum_i_8 ;
    wire bfn_4_14_0_;
    wire \b2v_inst11.mult1_un103_sum_i ;
    wire \b2v_inst11.mult1_un110_sum_cry_2 ;
    wire \b2v_inst11.mult1_un103_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_3 ;
    wire \b2v_inst11.mult1_un103_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_4 ;
    wire \b2v_inst11.mult1_un103_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_5 ;
    wire \b2v_inst11.mult1_un103_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un103_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un110_sum_cry_6 ;
    wire \b2v_inst11.mult1_un110_sum_axb_8 ;
    wire \b2v_inst11.mult1_un110_sum_cry_7 ;
    wire \b2v_inst11.mult1_un110_sum_s_8_cascade_ ;
    wire bfn_4_15_0_;
    wire \b2v_inst11.mult1_un117_sum_cry_2 ;
    wire \b2v_inst11.mult1_un110_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_3 ;
    wire \b2v_inst11.mult1_un110_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_4 ;
    wire \b2v_inst11.mult1_un110_sum_s_8 ;
    wire \b2v_inst11.mult1_un110_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_5 ;
    wire \b2v_inst11.mult1_un110_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un110_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un117_sum_cry_6 ;
    wire \b2v_inst11.mult1_un117_sum_axb_8 ;
    wire \b2v_inst11.mult1_un117_sum_cry_7 ;
    wire \b2v_inst11.mult1_un117_sum_s_8_cascade_ ;
    wire bfn_4_16_0_;
    wire \b2v_inst11.mult1_un166_sum_cry_0 ;
    wire \b2v_inst11.mult1_un166_sum_cry_1 ;
    wire \b2v_inst11.mult1_un166_sum_cry_2 ;
    wire \b2v_inst11.mult1_un166_sum_cry_3 ;
    wire G_2814;
    wire \b2v_inst11.mult1_un166_sum_cry_4 ;
    wire \b2v_inst11.mult1_un166_sum_cry_5 ;
    wire \b2v_inst11.un85_clk_100khz_0 ;
    wire \b2v_inst200.N_58_cascade_ ;
    wire \b2v_inst200.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst200.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst200.N_56 ;
    wire gpio_fpga_soc_1;
    wire \b2v_inst200.m6_i_0 ;
    wire N_411;
    wire \b2v_inst200.m6_i_0_cascade_ ;
    wire \b2v_inst200.count_RNI5RUP8Z0Z_8 ;
    wire \b2v_inst200.curr_state_3_0 ;
    wire \b2v_inst200.curr_stateZ0Z_2 ;
    wire \b2v_inst200.i4_mux_cascade_ ;
    wire \b2v_inst200.curr_state_i_2_cascade_ ;
    wire hda_sdo_atp;
    wire \b2v_inst200.N_3031_i ;
    wire \b2v_inst200.N_205 ;
    wire \b2v_inst200.curr_state_i_2 ;
    wire \b2v_inst200.N_205_cascade_ ;
    wire \b2v_inst200.HDA_SDO_ATP_0 ;
    wire \b2v_inst200.curr_stateZ0Z_0 ;
    wire \b2v_inst200.curr_stateZ0Z_1 ;
    wire \b2v_inst200.N_282 ;
    wire \b2v_inst200.curr_state_3_1 ;
    wire \b2v_inst16.curr_state_2_0 ;
    wire bfn_5_4_0_;
    wire \b2v_inst20.un4_counter_0 ;
    wire \b2v_inst20.un4_counter_2_and ;
    wire \b2v_inst20.un4_counter_1 ;
    wire \b2v_inst20.un4_counter_3_and ;
    wire \b2v_inst20.un4_counter_2 ;
    wire \b2v_inst20.un4_counter_4_and ;
    wire \b2v_inst20.un4_counter_3 ;
    wire \b2v_inst20.un4_counter_5_and ;
    wire \b2v_inst20.un4_counter_4 ;
    wire \b2v_inst20.un4_counter_5 ;
    wire \b2v_inst20.un4_counter_6 ;
    wire b2v_inst20_un4_counter_7;
    wire bfn_5_5_0_;
    wire \b2v_inst11.un1_dutycycle_53_axb_11_1 ;
    wire \b2v_inst11.un1_dutycycle_53_39_0_1_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_7 ;
    wire \b2v_inst20.un4_counter_6_and ;
    wire \b2v_inst11.un1_dutycycle_53_39_d_0_0 ;
    wire \b2v_inst11.dutycycle_RNITSFK3Z0Z_10_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI9LPN6Z0Z_10 ;
    wire \b2v_inst11.dutycycleZ0Z_10 ;
    wire \b2v_inst11.dutycycleZ0Z_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNITSFK3Z0Z_9_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9 ;
    wire \b2v_inst11.dutycycle_RNI9LPN6Z0Z_9_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_9 ;
    wire \b2v_inst11.un1_dutycycle_53_30_a1_0_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_44_2 ;
    wire \b2v_inst11.un1_dutycycle_53_5_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_6 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_4 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_8_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_9_1 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_11 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_7 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_8Z0Z_6 ;
    wire bfn_5_9_0_;
    wire \b2v_inst11.mult1_un47_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un47_sum_cry_2 ;
    wire \b2v_inst11.mult1_un47_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un47_sum_cry_3 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un47_sum_cry_4 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5 ;
    wire \b2v_inst11.mult1_un47_sum_l_fx_6 ;
    wire \b2v_inst11.mult1_un47_sum_i ;
    wire \b2v_inst11.un1_dutycycle_53_axb_12 ;
    wire \b2v_inst11.curr_stateZ0Z_0 ;
    wire \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \b2v_inst11.count_RNIZ0Z_8 ;
    wire \b2v_inst11.curr_state_4_0 ;
    wire \b2v_inst11.mult1_un47_sum_s_4_sf ;
    wire \b2v_inst11.mult1_un40_sum_i_l_ofx_4 ;
    wire \b2v_inst11.mult1_un40_sum_i_5 ;
    wire \b2v_inst11.mult1_un40_sum_i_5_cascade_ ;
    wire \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ;
    wire \b2v_inst11.mult1_un47_sum_s_6 ;
    wire \b2v_inst11.un1_dutycycle_53_i_29 ;
    wire \b2v_inst16.count_rst ;
    wire \b2v_inst16.count_4_10 ;
    wire \b2v_inst16.count_en ;
    wire \b2v_inst16.countZ0Z_10 ;
    wire \b2v_inst11.mult1_un110_sum_i ;
    wire \b2v_inst11.mult1_un117_sum_i_8 ;
    wire vccst_en;
    wire \b2v_inst11.un85_clk_100khz_4 ;
    wire \b2v_inst11.mult1_un124_sum_i_8 ;
    wire \b2v_inst11.un85_clk_100khz_2 ;
    wire \b2v_inst11.un85_clk_100khz_1 ;
    wire \b2v_inst11.mult1_un96_sum_i ;
    wire \b2v_inst11.mult1_un131_sum_i_8 ;
    wire \b2v_inst11.un85_clk_100khz_3 ;
    wire \b2v_inst11.mult1_un103_sum_s_8 ;
    wire \b2v_inst11.mult1_un103_sum_i_8 ;
    wire bfn_5_13_0_;
    wire \b2v_inst11.mult1_un124_sum_i ;
    wire \b2v_inst11.mult1_un131_sum_cry_2 ;
    wire \b2v_inst11.mult1_un131_sum_cry_3 ;
    wire \b2v_inst11.mult1_un131_sum_cry_4 ;
    wire \b2v_inst11.mult1_un131_sum_cry_5 ;
    wire \b2v_inst11.mult1_un131_sum_cry_6 ;
    wire \b2v_inst11.mult1_un131_sum_cry_7 ;
    wire \b2v_inst11.mult1_un131_sum_s_8_cascade_ ;
    wire bfn_5_14_0_;
    wire \b2v_inst11.mult1_un117_sum_i ;
    wire \b2v_inst11.mult1_un124_sum_cry_2 ;
    wire \b2v_inst11.mult1_un117_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_3 ;
    wire \b2v_inst11.mult1_un117_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_4 ;
    wire \b2v_inst11.mult1_un117_sum_s_8 ;
    wire \b2v_inst11.mult1_un117_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_5 ;
    wire \b2v_inst11.mult1_un117_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un117_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un131_sum_axb_8 ;
    wire \b2v_inst11.mult1_un124_sum_cry_6 ;
    wire \b2v_inst11.mult1_un124_sum_axb_8 ;
    wire \b2v_inst11.mult1_un124_sum_cry_7 ;
    wire \b2v_inst11.mult1_un124_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un124_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un131_sum_axb_7_l_fx ;
    wire \b2v_inst11.g3_0 ;
    wire bfn_5_15_0_;
    wire \b2v_inst11.mult1_un159_sum_cry_2_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_1 ;
    wire \b2v_inst11.mult1_un159_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_2 ;
    wire \b2v_inst11.mult1_un159_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_3 ;
    wire \b2v_inst11.mult1_un159_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_4 ;
    wire \b2v_inst11.mult1_un166_sum_axb_6 ;
    wire \b2v_inst11.mult1_un159_sum_cry_5 ;
    wire \b2v_inst11.mult1_un159_sum_cry_6 ;
    wire \b2v_inst11.mult1_un159_sum_s_7 ;
    wire \b2v_inst11.mult1_un124_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un159_sum_i ;
    wire bfn_6_2_0_;
    wire \b2v_inst20.counter_1_cry_1 ;
    wire \b2v_inst20.counter_1_cry_2 ;
    wire \b2v_inst20.counter_1_cry_3 ;
    wire \b2v_inst20.counter_1_cry_4 ;
    wire \b2v_inst20.counter_1_cry_5 ;
    wire \b2v_inst20.counter_1_cry_6 ;
    wire \b2v_inst20.counterZ0Z_8 ;
    wire \b2v_inst20.counter_1_cry_7 ;
    wire \b2v_inst20.counter_1_cry_8 ;
    wire \b2v_inst20.counterZ0Z_9 ;
    wire bfn_6_3_0_;
    wire \b2v_inst20.counterZ0Z_10 ;
    wire \b2v_inst20.counter_1_cry_9 ;
    wire \b2v_inst20.counterZ0Z_11 ;
    wire \b2v_inst20.counter_1_cry_10 ;
    wire \b2v_inst20.counterZ0Z_12 ;
    wire \b2v_inst20.counter_1_cry_11 ;
    wire \b2v_inst20.counterZ0Z_13 ;
    wire \b2v_inst20.counter_1_cry_12 ;
    wire \b2v_inst20.counterZ0Z_14 ;
    wire \b2v_inst20.counter_1_cry_13 ;
    wire \b2v_inst20.counterZ0Z_15 ;
    wire \b2v_inst20.counter_1_cry_14 ;
    wire \b2v_inst20.counterZ0Z_16 ;
    wire \b2v_inst20.counter_1_cry_15 ;
    wire \b2v_inst20.counter_1_cry_16 ;
    wire \b2v_inst20.counterZ0Z_17 ;
    wire bfn_6_4_0_;
    wire \b2v_inst20.counterZ0Z_18 ;
    wire \b2v_inst20.counter_1_cry_17 ;
    wire \b2v_inst20.counterZ0Z_19 ;
    wire \b2v_inst20.counter_1_cry_18 ;
    wire \b2v_inst20.counterZ0Z_20 ;
    wire \b2v_inst20.counter_1_cry_19 ;
    wire \b2v_inst20.counterZ0Z_21 ;
    wire \b2v_inst20.counter_1_cry_20 ;
    wire \b2v_inst20.counterZ0Z_22 ;
    wire \b2v_inst20.counter_1_cry_21 ;
    wire \b2v_inst20.counterZ0Z_23 ;
    wire \b2v_inst20.counter_1_cry_22 ;
    wire \b2v_inst20.counterZ0Z_24 ;
    wire \b2v_inst20.counter_1_cry_23 ;
    wire \b2v_inst20.counter_1_cry_24 ;
    wire \b2v_inst20.counterZ0Z_25 ;
    wire bfn_6_5_0_;
    wire \b2v_inst20.counterZ0Z_26 ;
    wire \b2v_inst20.counter_1_cry_25 ;
    wire \b2v_inst20.counterZ0Z_27 ;
    wire \b2v_inst20.counter_1_cry_26 ;
    wire \b2v_inst20.counter_1_cry_27 ;
    wire \b2v_inst20.counter_1_cry_28 ;
    wire \b2v_inst20.counter_1_cry_29 ;
    wire \b2v_inst20.counter_1_cry_30 ;
    wire \b2v_inst20.counterZ0Z_28 ;
    wire \b2v_inst20.counterZ0Z_29 ;
    wire \b2v_inst20.counterZ0Z_30 ;
    wire \b2v_inst20.counterZ0Z_31 ;
    wire \b2v_inst20.un4_counter_7_and ;
    wire \b2v_inst11.un1_dutycycle_53_9_1_1 ;
    wire \b2v_inst11.dutycycleZ1Z_5_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_8 ;
    wire \b2v_inst11.un1_dutycycle_53_3_0_tz ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_3_cascade_ ;
    wire \b2v_inst11.N_26_i_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_9_1 ;
    wire \b2v_inst11.dutycycleZ0Z_13 ;
    wire \b2v_inst11.dutycycleZ1Z_4 ;
    wire \b2v_inst11.dutycycleZ0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_8Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_4_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_8_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_11 ;
    wire \b2v_inst11.un1_dutycycle_53_axb_3_1_0_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_3_cascade_ ;
    wire \b2v_inst11.un1_i3_mux_cascade_ ;
    wire \b2v_inst11.d_i3_mux ;
    wire bfn_6_9_0_;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_1 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_2 ;
    wire \b2v_inst11.mult1_un124_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_2 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_5 ;
    wire \b2v_inst11.mult1_un117_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_3 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_7 ;
    wire \b2v_inst11.mult1_un110_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_4 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_5 ;
    wire \b2v_inst11.mult1_un103_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_5 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_10 ;
    wire \b2v_inst11.mult1_un96_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_6 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_7 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_11 ;
    wire \b2v_inst11.mult1_un89_sum ;
    wire bfn_6_10_0_;
    wire \b2v_inst11.dutycycle_RNIZ0Z_12 ;
    wire \b2v_inst11.mult1_un82_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_8 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_13 ;
    wire \b2v_inst11.mult1_un75_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_9 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_14 ;
    wire \b2v_inst11.mult1_un68_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_10 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_15 ;
    wire \b2v_inst11.mult1_un61_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_11 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_13 ;
    wire \b2v_inst11.mult1_un54_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_12 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_13 ;
    wire \b2v_inst11.mult1_un47_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_13 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_14 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ;
    wire bfn_6_11_0_;
    wire \b2v_inst11.CO2 ;
    wire \b2v_inst11.CO2_THRU_CO ;
    wire \b2v_inst11.mult1_un131_sum ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_14 ;
    wire \b2v_inst5.count_1_6 ;
    wire vr_ready_vccinaux;
    wire vr_ready_vccin;
    wire \b2v_inst11.mult1_un124_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un124_sum_s_8 ;
    wire \b2v_inst11.mult1_un131_sum_axb_4_l_fx ;
    wire \b2v_inst11.mult1_un138_sum ;
    wire bfn_6_13_0_;
    wire \b2v_inst11.mult1_un131_sum_i ;
    wire \b2v_inst11.mult1_un138_sum_cry_2_c ;
    wire \b2v_inst11.mult1_un131_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_3_c ;
    wire \b2v_inst11.mult1_un131_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_4_c ;
    wire \b2v_inst11.mult1_un131_sum_s_8 ;
    wire \b2v_inst11.mult1_un131_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_5_c ;
    wire \b2v_inst11.mult1_un131_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un131_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un138_sum_cry_6_c ;
    wire \b2v_inst11.mult1_un138_sum_axb_8 ;
    wire \b2v_inst11.mult1_un138_sum_cry_7 ;
    wire \b2v_inst11.mult1_un138_sum_s_8_cascade_ ;
    wire bfn_6_14_0_;
    wire \b2v_inst11.mult1_un138_sum_i ;
    wire \b2v_inst11.mult1_un145_sum_cry_2 ;
    wire \b2v_inst11.mult1_un138_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_3 ;
    wire \b2v_inst11.mult1_un138_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_4 ;
    wire \b2v_inst11.mult1_un138_sum_s_8 ;
    wire \b2v_inst11.mult1_un138_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_5 ;
    wire \b2v_inst11.mult1_un138_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un138_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un145_sum_cry_6 ;
    wire \b2v_inst11.mult1_un145_sum_axb_8 ;
    wire \b2v_inst11.mult1_un145_sum_cry_7 ;
    wire \b2v_inst11.mult1_un145_sum_s_8_cascade_ ;
    wire bfn_6_15_0_;
    wire \b2v_inst11.mult1_un152_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_2 ;
    wire \b2v_inst11.mult1_un145_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_3 ;
    wire \b2v_inst11.mult1_un145_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_4 ;
    wire \b2v_inst11.mult1_un145_sum_s_8 ;
    wire \b2v_inst11.mult1_un145_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_5 ;
    wire \b2v_inst11.mult1_un145_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un145_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un159_sum_axb_7 ;
    wire \b2v_inst11.mult1_un152_sum_cry_6 ;
    wire \b2v_inst11.mult1_un152_sum_axb_8 ;
    wire \b2v_inst11.mult1_un152_sum_cry_7 ;
    wire \b2v_inst11.mult1_un152_sum_s_8 ;
    wire \b2v_inst11.mult1_un152_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un152_sum_i_0_8 ;
    wire \b2v_inst36.count_rst_3_cascade_ ;
    wire \b2v_inst36.countZ0Z_11_cascade_ ;
    wire \b2v_inst36.count_2_11 ;
    wire \b2v_inst36.count_2_1 ;
    wire \b2v_inst36.count_2_15 ;
    wire \b2v_inst36.count_2_13 ;
    wire \b2v_inst36.count_2_14 ;
    wire \b2v_inst36.count_i_0 ;
    wire \b2v_inst5.count_1_7 ;
    wire \b2v_inst5.count_1_11 ;
    wire \b2v_inst5.countZ0Z_7_cascade_ ;
    wire \b2v_inst5.count_1_12 ;
    wire \b2v_inst20.counterZ0Z_7 ;
    wire \b2v_inst20.un4_counter_1_and ;
    wire \b2v_inst20.counter_1_cry_5_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_6 ;
    wire \b2v_inst20.counterZ0Z_1 ;
    wire \b2v_inst20.counterZ0Z_0 ;
    wire \b2v_inst20.un4_counter_0_and ;
    wire \b2v_inst20.counter_1_cry_4_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_5 ;
    wire \b2v_inst20.counter_1_cry_3_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_4 ;
    wire bfn_7_5_0_;
    wire \b2v_inst5.un2_count_1_cry_0 ;
    wire \b2v_inst5.un2_count_1_cry_1 ;
    wire \b2v_inst5.un2_count_1_cry_2 ;
    wire \b2v_inst5.un2_count_1_cry_3 ;
    wire \b2v_inst5.un2_count_1_cry_4 ;
    wire \b2v_inst5.count_rst_8 ;
    wire \b2v_inst5.un2_count_1_cry_5 ;
    wire \b2v_inst5.countZ0Z_7 ;
    wire \b2v_inst5.count_rst_7 ;
    wire \b2v_inst5.un2_count_1_cry_6 ;
    wire \b2v_inst5.un2_count_1_cry_7 ;
    wire bfn_7_6_0_;
    wire \b2v_inst5.un2_count_1_cry_8 ;
    wire \b2v_inst5.un2_count_1_cry_9 ;
    wire \b2v_inst5.un2_count_1_axb_11 ;
    wire \b2v_inst5.count_rst_3 ;
    wire \b2v_inst5.un2_count_1_cry_10 ;
    wire \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2 ;
    wire \b2v_inst5.un2_count_1_cry_11 ;
    wire \b2v_inst5.un2_count_1_cry_12 ;
    wire \b2v_inst5.un2_count_1_cry_13 ;
    wire \b2v_inst5.un2_count_1_cry_14 ;
    wire bfn_7_7_0_;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_4 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ;
    wire \b2v_inst11.dutycycleZ1Z_3 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9JZ0Z1 ;
    wire bfn_7_8_0_;
    wire \b2v_inst11.dutycycleZ0Z_1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJZ0Z1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ;
    wire \b2v_inst11.dutycycleZ0Z_4 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJZ0Z1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14 ;
    wire \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_3_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ;
    wire \b2v_inst11.dutycycle_e_1_3 ;
    wire \b2v_inst11.un1_clk_100khz_43_and_i_0_0_0 ;
    wire \b2v_inst11.dutycycle_e_1_3_cascade_ ;
    wire \b2v_inst11.dutycycle_0_3 ;
    wire \b2v_inst11.un1_clk_100khz_40_and_i_0_0_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIT35D7Z0Z_4 ;
    wire \b2v_inst11.N_155_N ;
    wire \b2v_inst11.dutycycle_en_11_cascade_ ;
    wire \b2v_inst11.N_158_N_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIT35D7Z0Z_15 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ;
    wire \b2v_inst11.dutycycle_RNIT35D7Z0Z_15_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_15 ;
    wire \b2v_inst11.dutycycleZ0Z_14 ;
    wire \b2v_inst11.dutycycle_en_11 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ;
    wire \b2v_inst11.dutycycleZ0Z_12 ;
    wire \b2v_inst11.dutycycleZ0Z_12_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_13 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_14 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19 ;
    wire \b2v_inst11.dutycycle_set_1_cascade_ ;
    wire \b2v_inst11.N_300 ;
    wire \b2v_inst11.N_300_0_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29 ;
    wire \b2v_inst11.dutycycle_set_0_0 ;
    wire \b2v_inst11.dutycycle_set_0_0_cascade_ ;
    wire \b2v_inst11.dutycycle_0_6 ;
    wire \b2v_inst11.dutycycle_0_5 ;
    wire \b2v_inst11.dutycycle_set_1 ;
    wire \b2v_inst11.dutycycle_eena_13_0 ;
    wire \b2v_inst11.N_200_i_cascade_ ;
    wire \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_3 ;
    wire \b2v_inst11.dutycycleZ1Z_5 ;
    wire \b2v_inst11.un1_clk_100khz_32_and_i_0_c ;
    wire \b2v_inst11.un1_clk_100khz_40_and_i_0_c ;
    wire \b2v_inst11.dutycycleZ0Z_3 ;
    wire \b2v_inst11.mult1_un145_sum ;
    wire \b2v_inst11.mult1_un145_sum_cascade_ ;
    wire \b2v_inst11.mult1_un145_sum_i ;
    wire \b2v_inst11.N_10 ;
    wire \b2v_inst11.count_clk_0_8 ;
    wire \b2v_inst11.count_clkZ0Z_8_cascade_ ;
    wire \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ;
    wire \b2v_inst11.N_379 ;
    wire \b2v_inst11.N_379_cascade_ ;
    wire \b2v_inst11.count_clk_0_9 ;
    wire \b2v_inst11.count_clkZ0Z_9_cascade_ ;
    wire \b2v_inst11.N_190 ;
    wire \b2v_inst11.count_clk_0_5 ;
    wire \b2v_inst11.count_clkZ0Z_5_cascade_ ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2 ;
    wire \b2v_inst11.count_clkZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_clk_0_1 ;
    wire \b2v_inst11.count_clkZ0Z_15_cascade_ ;
    wire \b2v_inst11.N_175 ;
    wire \b2v_inst11.count_clk_0_14 ;
    wire \b2v_inst11.count_clk_0_15 ;
    wire \b2v_inst36.un2_count_1_axb_3_cascade_ ;
    wire \b2v_inst36.count_rst_11 ;
    wire \b2v_inst36.count_rst_11_cascade_ ;
    wire \b2v_inst36.count_2_3 ;
    wire \b2v_inst36.count_rst_12_cascade_ ;
    wire \b2v_inst36.countZ0Z_2_cascade_ ;
    wire \b2v_inst36.count_2_2 ;
    wire \b2v_inst36.count_rst_7_cascade_ ;
    wire \b2v_inst36.count_rst_9_cascade_ ;
    wire \b2v_inst36.count_2_5 ;
    wire \b2v_inst36.count_2_7 ;
    wire \b2v_inst36.count_rst_7 ;
    wire \b2v_inst36.countZ0Z_5_cascade_ ;
    wire \b2v_inst36.count_2_0 ;
    wire \b2v_inst36.count_rst_14 ;
    wire \b2v_inst36.un2_count_1_axb_0 ;
    wire bfn_8_3_0_;
    wire \b2v_inst36.un2_count_1_axb_1 ;
    wire \b2v_inst36.count_rst_13 ;
    wire \b2v_inst36.un2_count_1_cry_0 ;
    wire \b2v_inst36.countZ0Z_2 ;
    wire \b2v_inst36.un2_count_1_cry_1_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_1 ;
    wire \b2v_inst36.un2_count_1_axb_3 ;
    wire \b2v_inst36.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_2 ;
    wire \b2v_inst36.un2_count_1_cry_3 ;
    wire \b2v_inst36.countZ0Z_5 ;
    wire \b2v_inst36.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_4 ;
    wire \b2v_inst36.un2_count_1_cry_5 ;
    wire \b2v_inst36.un2_count_1_axb_7 ;
    wire \b2v_inst36.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_6 ;
    wire \b2v_inst36.un2_count_1_cry_7 ;
    wire bfn_8_4_0_;
    wire \b2v_inst36.un2_count_1_cry_8 ;
    wire \b2v_inst36.un2_count_1_cry_9 ;
    wire \b2v_inst36.countZ0Z_11 ;
    wire \b2v_inst36.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_10 ;
    wire \b2v_inst36.un2_count_1_cry_11 ;
    wire \b2v_inst36.countZ0Z_13 ;
    wire \b2v_inst36.count_rst_1 ;
    wire \b2v_inst36.un2_count_1_cry_12 ;
    wire \b2v_inst36.countZ0Z_14 ;
    wire \b2v_inst36.count_rst_0 ;
    wire \b2v_inst36.un2_count_1_cry_13 ;
    wire \b2v_inst36.countZ0Z_15 ;
    wire \b2v_inst36.un2_count_1_cry_14 ;
    wire \b2v_inst36.count_rst ;
    wire \b2v_inst20.counter_1_cry_1_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_2 ;
    wire \b2v_inst36.curr_state_RNI3E27Z0Z_0_cascade_ ;
    wire dsw_pwrok;
    wire b2v_inst20_un4_counter_7_THRU_CO;
    wire \b2v_inst20.counter_1_cry_2_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_3 ;
    wire \b2v_inst5.countZ0Z_13_cascade_ ;
    wire \b2v_inst5.count_1_13 ;
    wire \b2v_inst5.count_i_0_cascade_ ;
    wire \b2v_inst5.count_rst_14 ;
    wire \b2v_inst5.count_1_0 ;
    wire \b2v_inst5.count_rst_14_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_0 ;
    wire \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2 ;
    wire \b2v_inst5.count_1_14 ;
    wire \b2v_inst5.countZ0Z_14 ;
    wire \b2v_inst5.count_i_0 ;
    wire \b2v_inst5.countZ0Z_14_cascade_ ;
    wire \b2v_inst5.countZ0Z_12 ;
    wire \b2v_inst5.count_rst_6 ;
    wire \b2v_inst5.count_rst_6_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_8 ;
    wire \b2v_inst5.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst5.un2_count_1_axb_8_cascade_ ;
    wire \b2v_inst5.count_1_8 ;
    wire \b2v_inst5.count_rst_10_cascade_ ;
    wire \b2v_inst5.countZ0Z_4 ;
    wire \b2v_inst5.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst5.countZ0Z_4_cascade_ ;
    wire \b2v_inst5.count_1_4 ;
    wire \b2v_inst5.un2_count_1_cry_12_THRU_CO ;
    wire \b2v_inst5.count_rst_1 ;
    wire \b2v_inst11.N_396_N_cascade_ ;
    wire \b2v_inst11.N_234_N_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_9 ;
    wire \b2v_inst11.dutycycle_rst_8 ;
    wire \b2v_inst11.dutycycleZ1Z_12 ;
    wire \b2v_inst11.dutycycle_eena_9_cascade_ ;
    wire \b2v_inst11.N_234_N ;
    wire \b2v_inst11.dutycycle_eena_7 ;
    wire \b2v_inst11.dutycycleZ1Z_11 ;
    wire \b2v_inst11.dutycycle_eena_7_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUFZ0Z1 ;
    wire \b2v_inst11.dutycycle_RNIT35D7Z0Z_13 ;
    wire \b2v_inst11.dutycycleZ0Z_11 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_11 ;
    wire \b2v_inst11.dutycycleZ0Z_7 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_5 ;
    wire \b2v_inst11.dutycycleZ0Z_6 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_11 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_9 ;
    wire \b2v_inst11.N_365_cascade_ ;
    wire \b2v_inst11.N_366_cascade_ ;
    wire \b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1 ;
    wire \b2v_inst11.dutycycleZ0Z_8 ;
    wire \b2v_inst11.N_153_N ;
    wire \b2v_inst11.g2_i_a6_0 ;
    wire \b2v_inst11.N_363 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ;
    wire \b2v_inst11.func_state_RNIDUQ02Z0Z_1_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0 ;
    wire \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf0_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf1 ;
    wire \b2v_inst11.N_14_0_cascade_ ;
    wire \b2v_inst11.g2_i_2 ;
    wire \b2v_inst11.func_state_RNI_6Z0Z_0 ;
    wire \b2v_inst11.N_395_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_ ;
    wire \b2v_inst11.g0_4_2 ;
    wire \b2v_inst11.g0_0_0 ;
    wire \b2v_inst11.un1_clk_100khz_36_and_i_o3_0_c_0 ;
    wire \b2v_inst11.g0_0_0_1 ;
    wire \b2v_inst11.func_state_RNI8H551Z0Z_0 ;
    wire \b2v_inst11.func_state_RNIDUQ02Z0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_7 ;
    wire \b2v_inst11.dutycycle_eena_5_d_1_1_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_5_0_1_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_36_and_i_0 ;
    wire \b2v_inst11.dutycycle_RNI2IQ6CZ0Z_7 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ;
    wire \b2v_inst11.count_clk_en_0 ;
    wire \b2v_inst11.N_328_cascade_ ;
    wire \b2v_inst11.count_clk_RNI_0Z0Z_0 ;
    wire \b2v_inst11.count_clk_en_cascade_ ;
    wire \b2v_inst11.N_218 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_329_N_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_0 ;
    wire \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7_cascade_ ;
    wire \b2v_inst11.count_clk_0_2 ;
    wire \b2v_inst11.count_clk_0_3 ;
    wire \b2v_inst11.count_clk_0_4 ;
    wire \b2v_inst11.count_clk_0_6 ;
    wire bfn_8_15_0_;
    wire \b2v_inst11.count_clkZ0Z_2 ;
    wire \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_1 ;
    wire \b2v_inst11.count_clkZ0Z_3 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2 ;
    wire \b2v_inst11.count_clkZ0Z_4 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3 ;
    wire \b2v_inst11.count_clkZ0Z_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4 ;
    wire \b2v_inst11.count_clkZ0Z_6 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6 ;
    wire \b2v_inst11.count_clkZ0Z_8 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8_cZ0 ;
    wire \b2v_inst11.count_clkZ0Z_9 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ;
    wire bfn_8_16_0_;
    wire \b2v_inst11.un1_count_clk_2_cry_9_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_10 ;
    wire \b2v_inst11.un1_count_clk_2_cry_11 ;
    wire \b2v_inst11.un1_count_clk_2_cry_12 ;
    wire \b2v_inst11.count_clkZ0Z_14 ;
    wire \b2v_inst11.count_clk_1_14 ;
    wire \b2v_inst11.un1_count_clk_2_cry_13 ;
    wire \b2v_inst11.count_clkZ0Z_15 ;
    wire \b2v_inst11.un1_count_clk_2_cry_14 ;
    wire \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ;
    wire \b2v_inst11.count_clk_0_11 ;
    wire \b2v_inst11.count_clk_1_11 ;
    wire \b2v_inst36.curr_state_7_0_cascade_ ;
    wire \b2v_inst36.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst36.curr_state_0_0 ;
    wire \b2v_inst36.curr_state_0_1 ;
    wire \b2v_inst36.curr_state_7_1 ;
    wire \b2v_inst36.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst36.DSW_PWROK_0 ;
    wire \b2v_inst36.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst36.count_2_8 ;
    wire \b2v_inst36.count_rst_6 ;
    wire \b2v_inst36.countZ0Z_8 ;
    wire \b2v_inst36.countZ0Z_8_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_5 ;
    wire \b2v_inst36.un12_clk_100khz_4 ;
    wire \b2v_inst36.un12_clk_100khz_6_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_7 ;
    wire \b2v_inst36.un12_clk_100khz_9 ;
    wire \b2v_inst36.un12_clk_100khz_13_cascade_ ;
    wire \b2v_inst36.N_1_i_cascade_ ;
    wire \b2v_inst36.count_rst_4 ;
    wire \b2v_inst36.count_rst_4_cascade_ ;
    wire \b2v_inst36.un2_count_1_axb_10 ;
    wire \b2v_inst36.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst36.un2_count_1_axb_10_cascade_ ;
    wire \b2v_inst36.N_1_i ;
    wire \b2v_inst36.count_2_10 ;
    wire \b2v_inst36.un2_count_1_axb_6 ;
    wire \b2v_inst36.count_rst_10 ;
    wire \b2v_inst36.count_2_4 ;
    wire \b2v_inst36.countZ0Z_4 ;
    wire \b2v_inst36.count_rst_8 ;
    wire \b2v_inst36.countZ0Z_4_cascade_ ;
    wire \b2v_inst36.count_2_6 ;
    wire \b2v_inst36.un12_clk_100khz_0 ;
    wire \b2v_inst36.un2_count_1_axb_12 ;
    wire \b2v_inst36.count_2_12 ;
    wire \b2v_inst36.count_rst_2 ;
    wire \b2v_inst36.un12_clk_100khz_1 ;
    wire \b2v_inst5.count_rst_13 ;
    wire \b2v_inst5.count_1_1 ;
    wire \b2v_inst5.count_rst_12 ;
    wire \b2v_inst5.count_1_2 ;
    wire \b2v_inst5.count_rst_11 ;
    wire \b2v_inst5.count_1_3 ;
    wire \b2v_inst5.countZ0Z_3 ;
    wire \b2v_inst5.countZ0Z_13 ;
    wire \b2v_inst5.countZ0Z_1 ;
    wire \b2v_inst5.countZ0Z_3_cascade_ ;
    wire \b2v_inst5.countZ0Z_2 ;
    wire \b2v_inst5.un12_clk_100khz_11 ;
    wire \b2v_inst5.un12_clk_100khz_4 ;
    wire \b2v_inst5.un12_clk_100khz_5_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_10_cascade_ ;
    wire \b2v_inst5.count_1_10 ;
    wire \b2v_inst5.un12_clk_100khz_1 ;
    wire \b2v_inst5.countZ0Z_5 ;
    wire \b2v_inst5.un12_clk_100khz_9 ;
    wire \b2v_inst5.countZ0Z_6 ;
    wire \b2v_inst5.un12_clk_100khz_12 ;
    wire \b2v_inst5.countZ0Z_9_cascade_ ;
    wire \b2v_inst5.count_1_9 ;
    wire \b2v_inst5.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst5.un2_count_1_axb_10 ;
    wire \b2v_inst5.count_rst_4 ;
    wire \b2v_inst5.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst5.curr_state_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_ ;
    wire \b2v_inst5.countZ0Z_15 ;
    wire \b2v_inst5.count_rst ;
    wire \b2v_inst5.count_1_15 ;
    wire \b2v_inst5.curr_stateZ0Z_1 ;
    wire \b2v_inst5.countZ0Z_9 ;
    wire \b2v_inst5.un2_count_1_cry_8_THRU_CO ;
    wire \b2v_inst5.N_1_i ;
    wire \b2v_inst5.count_rst_5 ;
    wire \b2v_inst5.count_rst_9 ;
    wire \b2v_inst5.count_1_5 ;
    wire \b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ;
    wire \b2v_inst5.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst5.m4_0 ;
    wire \b2v_inst5.N_2898_i_cascade_ ;
    wire N_413;
    wire \b2v_inst5.curr_state_0_0 ;
    wire \b2v_inst5.curr_stateZ0Z_0 ;
    wire \b2v_inst5.curr_state_RNIZ0Z_1 ;
    wire \b2v_inst5.N_2898_i ;
    wire \b2v_inst5.count_0_sqmuxa ;
    wire \b2v_inst11.N_172_i ;
    wire \b2v_inst11.un1_clk_100khz_2_i_o3_out ;
    wire \b2v_inst11.N_19_cascade_ ;
    wire rsmrstn_cascade_;
    wire SYNTHESIZED_WIRE_1keep_3_fast;
    wire \b2v_inst11.N_168_cascade_ ;
    wire curr_state_RNID8DP1_0_0;
    wire RSMRSTn_0;
    wire \b2v_inst11.count_clk_RNIDQ4A1Z0Z_6_cascade_ ;
    wire \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0 ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_ ;
    wire \b2v_inst11.N_186_i_cascade_ ;
    wire \b2v_inst11.N_115_f0_cascade_ ;
    wire \b2v_inst11.N_381 ;
    wire \b2v_inst11.g0_i_a7_1_2 ;
    wire \b2v_inst16.curr_state_RNIUCAD1Z0Z_0 ;
    wire \b2v_inst16.curr_stateZ0Z_1 ;
    wire \b2v_inst16.N_268 ;
    wire \b2v_inst11.N_395 ;
    wire \b2v_inst11.N_159 ;
    wire \b2v_inst11.N_159_cascade_ ;
    wire \b2v_inst11.N_425 ;
    wire \b2v_inst11.g2 ;
    wire \b2v_inst11.N_366 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_0_cascade_ ;
    wire \b2v_inst11.N_406_cascade_ ;
    wire \b2v_inst11.func_stateZ1Z_0 ;
    wire \b2v_inst11.func_state_enZ0_cascade_ ;
    wire \b2v_inst11.func_state_cascade_ ;
    wire \b2v_inst11.N_428 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0_cascade_ ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_0 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ;
    wire \b2v_inst11.N_369 ;
    wire \b2v_inst11.func_state_1_m2_ns_1_1_0_cascade_ ;
    wire \b2v_inst11.func_state_1_m2_ns_1_0_cascade_ ;
    wire \b2v_inst11.func_state_1_m2_0 ;
    wire \b2v_inst11.N_327 ;
    wire \b2v_inst11.func_state_1_m2_ns_1_1_1 ;
    wire \b2v_inst11.N_382_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_2 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_0 ;
    wire \b2v_inst11.un1_func_state25_6_0_a3_1 ;
    wire \b2v_inst11.N_406 ;
    wire \b2v_inst11.func_state_1_m2_ns_1_1 ;
    wire \b2v_inst11.func_state_1_m2_1_cascade_ ;
    wire \b2v_inst11.func_stateZ0Z_0_cascade_ ;
    wire \b2v_inst11.N_337 ;
    wire \b2v_inst11.N_338_cascade_ ;
    wire \b2v_inst11.N_76 ;
    wire \b2v_inst11.func_state_enZ0 ;
    wire \b2v_inst11.func_state_1_m2_1 ;
    wire \b2v_inst11.func_stateZ0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_5 ;
    wire \b2v_inst11.func_state_1_m2s2_i_0 ;
    wire \b2v_inst11.count_clkZ0Z_1 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_0 ;
    wire \b2v_inst11.count_clkZ0Z_0 ;
    wire \b2v_inst11.func_state_RNINIV94_0_0 ;
    wire \b2v_inst11.count_clk_0_0 ;
    wire \b2v_inst11.count_clkZ0Z_7 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ;
    wire \b2v_inst11.count_clk_0_7 ;
    wire \b2v_inst11.count_clk_0_10 ;
    wire \b2v_inst11.count_clk_1_10 ;
    wire \b2v_inst11.count_clkZ0Z_13 ;
    wire \b2v_inst11.count_clkZ0Z_11 ;
    wire \b2v_inst11.count_clkZ0Z_13_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_10 ;
    wire \b2v_inst11.un2_count_clk_17_0_o2_4 ;
    wire \b2v_inst11.count_clk_1_12 ;
    wire \b2v_inst11.count_clk_0_12 ;
    wire \b2v_inst11.count_clkZ0Z_12 ;
    wire \b2v_inst11.count_clk_1_13 ;
    wire \b2v_inst11.count_clk_0_13 ;
    wire \b2v_inst11.count_clk_en ;
    wire bfn_11_1_0_;
    wire \b2v_inst6.un2_count_1_cry_1 ;
    wire \b2v_inst6.un2_count_1_cry_2 ;
    wire \b2v_inst6.un2_count_1_cry_3 ;
    wire \b2v_inst6.un2_count_1_cry_4 ;
    wire \b2v_inst6.un2_count_1_cry_5 ;
    wire \b2v_inst6.un2_count_1_cry_6 ;
    wire \b2v_inst6.un2_count_1_cry_7 ;
    wire \b2v_inst6.un2_count_1_cry_8 ;
    wire bfn_11_2_0_;
    wire \b2v_inst6.un2_count_1_cry_9 ;
    wire \b2v_inst6.un2_count_1_cry_10 ;
    wire \b2v_inst6.un2_count_1_cry_11 ;
    wire \b2v_inst6.un2_count_1_cry_12 ;
    wire \b2v_inst6.un2_count_1_cry_13 ;
    wire \b2v_inst6.un2_count_1_cry_14 ;
    wire \b2v_inst6.count_0_15 ;
    wire \b2v_inst6.count_rst ;
    wire \b2v_inst6.countZ0Z_15 ;
    wire \b2v_inst6.countZ0Z_15_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_7 ;
    wire \b2v_inst6.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst6.un2_count_1_axb_7_cascade_ ;
    wire \b2v_inst6.count_rst_7 ;
    wire \b2v_inst6.count_0_7 ;
    wire \b2v_inst6.count_rst_7_cascade_ ;
    wire \b2v_inst6.count_en_cascade_ ;
    wire \b2v_inst6.countZ0Z_6 ;
    wire \b2v_inst6.countZ0Z_6_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_0_0_cascade_ ;
    wire \b2v_inst36.curr_stateZ0Z_1 ;
    wire \b2v_inst36.curr_stateZ0Z_0 ;
    wire v33dsw_ok;
    wire \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_ ;
    wire \b2v_inst36.countZ0Z_9 ;
    wire \b2v_inst36.count_rst_5 ;
    wire \b2v_inst36.count_2_9 ;
    wire \b2v_inst36.curr_state_RNINSDSZ0Z_0 ;
    wire \b2v_inst36.count_0_sqmuxa ;
    wire \b2v_inst6.count_0_10 ;
    wire \b2v_inst6.count_rst_4 ;
    wire \b2v_inst6.un2_count_1_axb_10 ;
    wire v33a_ok;
    wire vccst_cpu_ok;
    wire v1p8a_ok;
    wire v5a_ok;
    wire \b2v_inst6.count_rst_5_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_9 ;
    wire \b2v_inst6.un2_count_1_cry_8_THRU_CO ;
    wire \b2v_inst6.un2_count_1_axb_9_cascade_ ;
    wire \b2v_inst6.count_rst_6_cascade_ ;
    wire \b2v_inst6.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst6.countZ0Z_8_cascade_ ;
    wire \b2v_inst6.count_0_8 ;
    wire \b2v_inst6.curr_state_1_0 ;
    wire \b2v_inst6.curr_state_7_0_cascade_ ;
    wire \b2v_inst6.N_42 ;
    wire \b2v_inst6.curr_state_1_1 ;
    wire \b2v_inst6.N_42_cascade_ ;
    wire \b2v_inst6.curr_stateZ0Z_1 ;
    wire \b2v_inst6.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst6.N_3053_i_cascade_ ;
    wire \b2v_inst6.N_3034_i ;
    wire \b2v_inst6.N_3034_i_cascade_ ;
    wire \b2v_inst6.curr_state_RNIUP4B1Z0Z_0_cascade_ ;
    wire \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ;
    wire N_222;
    wire \b2v_inst6.curr_stateZ0Z_0 ;
    wire \b2v_inst6.N_3053_i ;
    wire \b2v_inst6.N_192 ;
    wire N_241;
    wire \b2v_inst6.N_276_0 ;
    wire \b2v_inst6.curr_state_RNIUP4B1Z0Z_0 ;
    wire \b2v_inst6.delayed_vccin_vccinaux_ok_0 ;
    wire \b2v_inst11.N_9 ;
    wire \b2v_inst11.N_172_cascade_ ;
    wire \b2v_inst11.g0_i_a7_1_3 ;
    wire \b2v_inst11.g0_i_0_cascade_ ;
    wire SYNTHESIZED_WIRE_1keep_3_rep1;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8 ;
    wire \b2v_inst11.N_295_cascade_ ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3_out ;
    wire \b2v_inst11.N_355 ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2 ;
    wire \b2v_inst11.dutycycleZ0Z_2_cascade_ ;
    wire \b2v_inst11.mult1_un152_sum_i ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_0_2 ;
    wire \b2v_inst11.N_168 ;
    wire \b2v_inst11.dutycycle_RNIAEUL3Z0Z_2 ;
    wire \b2v_inst11.dutycycleZ1Z_2 ;
    wire \b2v_inst11.dutycycleZ1Z_6 ;
    wire \b2v_inst11.N_365 ;
    wire \b2v_inst11.func_state_RNI_2Z0Z_1 ;
    wire \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_ ;
    wire \b2v_inst11.N_186_i ;
    wire \b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2 ;
    wire \b2v_inst11.func_state_1_ss0_i_0_o3_0_cascade_ ;
    wire \b2v_inst11.N_430 ;
    wire SYNTHESIZED_WIRE_1keep_3;
    wire \b2v_inst11.N_161 ;
    wire \b2v_inst11.N_339 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ;
    wire \b2v_inst11.dutycycle_1_0_1_cascade_ ;
    wire \b2v_inst11.dutycycle_eena ;
    wire \b2v_inst11.dutycycleZ1Z_0 ;
    wire \b2v_inst11.dutycycle_eena_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_0 ;
    wire \b2v_inst11.dutycycleZ0Z_0_cascade_ ;
    wire \b2v_inst11.dutycycle_1_0_0 ;
    wire \b2v_inst11.N_119_f0_1 ;
    wire \b2v_inst11.dutycycle ;
    wire \b2v_inst11.dutycycle_eena_0 ;
    wire G_146;
    wire \b2v_inst11.dutycycle_1_0_1 ;
    wire \b2v_inst11.dutycycle_eena_0_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_1 ;
    wire \b2v_inst11.N_224_iZ0 ;
    wire \b2v_inst11.count_off_1_0_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_330_N ;
    wire \b2v_inst11.func_state ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_0 ;
    wire \b2v_inst11.N_382 ;
    wire \b2v_inst11.count_clk_RNI_0Z0Z_1 ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ;
    wire \b2v_inst11.N_315_cascade_ ;
    wire \b2v_inst11.count_clk_RNIDQ4A1Z0Z_7 ;
    wire \b2v_inst11.N_125_cascade_ ;
    wire \b2v_inst11.N_382_N ;
    wire bfn_11_13_0_;
    wire \b2v_inst11.un3_count_off_1_cry_1 ;
    wire \b2v_inst11.un3_count_off_1_cry_2 ;
    wire \b2v_inst11.un3_count_off_1_cry_3 ;
    wire \b2v_inst11.un3_count_off_1_cry_4 ;
    wire \b2v_inst11.un3_count_off_1_cry_5 ;
    wire \b2v_inst11.un3_count_off_1_cry_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_7 ;
    wire \b2v_inst11.un3_count_off_1_cry_8 ;
    wire bfn_11_14_0_;
    wire \b2v_inst11.un3_count_off_1_cry_9 ;
    wire \b2v_inst11.un3_count_off_1_cry_10 ;
    wire \b2v_inst11.un3_count_off_1_cry_11 ;
    wire \b2v_inst11.un3_count_off_1_cry_12 ;
    wire \b2v_inst11.un3_count_off_1_cry_13 ;
    wire \b2v_inst11.un3_count_off_1_cry_14 ;
    wire \b2v_inst11.count_off_1_14 ;
    wire \b2v_inst11.count_off_0_14 ;
    wire \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DTZ0Z63 ;
    wire \b2v_inst11.count_off_0_15 ;
    wire \b2v_inst11.count_off_1_6 ;
    wire \b2v_inst11.count_off_0_6 ;
    wire \b2v_inst11.count_off_1_7 ;
    wire \b2v_inst11.count_off_0_7 ;
    wire \b2v_inst11.count_off_1_8 ;
    wire \b2v_inst11.count_off_0_8 ;
    wire \b2v_inst6.count_rst_10_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_4 ;
    wire \b2v_inst6.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst6.un2_count_1_axb_4_cascade_ ;
    wire \b2v_inst6.count_rst_10 ;
    wire \b2v_inst6.count_0_4 ;
    wire \b2v_inst6.count_rst_11_cascade_ ;
    wire \b2v_inst6.countZ0Z_3 ;
    wire \b2v_inst6.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst6.countZ0Z_3_cascade_ ;
    wire \b2v_inst6.count_0_3 ;
    wire \b2v_inst6.un2_count_1_axb_2 ;
    wire \b2v_inst6.count_0_14 ;
    wire \b2v_inst6.un2_count_1_cry_13_c_RNI06SPZ0Z1 ;
    wire \b2v_inst6.countZ0Z_14 ;
    wire \b2v_inst6.count_0_2 ;
    wire \b2v_inst6.countZ0Z_14_cascade_ ;
    wire \b2v_inst6.count_rst_12 ;
    wire \b2v_inst6.un2_count_1_axb_12 ;
    wire \b2v_inst6.count_rst_2 ;
    wire \b2v_inst6.count_0_12 ;
    wire \b2v_inst6.count_rst_1 ;
    wire \b2v_inst6.count_0_13 ;
    wire \b2v_inst6.un2_count_1_axb_13 ;
    wire \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ;
    wire \b2v_inst6.count_0_6 ;
    wire \b2v_inst6.N_394_cascade_ ;
    wire \b2v_inst6.count_rst_9_cascade_ ;
    wire \b2v_inst6.countZ0Z_5 ;
    wire \b2v_inst6.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst6.countZ0Z_5_cascade_ ;
    wire \b2v_inst6.count_0_5 ;
    wire \b2v_inst6.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst6.N_394 ;
    wire \b2v_inst6.count_rst_3_cascade_ ;
    wire \b2v_inst6.count_0_11 ;
    wire \b2v_inst6.count_RNIM6FE1Z0Z_0 ;
    wire \b2v_inst6.countZ0Z_0_cascade_ ;
    wire \b2v_inst6.countZ0Z_11 ;
    wire \b2v_inst6.count_rst_13_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_5_0 ;
    wire \b2v_inst6.count_1_i_a3_6_0 ;
    wire \b2v_inst6.count_1_i_a3_3_0_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_7_0 ;
    wire \b2v_inst6.count_1_i_a3_1_0 ;
    wire \b2v_inst6.count_1_i_a3_12_0_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_2_0 ;
    wire \b2v_inst6.N_389 ;
    wire \b2v_inst6.N_389_cascade_ ;
    wire \b2v_inst6.count_0_0 ;
    wire \b2v_inst6.count_rst_13 ;
    wire \b2v_inst6.un2_count_1_axb_1 ;
    wire \b2v_inst6.un2_count_1_axb_1_cascade_ ;
    wire \b2v_inst6.count_0_1 ;
    wire \b2v_inst6.curr_state_RNIM6FE1Z0Z_1 ;
    wire \b2v_inst6.count_rst_5 ;
    wire \b2v_inst6.count_0_9 ;
    wire \b2v_inst6.countZ0Z_8 ;
    wire \b2v_inst6.count_en ;
    wire \b2v_inst6.count_1_i_a3_4_0 ;
    wire \b2v_inst5.N_51 ;
    wire \b2v_inst5.curr_state_0_1 ;
    wire N_606_g;
    wire \b2v_inst6.countZ0Z_0 ;
    wire \b2v_inst6.N_3036_i ;
    wire CONSTANT_ONE_NET;
    wire v5s_ok;
    wire v33s_ok;
    wire SYNTHESIZED_WIRE_8;
    wire vccinaux_en;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_0 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_0_cascade_ ;
    wire slp_s4n;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_0 ;
    wire \b2v_inst11.un1_dutycycle_172_m1_ns_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_172_m1 ;
    wire \b2v_inst11.g0_i_2 ;
    wire \b2v_inst11.g0_0_0Z0Z_0_cascade_ ;
    wire \b2v_inst11.g0_13_1_cascade_ ;
    wire \b2v_inst11.N_4690_0_0_cascade_ ;
    wire \b2v_inst11.N_19_0 ;
    wire \b2v_inst11.N_19_1 ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ;
    wire \b2v_inst11.un1_dutycycle_172_m0 ;
    wire \b2v_inst11.g3_3 ;
    wire \b2v_inst11.N_172 ;
    wire \b2v_inst11.N_200_i ;
    wire \b2v_inst11.N_3099_0_0 ;
    wire \b2v_inst11.dutycycleZ0Z_2 ;
    wire \b2v_inst11.N_237 ;
    wire \b2v_inst11.N_293_0_0 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_6 ;
    wire \b2v_inst11.g2_1_0 ;
    wire \b2v_inst11.dutycycleZ0Z_5 ;
    wire \b2v_inst11.func_stateZ0Z_0 ;
    wire G_6_i_a3_1;
    wire N_5_cascade_;
    wire v5s_enn;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_rn_1 ;
    wire b2v_inst11_un1_clk_100khz_52_and_i_0_cascade_;
    wire \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_sn ;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_0_cascade_ ;
    wire \b2v_inst11.N_6063_0_0 ;
    wire \b2v_inst11.dutycycle_eena_14_0_0 ;
    wire slp_s3n;
    wire gpio_fpga_soc_4;
    wire rsmrstn;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0 ;
    wire \b2v_inst11.N_2946_i ;
    wire \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_5 ;
    wire \b2v_inst11.g0_1_1 ;
    wire vddq_ok;
    wire VCCST_EN_i_0_o3_0;
    wire \b2v_inst16.N_208_0 ;
    wire \b2v_inst11.count_off_1_1 ;
    wire \b2v_inst11.count_offZ0Z_6 ;
    wire \b2v_inst11.count_offZ0Z_5 ;
    wire \b2v_inst11.count_offZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_offZ0Z_2 ;
    wire \b2v_inst11.un34_clk_100khz_9_cascade_ ;
    wire \b2v_inst11.count_off_RNI_0Z0Z_1 ;
    wire \b2v_inst11.count_offZ0Z_15 ;
    wire \b2v_inst11.count_offZ0Z_13 ;
    wire \b2v_inst11.count_offZ0Z_14 ;
    wire \b2v_inst11.un34_clk_100khz_10 ;
    wire \b2v_inst11.count_offZ0Z_7 ;
    wire \b2v_inst11.count_offZ0Z_8 ;
    wire \b2v_inst11.count_offZ0Z_3 ;
    wire \b2v_inst11.count_offZ0Z_4 ;
    wire \b2v_inst11.un34_clk_100khz_8 ;
    wire \b2v_inst11.count_offZ0Z_1 ;
    wire \b2v_inst11.count_off_0_1 ;
    wire \b2v_inst11.count_offZ0Z_0 ;
    wire \b2v_inst11.N_125 ;
    wire \b2v_inst11.count_off_0_0 ;
    wire \b2v_inst11.count_off_0_9 ;
    wire \b2v_inst11.count_off_1_9 ;
    wire \b2v_inst11.count_offZ0Z_9 ;
    wire \b2v_inst11.count_offZ0Z_9_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_11 ;
    wire \b2v_inst11.count_offZ0Z_10 ;
    wire \b2v_inst11.count_off_1_10 ;
    wire \b2v_inst11.count_off_0_10 ;
    wire \b2v_inst11.count_offZ0Z_11 ;
    wire \b2v_inst11.count_off_1_11 ;
    wire \b2v_inst11.count_off_0_11 ;
    wire \b2v_inst11.count_offZ0Z_12 ;
    wire \b2v_inst11.count_off_1_12 ;
    wire \b2v_inst11.count_off_0_12 ;
    wire \b2v_inst11.count_off_1_13 ;
    wire \b2v_inst11.count_off_0_13 ;
    wire \b2v_inst11.count_off_1_2 ;
    wire \b2v_inst11.count_off_0_2 ;
    wire \b2v_inst11.count_off_1_3 ;
    wire \b2v_inst11.count_off_0_3 ;
    wire \b2v_inst11.count_off_1_4 ;
    wire \b2v_inst11.count_off_0_4 ;
    wire \b2v_inst11.count_off_1_5 ;
    wire \b2v_inst11.count_off_0_5 ;
    wire fpga_osc;
    wire \b2v_inst11.dutycycle_RNIHJNV7Z0Z_0 ;
    wire _gnd_net_;

    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__37287),
            .DIN(N__37286),
            .DOUT(N__37285),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__37287),
            .PADOUT(N__37286),
            .PADIN(N__37285),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccinaux),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__37278),
            .DIN(N__37277),
            .DOUT(N__37276),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__37278),
            .PADOUT(N__37277),
            .PADIN(N__37276),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__37269),
            .DIN(N__37268),
            .DOUT(N__37267),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__37269),
            .PADOUT(N__37268),
            .PADIN(N__37267),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__37260),
            .DIN(N__37259),
            .DOUT(N__37258),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__37260),
            .PADOUT(N__37259),
            .PADIN(N__37258),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18191),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__37251),
            .DIN(N__37250),
            .DOUT(N__37249),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__37251),
            .PADOUT(N__37250),
            .PADIN(N__37249),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__37242),
            .DIN(N__37241),
            .DOUT(N__37240),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__37242),
            .PADOUT(N__37241),
            .PADIN(N__37240),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__37233),
            .DIN(N__37232),
            .DOUT(N__37231),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__37233),
            .PADOUT(N__37232),
            .PADIN(N__37231),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__37224),
            .DIN(N__37223),
            .DOUT(N__37222),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__37224),
            .PADOUT(N__37223),
            .PADIN(N__37222),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__37215),
            .DIN(N__37214),
            .DOUT(N__37213),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__37215),
            .PADOUT(N__37214),
            .PADIN(N__37213),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34945),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__37206),
            .DIN(N__37205),
            .DOUT(N__37204),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__37206),
            .PADOUT(N__37205),
            .PADIN(N__37204),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__37197),
            .DIN(N__37196),
            .DOUT(N__37195),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__37197),
            .PADOUT(N__37196),
            .PADIN(N__37195),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__37188),
            .DIN(N__37187),
            .DOUT(N__37186),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__37188),
            .PADOUT(N__37187),
            .PADIN(N__37186),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17168),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__37179),
            .DIN(N__37178),
            .DOUT(N__37177),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__37179),
            .PADOUT(N__37178),
            .PADIN(N__37177),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__37170),
            .DIN(N__37169),
            .DOUT(N__37168),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__37170),
            .PADOUT(N__37169),
            .PADIN(N__37168),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__37161),
            .DIN(N__37160),
            .DOUT(N__37159),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__37161),
            .PADOUT(N__37160),
            .PADIN(N__37159),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__37152),
            .DIN(N__37151),
            .DOUT(N__37150),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__37152),
            .PADOUT(N__37151),
            .PADIN(N__37150),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__37143),
            .DIN(N__37142),
            .DOUT(N__37141),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__37143),
            .PADOUT(N__37142),
            .PADIN(N__37141),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19916),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__37134),
            .DIN(N__37133),
            .DOUT(N__37132),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__37134),
            .PADOUT(N__37133),
            .PADIN(N__37132),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33dsw_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__37125),
            .DIN(N__37124),
            .DOUT(N__37123),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__37125),
            .PADOUT(N__37124),
            .PADIN(N__37123),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__37116),
            .DIN(N__37115),
            .DOUT(N__37114),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__37116),
            .PADOUT(N__37115),
            .PADIN(N__37114),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__37107),
            .DIN(N__37106),
            .DOUT(N__37105),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__37107),
            .PADOUT(N__37106),
            .PADIN(N__37105),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__37098),
            .DIN(N__37097),
            .DOUT(N__37096),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__37098),
            .PADOUT(N__37097),
            .PADIN(N__37096),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__37089),
            .DIN(N__37088),
            .DOUT(N__37087),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__37089),
            .PADOUT(N__37088),
            .PADIN(N__37087),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__37080),
            .DIN(N__37079),
            .DOUT(N__37078),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__37080),
            .PADOUT(N__37079),
            .PADIN(N__37078),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__37071),
            .DIN(N__37070),
            .DOUT(N__37069),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__37071),
            .PADOUT(N__37070),
            .PADIN(N__37069),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34319),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__37062),
            .DIN(N__37061),
            .DOUT(N__37060),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__37062),
            .PADOUT(N__37061),
            .PADIN(N__37060),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__37053),
            .DIN(N__37052),
            .DOUT(N__37051),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__37053),
            .PADOUT(N__37052),
            .PADIN(N__37051),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17344),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__37044),
            .DIN(N__37043),
            .DOUT(N__37042),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__37044),
            .PADOUT(N__37043),
            .PADIN(N__37042),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17354),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__37035),
            .DIN(N__37034),
            .DOUT(N__37033),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__37035),
            .PADOUT(N__37034),
            .PADIN(N__37033),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__37026),
            .DIN(N__37025),
            .DOUT(N__37024),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__37026),
            .PADOUT(N__37025),
            .PADIN(N__37024),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__37017),
            .DIN(N__37016),
            .DOUT(N__37015),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__37017),
            .PADOUT(N__37016),
            .PADIN(N__37015),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__37008),
            .DIN(N__37007),
            .DOUT(N__37006),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__37008),
            .PADOUT(N__37007),
            .PADIN(N__37006),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__36999),
            .DIN(N__36998),
            .DOUT(N__36997),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__36999),
            .PADOUT(N__36998),
            .PADIN(N__36997),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__36990),
            .DIN(N__36989),
            .DOUT(N__36988),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__36990),
            .PADOUT(N__36989),
            .PADIN(N__36988),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19379),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__36981),
            .DIN(N__36980),
            .DOUT(N__36979),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__36981),
            .PADOUT(N__36980),
            .PADIN(N__36979),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__36972),
            .DIN(N__36971),
            .DOUT(N__36970),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__36972),
            .PADOUT(N__36971),
            .PADIN(N__36970),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17771),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__36963),
            .DIN(N__36962),
            .DOUT(N__36961),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__36963),
            .PADOUT(N__36962),
            .PADIN(N__36961),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__36954),
            .DIN(N__36953),
            .DOUT(N__36952),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__36954),
            .PADOUT(N__36953),
            .PADIN(N__36952),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__36945),
            .DIN(N__36944),
            .DOUT(N__36943),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__36945),
            .PADOUT(N__36944),
            .PADIN(N__36943),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__36936),
            .DIN(N__36935),
            .DOUT(N__36934),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__36936),
            .PADOUT(N__36935),
            .PADIN(N__36934),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__36927),
            .DIN(N__36926),
            .DOUT(N__36925),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__36927),
            .PADOUT(N__36926),
            .PADIN(N__36925),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32938),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__36918),
            .DIN(N__36917),
            .DOUT(N__36916),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__36918),
            .PADOUT(N__36917),
            .PADIN(N__36916),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__36909),
            .DIN(N__36908),
            .DOUT(N__36907),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__36909),
            .PADOUT(N__36908),
            .PADIN(N__36907),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34946),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__36900),
            .DIN(N__36899),
            .DOUT(N__36898),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__36900),
            .PADOUT(N__36899),
            .PADIN(N__36898),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__36891),
            .DIN(N__36890),
            .DOUT(N__36889),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__36891),
            .PADOUT(N__36890),
            .PADIN(N__36889),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24212),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__36882),
            .DIN(N__36881),
            .DOUT(N__36880),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__36882),
            .PADOUT(N__36881),
            .PADIN(N__36880),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32060),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__36873),
            .DIN(N__36872),
            .DOUT(N__36871),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__36873),
            .PADOUT(N__36872),
            .PADIN(N__36871),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__36864),
            .DIN(N__36863),
            .DOUT(N__36862),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__36864),
            .PADOUT(N__36863),
            .PADIN(N__36862),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__36855),
            .DIN(N__36854),
            .DOUT(N__36853),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__36855),
            .PADOUT(N__36854),
            .PADIN(N__36853),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__36846),
            .DIN(N__36845),
            .DOUT(N__36844),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__36846),
            .PADOUT(N__36845),
            .PADIN(N__36844),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__36837),
            .DIN(N__36836),
            .DOUT(N__36835),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__36837),
            .PADOUT(N__36836),
            .PADIN(N__36835),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32951),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__36828),
            .DIN(N__36827),
            .DOUT(N__36826),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__36828),
            .PADOUT(N__36827),
            .PADIN(N__36826),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__36819),
            .DIN(N__36818),
            .DOUT(N__36817),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__36819),
            .PADOUT(N__36818),
            .PADIN(N__36817),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__36810),
            .DIN(N__36809),
            .DOUT(N__36808),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__36810),
            .PADOUT(N__36809),
            .PADIN(N__36808),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__36801),
            .DIN(N__36800),
            .DOUT(N__36799),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__36801),
            .PADOUT(N__36800),
            .PADIN(N__36799),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__36792),
            .DIN(N__36791),
            .DOUT(N__36790),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__36792),
            .PADOUT(N__36791),
            .PADIN(N__36790),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__36783),
            .DIN(N__36782),
            .DOUT(N__36781),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__36783),
            .PADOUT(N__36782),
            .PADIN(N__36781),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__36774),
            .DIN(N__36773),
            .DOUT(N__36772),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__36774),
            .PADOUT(N__36773),
            .PADIN(N__36772),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17337),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__36765),
            .DIN(N__36764),
            .DOUT(N__36763),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__36765),
            .PADOUT(N__36764),
            .PADIN(N__36763),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__8563 (
            .O(N__36746),
            .I(N__36743));
    LocalMux I__8562 (
            .O(N__36743),
            .I(N__36739));
    InMux I__8561 (
            .O(N__36742),
            .I(N__36736));
    Span4Mux_h I__8560 (
            .O(N__36739),
            .I(N__36733));
    LocalMux I__8559 (
            .O(N__36736),
            .I(\b2v_inst11.count_off_1_3 ));
    Odrv4 I__8558 (
            .O(N__36733),
            .I(\b2v_inst11.count_off_1_3 ));
    InMux I__8557 (
            .O(N__36728),
            .I(N__36725));
    LocalMux I__8556 (
            .O(N__36725),
            .I(N__36722));
    Odrv4 I__8555 (
            .O(N__36722),
            .I(\b2v_inst11.count_off_0_3 ));
    InMux I__8554 (
            .O(N__36719),
            .I(N__36716));
    LocalMux I__8553 (
            .O(N__36716),
            .I(N__36712));
    InMux I__8552 (
            .O(N__36715),
            .I(N__36709));
    Span4Mux_h I__8551 (
            .O(N__36712),
            .I(N__36706));
    LocalMux I__8550 (
            .O(N__36709),
            .I(\b2v_inst11.count_off_1_4 ));
    Odrv4 I__8549 (
            .O(N__36706),
            .I(\b2v_inst11.count_off_1_4 ));
    InMux I__8548 (
            .O(N__36701),
            .I(N__36698));
    LocalMux I__8547 (
            .O(N__36698),
            .I(N__36695));
    Odrv4 I__8546 (
            .O(N__36695),
            .I(\b2v_inst11.count_off_0_4 ));
    InMux I__8545 (
            .O(N__36692),
            .I(N__36689));
    LocalMux I__8544 (
            .O(N__36689),
            .I(N__36685));
    InMux I__8543 (
            .O(N__36688),
            .I(N__36682));
    Span4Mux_s3_v I__8542 (
            .O(N__36685),
            .I(N__36679));
    LocalMux I__8541 (
            .O(N__36682),
            .I(\b2v_inst11.count_off_1_5 ));
    Odrv4 I__8540 (
            .O(N__36679),
            .I(\b2v_inst11.count_off_1_5 ));
    InMux I__8539 (
            .O(N__36674),
            .I(N__36671));
    LocalMux I__8538 (
            .O(N__36671),
            .I(N__36668));
    Odrv4 I__8537 (
            .O(N__36668),
            .I(\b2v_inst11.count_off_0_5 ));
    ClkMux I__8536 (
            .O(N__36665),
            .I(N__36662));
    LocalMux I__8535 (
            .O(N__36662),
            .I(N__36658));
    ClkMux I__8534 (
            .O(N__36661),
            .I(N__36653));
    Span4Mux_s3_h I__8533 (
            .O(N__36658),
            .I(N__36649));
    ClkMux I__8532 (
            .O(N__36657),
            .I(N__36646));
    ClkMux I__8531 (
            .O(N__36656),
            .I(N__36643));
    LocalMux I__8530 (
            .O(N__36653),
            .I(N__36640));
    ClkMux I__8529 (
            .O(N__36652),
            .I(N__36637));
    Span4Mux_h I__8528 (
            .O(N__36649),
            .I(N__36628));
    LocalMux I__8527 (
            .O(N__36646),
            .I(N__36628));
    LocalMux I__8526 (
            .O(N__36643),
            .I(N__36628));
    Span4Mux_v I__8525 (
            .O(N__36640),
            .I(N__36623));
    LocalMux I__8524 (
            .O(N__36637),
            .I(N__36623));
    ClkMux I__8523 (
            .O(N__36636),
            .I(N__36620));
    ClkMux I__8522 (
            .O(N__36635),
            .I(N__36615));
    Span4Mux_v I__8521 (
            .O(N__36628),
            .I(N__36608));
    Span4Mux_h I__8520 (
            .O(N__36623),
            .I(N__36608));
    LocalMux I__8519 (
            .O(N__36620),
            .I(N__36608));
    ClkMux I__8518 (
            .O(N__36619),
            .I(N__36605));
    ClkMux I__8517 (
            .O(N__36618),
            .I(N__36599));
    LocalMux I__8516 (
            .O(N__36615),
            .I(N__36593));
    Span4Mux_v I__8515 (
            .O(N__36608),
            .I(N__36593));
    LocalMux I__8514 (
            .O(N__36605),
            .I(N__36590));
    ClkMux I__8513 (
            .O(N__36604),
            .I(N__36587));
    ClkMux I__8512 (
            .O(N__36603),
            .I(N__36583));
    ClkMux I__8511 (
            .O(N__36602),
            .I(N__36576));
    LocalMux I__8510 (
            .O(N__36599),
            .I(N__36572));
    ClkMux I__8509 (
            .O(N__36598),
            .I(N__36569));
    IoSpan4Mux I__8508 (
            .O(N__36593),
            .I(N__36565));
    Span4Mux_v I__8507 (
            .O(N__36590),
            .I(N__36560));
    LocalMux I__8506 (
            .O(N__36587),
            .I(N__36560));
    ClkMux I__8505 (
            .O(N__36586),
            .I(N__36557));
    LocalMux I__8504 (
            .O(N__36583),
            .I(N__36553));
    ClkMux I__8503 (
            .O(N__36582),
            .I(N__36549));
    ClkMux I__8502 (
            .O(N__36581),
            .I(N__36546));
    ClkMux I__8501 (
            .O(N__36580),
            .I(N__36543));
    ClkMux I__8500 (
            .O(N__36579),
            .I(N__36538));
    LocalMux I__8499 (
            .O(N__36576),
            .I(N__36535));
    ClkMux I__8498 (
            .O(N__36575),
            .I(N__36532));
    Span4Mux_v I__8497 (
            .O(N__36572),
            .I(N__36527));
    LocalMux I__8496 (
            .O(N__36569),
            .I(N__36524));
    ClkMux I__8495 (
            .O(N__36568),
            .I(N__36521));
    Span4Mux_s1_h I__8494 (
            .O(N__36565),
            .I(N__36514));
    Span4Mux_h I__8493 (
            .O(N__36560),
            .I(N__36514));
    LocalMux I__8492 (
            .O(N__36557),
            .I(N__36514));
    ClkMux I__8491 (
            .O(N__36556),
            .I(N__36511));
    IoSpan4Mux I__8490 (
            .O(N__36553),
            .I(N__36507));
    ClkMux I__8489 (
            .O(N__36552),
            .I(N__36504));
    LocalMux I__8488 (
            .O(N__36549),
            .I(N__36498));
    LocalMux I__8487 (
            .O(N__36546),
            .I(N__36498));
    LocalMux I__8486 (
            .O(N__36543),
            .I(N__36495));
    ClkMux I__8485 (
            .O(N__36542),
            .I(N__36492));
    ClkMux I__8484 (
            .O(N__36541),
            .I(N__36486));
    LocalMux I__8483 (
            .O(N__36538),
            .I(N__36482));
    Span4Mux_s2_v I__8482 (
            .O(N__36535),
            .I(N__36474));
    LocalMux I__8481 (
            .O(N__36532),
            .I(N__36474));
    ClkMux I__8480 (
            .O(N__36531),
            .I(N__36471));
    ClkMux I__8479 (
            .O(N__36530),
            .I(N__36465));
    Span4Mux_v I__8478 (
            .O(N__36527),
            .I(N__36454));
    Span4Mux_s1_h I__8477 (
            .O(N__36524),
            .I(N__36454));
    LocalMux I__8476 (
            .O(N__36521),
            .I(N__36454));
    Span4Mux_h I__8475 (
            .O(N__36514),
            .I(N__36454));
    LocalMux I__8474 (
            .O(N__36511),
            .I(N__36454));
    ClkMux I__8473 (
            .O(N__36510),
            .I(N__36451));
    Span4Mux_s2_h I__8472 (
            .O(N__36507),
            .I(N__36442));
    LocalMux I__8471 (
            .O(N__36504),
            .I(N__36442));
    ClkMux I__8470 (
            .O(N__36503),
            .I(N__36439));
    Span4Mux_v I__8469 (
            .O(N__36498),
            .I(N__36429));
    Span4Mux_v I__8468 (
            .O(N__36495),
            .I(N__36429));
    LocalMux I__8467 (
            .O(N__36492),
            .I(N__36429));
    ClkMux I__8466 (
            .O(N__36491),
            .I(N__36426));
    ClkMux I__8465 (
            .O(N__36490),
            .I(N__36423));
    ClkMux I__8464 (
            .O(N__36489),
            .I(N__36417));
    LocalMux I__8463 (
            .O(N__36486),
            .I(N__36413));
    ClkMux I__8462 (
            .O(N__36485),
            .I(N__36410));
    Span4Mux_s1_h I__8461 (
            .O(N__36482),
            .I(N__36407));
    ClkMux I__8460 (
            .O(N__36481),
            .I(N__36404));
    ClkMux I__8459 (
            .O(N__36480),
            .I(N__36398));
    ClkMux I__8458 (
            .O(N__36479),
            .I(N__36395));
    Span4Mux_v I__8457 (
            .O(N__36474),
            .I(N__36389));
    LocalMux I__8456 (
            .O(N__36471),
            .I(N__36389));
    ClkMux I__8455 (
            .O(N__36470),
            .I(N__36386));
    ClkMux I__8454 (
            .O(N__36469),
            .I(N__36383));
    ClkMux I__8453 (
            .O(N__36468),
            .I(N__36380));
    LocalMux I__8452 (
            .O(N__36465),
            .I(N__36377));
    Span4Mux_v I__8451 (
            .O(N__36454),
            .I(N__36372));
    LocalMux I__8450 (
            .O(N__36451),
            .I(N__36372));
    ClkMux I__8449 (
            .O(N__36450),
            .I(N__36369));
    ClkMux I__8448 (
            .O(N__36449),
            .I(N__36364));
    ClkMux I__8447 (
            .O(N__36448),
            .I(N__36361));
    ClkMux I__8446 (
            .O(N__36447),
            .I(N__36357));
    Span4Mux_s3_v I__8445 (
            .O(N__36442),
            .I(N__36351));
    LocalMux I__8444 (
            .O(N__36439),
            .I(N__36351));
    ClkMux I__8443 (
            .O(N__36438),
            .I(N__36346));
    ClkMux I__8442 (
            .O(N__36437),
            .I(N__36343));
    ClkMux I__8441 (
            .O(N__36436),
            .I(N__36340));
    Span4Mux_v I__8440 (
            .O(N__36429),
            .I(N__36332));
    LocalMux I__8439 (
            .O(N__36426),
            .I(N__36332));
    LocalMux I__8438 (
            .O(N__36423),
            .I(N__36332));
    ClkMux I__8437 (
            .O(N__36422),
            .I(N__36329));
    ClkMux I__8436 (
            .O(N__36421),
            .I(N__36326));
    ClkMux I__8435 (
            .O(N__36420),
            .I(N__36323));
    LocalMux I__8434 (
            .O(N__36417),
            .I(N__36319));
    ClkMux I__8433 (
            .O(N__36416),
            .I(N__36316));
    Span4Mux_h I__8432 (
            .O(N__36413),
            .I(N__36309));
    LocalMux I__8431 (
            .O(N__36410),
            .I(N__36309));
    Span4Mux_h I__8430 (
            .O(N__36407),
            .I(N__36304));
    LocalMux I__8429 (
            .O(N__36404),
            .I(N__36304));
    ClkMux I__8428 (
            .O(N__36403),
            .I(N__36301));
    ClkMux I__8427 (
            .O(N__36402),
            .I(N__36298));
    ClkMux I__8426 (
            .O(N__36401),
            .I(N__36295));
    LocalMux I__8425 (
            .O(N__36398),
            .I(N__36292));
    LocalMux I__8424 (
            .O(N__36395),
            .I(N__36288));
    ClkMux I__8423 (
            .O(N__36394),
            .I(N__36285));
    Span4Mux_v I__8422 (
            .O(N__36389),
            .I(N__36280));
    LocalMux I__8421 (
            .O(N__36386),
            .I(N__36280));
    LocalMux I__8420 (
            .O(N__36383),
            .I(N__36277));
    LocalMux I__8419 (
            .O(N__36380),
            .I(N__36274));
    Span4Mux_s1_h I__8418 (
            .O(N__36377),
            .I(N__36267));
    Span4Mux_s1_v I__8417 (
            .O(N__36372),
            .I(N__36267));
    LocalMux I__8416 (
            .O(N__36369),
            .I(N__36267));
    ClkMux I__8415 (
            .O(N__36368),
            .I(N__36264));
    ClkMux I__8414 (
            .O(N__36367),
            .I(N__36260));
    LocalMux I__8413 (
            .O(N__36364),
            .I(N__36257));
    LocalMux I__8412 (
            .O(N__36361),
            .I(N__36254));
    ClkMux I__8411 (
            .O(N__36360),
            .I(N__36251));
    LocalMux I__8410 (
            .O(N__36357),
            .I(N__36248));
    ClkMux I__8409 (
            .O(N__36356),
            .I(N__36245));
    Span4Mux_v I__8408 (
            .O(N__36351),
            .I(N__36241));
    ClkMux I__8407 (
            .O(N__36350),
            .I(N__36238));
    ClkMux I__8406 (
            .O(N__36349),
            .I(N__36235));
    LocalMux I__8405 (
            .O(N__36346),
            .I(N__36231));
    LocalMux I__8404 (
            .O(N__36343),
            .I(N__36228));
    LocalMux I__8403 (
            .O(N__36340),
            .I(N__36225));
    ClkMux I__8402 (
            .O(N__36339),
            .I(N__36222));
    Span4Mux_v I__8401 (
            .O(N__36332),
            .I(N__36213));
    LocalMux I__8400 (
            .O(N__36329),
            .I(N__36213));
    LocalMux I__8399 (
            .O(N__36326),
            .I(N__36213));
    LocalMux I__8398 (
            .O(N__36323),
            .I(N__36213));
    ClkMux I__8397 (
            .O(N__36322),
            .I(N__36210));
    Span4Mux_s3_v I__8396 (
            .O(N__36319),
            .I(N__36202));
    LocalMux I__8395 (
            .O(N__36316),
            .I(N__36202));
    ClkMux I__8394 (
            .O(N__36315),
            .I(N__36199));
    ClkMux I__8393 (
            .O(N__36314),
            .I(N__36195));
    Span4Mux_v I__8392 (
            .O(N__36309),
            .I(N__36185));
    Span4Mux_v I__8391 (
            .O(N__36304),
            .I(N__36185));
    LocalMux I__8390 (
            .O(N__36301),
            .I(N__36185));
    LocalMux I__8389 (
            .O(N__36298),
            .I(N__36182));
    LocalMux I__8388 (
            .O(N__36295),
            .I(N__36179));
    Span4Mux_s1_h I__8387 (
            .O(N__36292),
            .I(N__36176));
    ClkMux I__8386 (
            .O(N__36291),
            .I(N__36173));
    Span4Mux_v I__8385 (
            .O(N__36288),
            .I(N__36168));
    LocalMux I__8384 (
            .O(N__36285),
            .I(N__36168));
    Span4Mux_v I__8383 (
            .O(N__36280),
            .I(N__36156));
    Span4Mux_s2_h I__8382 (
            .O(N__36277),
            .I(N__36156));
    Span4Mux_s2_h I__8381 (
            .O(N__36274),
            .I(N__36156));
    Span4Mux_h I__8380 (
            .O(N__36267),
            .I(N__36156));
    LocalMux I__8379 (
            .O(N__36264),
            .I(N__36156));
    ClkMux I__8378 (
            .O(N__36263),
            .I(N__36153));
    LocalMux I__8377 (
            .O(N__36260),
            .I(N__36150));
    Span4Mux_s2_h I__8376 (
            .O(N__36257),
            .I(N__36139));
    Span4Mux_h I__8375 (
            .O(N__36254),
            .I(N__36139));
    LocalMux I__8374 (
            .O(N__36251),
            .I(N__36139));
    Span4Mux_h I__8373 (
            .O(N__36248),
            .I(N__36139));
    LocalMux I__8372 (
            .O(N__36245),
            .I(N__36139));
    ClkMux I__8371 (
            .O(N__36244),
            .I(N__36136));
    Span4Mux_v I__8370 (
            .O(N__36241),
            .I(N__36131));
    LocalMux I__8369 (
            .O(N__36238),
            .I(N__36131));
    LocalMux I__8368 (
            .O(N__36235),
            .I(N__36128));
    ClkMux I__8367 (
            .O(N__36234),
            .I(N__36125));
    Span4Mux_h I__8366 (
            .O(N__36231),
            .I(N__36116));
    Span4Mux_v I__8365 (
            .O(N__36228),
            .I(N__36116));
    Span4Mux_h I__8364 (
            .O(N__36225),
            .I(N__36116));
    LocalMux I__8363 (
            .O(N__36222),
            .I(N__36116));
    IoSpan4Mux I__8362 (
            .O(N__36213),
            .I(N__36113));
    LocalMux I__8361 (
            .O(N__36210),
            .I(N__36110));
    ClkMux I__8360 (
            .O(N__36209),
            .I(N__36107));
    ClkMux I__8359 (
            .O(N__36208),
            .I(N__36104));
    ClkMux I__8358 (
            .O(N__36207),
            .I(N__36100));
    Span4Mux_v I__8357 (
            .O(N__36202),
            .I(N__36096));
    LocalMux I__8356 (
            .O(N__36199),
            .I(N__36093));
    ClkMux I__8355 (
            .O(N__36198),
            .I(N__36090));
    LocalMux I__8354 (
            .O(N__36195),
            .I(N__36087));
    ClkMux I__8353 (
            .O(N__36194),
            .I(N__36084));
    ClkMux I__8352 (
            .O(N__36193),
            .I(N__36081));
    ClkMux I__8351 (
            .O(N__36192),
            .I(N__36078));
    Span4Mux_v I__8350 (
            .O(N__36185),
            .I(N__36075));
    Span4Mux_s1_h I__8349 (
            .O(N__36182),
            .I(N__36072));
    Span4Mux_s2_h I__8348 (
            .O(N__36179),
            .I(N__36065));
    Span4Mux_h I__8347 (
            .O(N__36176),
            .I(N__36065));
    LocalMux I__8346 (
            .O(N__36173),
            .I(N__36065));
    Span4Mux_v I__8345 (
            .O(N__36168),
            .I(N__36062));
    ClkMux I__8344 (
            .O(N__36167),
            .I(N__36059));
    Span4Mux_h I__8343 (
            .O(N__36156),
            .I(N__36054));
    LocalMux I__8342 (
            .O(N__36153),
            .I(N__36054));
    Span4Mux_s2_h I__8341 (
            .O(N__36150),
            .I(N__36047));
    Span4Mux_v I__8340 (
            .O(N__36139),
            .I(N__36047));
    LocalMux I__8339 (
            .O(N__36136),
            .I(N__36047));
    Span4Mux_v I__8338 (
            .O(N__36131),
            .I(N__36040));
    Span4Mux_s2_h I__8337 (
            .O(N__36128),
            .I(N__36040));
    LocalMux I__8336 (
            .O(N__36125),
            .I(N__36040));
    Span4Mux_v I__8335 (
            .O(N__36116),
            .I(N__36031));
    IoSpan4Mux I__8334 (
            .O(N__36113),
            .I(N__36031));
    Span4Mux_v I__8333 (
            .O(N__36110),
            .I(N__36031));
    LocalMux I__8332 (
            .O(N__36107),
            .I(N__36031));
    LocalMux I__8331 (
            .O(N__36104),
            .I(N__36028));
    ClkMux I__8330 (
            .O(N__36103),
            .I(N__36025));
    LocalMux I__8329 (
            .O(N__36100),
            .I(N__36021));
    ClkMux I__8328 (
            .O(N__36099),
            .I(N__36018));
    Span4Mux_h I__8327 (
            .O(N__36096),
            .I(N__36011));
    Span4Mux_v I__8326 (
            .O(N__36093),
            .I(N__36011));
    LocalMux I__8325 (
            .O(N__36090),
            .I(N__36011));
    Span4Mux_h I__8324 (
            .O(N__36087),
            .I(N__36002));
    LocalMux I__8323 (
            .O(N__36084),
            .I(N__36002));
    LocalMux I__8322 (
            .O(N__36081),
            .I(N__36002));
    LocalMux I__8321 (
            .O(N__36078),
            .I(N__36002));
    Span4Mux_v I__8320 (
            .O(N__36075),
            .I(N__35994));
    Span4Mux_h I__8319 (
            .O(N__36072),
            .I(N__35994));
    Span4Mux_h I__8318 (
            .O(N__36065),
            .I(N__35994));
    Span4Mux_v I__8317 (
            .O(N__36062),
            .I(N__35989));
    LocalMux I__8316 (
            .O(N__36059),
            .I(N__35989));
    Span4Mux_h I__8315 (
            .O(N__36054),
            .I(N__35986));
    IoSpan4Mux I__8314 (
            .O(N__36047),
            .I(N__35979));
    IoSpan4Mux I__8313 (
            .O(N__36040),
            .I(N__35979));
    IoSpan4Mux I__8312 (
            .O(N__36031),
            .I(N__35979));
    Span4Mux_h I__8311 (
            .O(N__36028),
            .I(N__35974));
    LocalMux I__8310 (
            .O(N__36025),
            .I(N__35974));
    ClkMux I__8309 (
            .O(N__36024),
            .I(N__35971));
    Span12Mux_s5_h I__8308 (
            .O(N__36021),
            .I(N__35962));
    LocalMux I__8307 (
            .O(N__36018),
            .I(N__35962));
    Sp12to4 I__8306 (
            .O(N__36011),
            .I(N__35962));
    Sp12to4 I__8305 (
            .O(N__36002),
            .I(N__35962));
    ClkMux I__8304 (
            .O(N__36001),
            .I(N__35959));
    Odrv4 I__8303 (
            .O(N__35994),
            .I(fpga_osc));
    Odrv4 I__8302 (
            .O(N__35989),
            .I(fpga_osc));
    Odrv4 I__8301 (
            .O(N__35986),
            .I(fpga_osc));
    Odrv4 I__8300 (
            .O(N__35979),
            .I(fpga_osc));
    Odrv4 I__8299 (
            .O(N__35974),
            .I(fpga_osc));
    LocalMux I__8298 (
            .O(N__35971),
            .I(fpga_osc));
    Odrv12 I__8297 (
            .O(N__35962),
            .I(fpga_osc));
    LocalMux I__8296 (
            .O(N__35959),
            .I(fpga_osc));
    CEMux I__8295 (
            .O(N__35942),
            .I(N__35931));
    CEMux I__8294 (
            .O(N__35941),
            .I(N__35926));
    CEMux I__8293 (
            .O(N__35940),
            .I(N__35923));
    CEMux I__8292 (
            .O(N__35939),
            .I(N__35920));
    CEMux I__8291 (
            .O(N__35938),
            .I(N__35917));
    InMux I__8290 (
            .O(N__35937),
            .I(N__35908));
    InMux I__8289 (
            .O(N__35936),
            .I(N__35908));
    InMux I__8288 (
            .O(N__35935),
            .I(N__35908));
    InMux I__8287 (
            .O(N__35934),
            .I(N__35908));
    LocalMux I__8286 (
            .O(N__35931),
            .I(N__35905));
    InMux I__8285 (
            .O(N__35930),
            .I(N__35902));
    InMux I__8284 (
            .O(N__35929),
            .I(N__35899));
    LocalMux I__8283 (
            .O(N__35926),
            .I(N__35892));
    LocalMux I__8282 (
            .O(N__35923),
            .I(N__35883));
    LocalMux I__8281 (
            .O(N__35920),
            .I(N__35880));
    LocalMux I__8280 (
            .O(N__35917),
            .I(N__35875));
    LocalMux I__8279 (
            .O(N__35908),
            .I(N__35875));
    Span4Mux_s3_v I__8278 (
            .O(N__35905),
            .I(N__35868));
    LocalMux I__8277 (
            .O(N__35902),
            .I(N__35868));
    LocalMux I__8276 (
            .O(N__35899),
            .I(N__35868));
    InMux I__8275 (
            .O(N__35898),
            .I(N__35859));
    InMux I__8274 (
            .O(N__35897),
            .I(N__35859));
    InMux I__8273 (
            .O(N__35896),
            .I(N__35859));
    InMux I__8272 (
            .O(N__35895),
            .I(N__35859));
    Span4Mux_s2_h I__8271 (
            .O(N__35892),
            .I(N__35856));
    InMux I__8270 (
            .O(N__35891),
            .I(N__35843));
    InMux I__8269 (
            .O(N__35890),
            .I(N__35843));
    InMux I__8268 (
            .O(N__35889),
            .I(N__35843));
    InMux I__8267 (
            .O(N__35888),
            .I(N__35843));
    InMux I__8266 (
            .O(N__35887),
            .I(N__35843));
    InMux I__8265 (
            .O(N__35886),
            .I(N__35843));
    Span4Mux_s0_h I__8264 (
            .O(N__35883),
            .I(N__35834));
    Span4Mux_v I__8263 (
            .O(N__35880),
            .I(N__35834));
    Span4Mux_s3_v I__8262 (
            .O(N__35875),
            .I(N__35834));
    Span4Mux_v I__8261 (
            .O(N__35868),
            .I(N__35834));
    LocalMux I__8260 (
            .O(N__35859),
            .I(N__35831));
    Odrv4 I__8259 (
            .O(N__35856),
            .I(\b2v_inst11.dutycycle_RNIHJNV7Z0Z_0 ));
    LocalMux I__8258 (
            .O(N__35843),
            .I(\b2v_inst11.dutycycle_RNIHJNV7Z0Z_0 ));
    Odrv4 I__8257 (
            .O(N__35834),
            .I(\b2v_inst11.dutycycle_RNIHJNV7Z0Z_0 ));
    Odrv4 I__8256 (
            .O(N__35831),
            .I(\b2v_inst11.dutycycle_RNIHJNV7Z0Z_0 ));
    CascadeMux I__8255 (
            .O(N__35822),
            .I(\b2v_inst11.count_offZ0Z_9_cascade_ ));
    InMux I__8254 (
            .O(N__35819),
            .I(N__35816));
    LocalMux I__8253 (
            .O(N__35816),
            .I(\b2v_inst11.un34_clk_100khz_11 ));
    CascadeMux I__8252 (
            .O(N__35813),
            .I(N__35809));
    InMux I__8251 (
            .O(N__35812),
            .I(N__35806));
    InMux I__8250 (
            .O(N__35809),
            .I(N__35803));
    LocalMux I__8249 (
            .O(N__35806),
            .I(\b2v_inst11.count_offZ0Z_10 ));
    LocalMux I__8248 (
            .O(N__35803),
            .I(\b2v_inst11.count_offZ0Z_10 ));
    InMux I__8247 (
            .O(N__35798),
            .I(N__35792));
    InMux I__8246 (
            .O(N__35797),
            .I(N__35792));
    LocalMux I__8245 (
            .O(N__35792),
            .I(\b2v_inst11.count_off_1_10 ));
    InMux I__8244 (
            .O(N__35789),
            .I(N__35786));
    LocalMux I__8243 (
            .O(N__35786),
            .I(\b2v_inst11.count_off_0_10 ));
    InMux I__8242 (
            .O(N__35783),
            .I(N__35779));
    InMux I__8241 (
            .O(N__35782),
            .I(N__35776));
    LocalMux I__8240 (
            .O(N__35779),
            .I(\b2v_inst11.count_offZ0Z_11 ));
    LocalMux I__8239 (
            .O(N__35776),
            .I(\b2v_inst11.count_offZ0Z_11 ));
    InMux I__8238 (
            .O(N__35771),
            .I(N__35765));
    InMux I__8237 (
            .O(N__35770),
            .I(N__35765));
    LocalMux I__8236 (
            .O(N__35765),
            .I(\b2v_inst11.count_off_1_11 ));
    InMux I__8235 (
            .O(N__35762),
            .I(N__35759));
    LocalMux I__8234 (
            .O(N__35759),
            .I(\b2v_inst11.count_off_0_11 ));
    InMux I__8233 (
            .O(N__35756),
            .I(N__35752));
    InMux I__8232 (
            .O(N__35755),
            .I(N__35749));
    LocalMux I__8231 (
            .O(N__35752),
            .I(\b2v_inst11.count_offZ0Z_12 ));
    LocalMux I__8230 (
            .O(N__35749),
            .I(\b2v_inst11.count_offZ0Z_12 ));
    InMux I__8229 (
            .O(N__35744),
            .I(N__35740));
    InMux I__8228 (
            .O(N__35743),
            .I(N__35737));
    LocalMux I__8227 (
            .O(N__35740),
            .I(\b2v_inst11.count_off_1_12 ));
    LocalMux I__8226 (
            .O(N__35737),
            .I(\b2v_inst11.count_off_1_12 ));
    InMux I__8225 (
            .O(N__35732),
            .I(N__35729));
    LocalMux I__8224 (
            .O(N__35729),
            .I(\b2v_inst11.count_off_0_12 ));
    InMux I__8223 (
            .O(N__35726),
            .I(N__35722));
    InMux I__8222 (
            .O(N__35725),
            .I(N__35719));
    LocalMux I__8221 (
            .O(N__35722),
            .I(N__35716));
    LocalMux I__8220 (
            .O(N__35719),
            .I(\b2v_inst11.count_off_1_13 ));
    Odrv4 I__8219 (
            .O(N__35716),
            .I(\b2v_inst11.count_off_1_13 ));
    InMux I__8218 (
            .O(N__35711),
            .I(N__35708));
    LocalMux I__8217 (
            .O(N__35708),
            .I(N__35705));
    Span4Mux_h I__8216 (
            .O(N__35705),
            .I(N__35702));
    Odrv4 I__8215 (
            .O(N__35702),
            .I(\b2v_inst11.count_off_0_13 ));
    InMux I__8214 (
            .O(N__35699),
            .I(N__35696));
    LocalMux I__8213 (
            .O(N__35696),
            .I(N__35692));
    InMux I__8212 (
            .O(N__35695),
            .I(N__35689));
    Span4Mux_h I__8211 (
            .O(N__35692),
            .I(N__35686));
    LocalMux I__8210 (
            .O(N__35689),
            .I(\b2v_inst11.count_off_1_2 ));
    Odrv4 I__8209 (
            .O(N__35686),
            .I(\b2v_inst11.count_off_1_2 ));
    InMux I__8208 (
            .O(N__35681),
            .I(N__35678));
    LocalMux I__8207 (
            .O(N__35678),
            .I(N__35675));
    Odrv4 I__8206 (
            .O(N__35675),
            .I(\b2v_inst11.count_off_0_2 ));
    InMux I__8205 (
            .O(N__35672),
            .I(N__35668));
    InMux I__8204 (
            .O(N__35671),
            .I(N__35665));
    LocalMux I__8203 (
            .O(N__35668),
            .I(N__35662));
    LocalMux I__8202 (
            .O(N__35665),
            .I(N__35659));
    Odrv4 I__8201 (
            .O(N__35662),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    Odrv4 I__8200 (
            .O(N__35659),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    InMux I__8199 (
            .O(N__35654),
            .I(N__35650));
    InMux I__8198 (
            .O(N__35653),
            .I(N__35647));
    LocalMux I__8197 (
            .O(N__35650),
            .I(N__35644));
    LocalMux I__8196 (
            .O(N__35647),
            .I(N__35641));
    Span4Mux_v I__8195 (
            .O(N__35644),
            .I(N__35638));
    Span4Mux_s2_h I__8194 (
            .O(N__35641),
            .I(N__35635));
    Odrv4 I__8193 (
            .O(N__35638),
            .I(\b2v_inst11.count_offZ0Z_5 ));
    Odrv4 I__8192 (
            .O(N__35635),
            .I(\b2v_inst11.count_offZ0Z_5 ));
    CascadeMux I__8191 (
            .O(N__35630),
            .I(\b2v_inst11.count_offZ0Z_1_cascade_ ));
    InMux I__8190 (
            .O(N__35627),
            .I(N__35623));
    InMux I__8189 (
            .O(N__35626),
            .I(N__35620));
    LocalMux I__8188 (
            .O(N__35623),
            .I(N__35617));
    LocalMux I__8187 (
            .O(N__35620),
            .I(N__35614));
    Span4Mux_v I__8186 (
            .O(N__35617),
            .I(N__35611));
    Span4Mux_s2_h I__8185 (
            .O(N__35614),
            .I(N__35608));
    Odrv4 I__8184 (
            .O(N__35611),
            .I(\b2v_inst11.count_offZ0Z_2 ));
    Odrv4 I__8183 (
            .O(N__35608),
            .I(\b2v_inst11.count_offZ0Z_2 ));
    CascadeMux I__8182 (
            .O(N__35603),
            .I(\b2v_inst11.un34_clk_100khz_9_cascade_ ));
    InMux I__8181 (
            .O(N__35600),
            .I(N__35596));
    CascadeMux I__8180 (
            .O(N__35599),
            .I(N__35591));
    LocalMux I__8179 (
            .O(N__35596),
            .I(N__35588));
    InMux I__8178 (
            .O(N__35595),
            .I(N__35578));
    InMux I__8177 (
            .O(N__35594),
            .I(N__35578));
    InMux I__8176 (
            .O(N__35591),
            .I(N__35574));
    Span4Mux_v I__8175 (
            .O(N__35588),
            .I(N__35571));
    InMux I__8174 (
            .O(N__35587),
            .I(N__35568));
    InMux I__8173 (
            .O(N__35586),
            .I(N__35561));
    InMux I__8172 (
            .O(N__35585),
            .I(N__35561));
    InMux I__8171 (
            .O(N__35584),
            .I(N__35561));
    InMux I__8170 (
            .O(N__35583),
            .I(N__35558));
    LocalMux I__8169 (
            .O(N__35578),
            .I(N__35555));
    InMux I__8168 (
            .O(N__35577),
            .I(N__35552));
    LocalMux I__8167 (
            .O(N__35574),
            .I(N__35549));
    Span4Mux_v I__8166 (
            .O(N__35571),
            .I(N__35542));
    LocalMux I__8165 (
            .O(N__35568),
            .I(N__35542));
    LocalMux I__8164 (
            .O(N__35561),
            .I(N__35542));
    LocalMux I__8163 (
            .O(N__35558),
            .I(N__35537));
    Span4Mux_h I__8162 (
            .O(N__35555),
            .I(N__35537));
    LocalMux I__8161 (
            .O(N__35552),
            .I(\b2v_inst11.count_off_RNI_0Z0Z_1 ));
    Odrv12 I__8160 (
            .O(N__35549),
            .I(\b2v_inst11.count_off_RNI_0Z0Z_1 ));
    Odrv4 I__8159 (
            .O(N__35542),
            .I(\b2v_inst11.count_off_RNI_0Z0Z_1 ));
    Odrv4 I__8158 (
            .O(N__35537),
            .I(\b2v_inst11.count_off_RNI_0Z0Z_1 ));
    InMux I__8157 (
            .O(N__35528),
            .I(N__35525));
    LocalMux I__8156 (
            .O(N__35525),
            .I(N__35521));
    InMux I__8155 (
            .O(N__35524),
            .I(N__35518));
    Odrv4 I__8154 (
            .O(N__35521),
            .I(\b2v_inst11.count_offZ0Z_15 ));
    LocalMux I__8153 (
            .O(N__35518),
            .I(\b2v_inst11.count_offZ0Z_15 ));
    InMux I__8152 (
            .O(N__35513),
            .I(N__35510));
    LocalMux I__8151 (
            .O(N__35510),
            .I(N__35507));
    Span4Mux_s2_h I__8150 (
            .O(N__35507),
            .I(N__35503));
    InMux I__8149 (
            .O(N__35506),
            .I(N__35500));
    Span4Mux_h I__8148 (
            .O(N__35503),
            .I(N__35497));
    LocalMux I__8147 (
            .O(N__35500),
            .I(N__35494));
    Odrv4 I__8146 (
            .O(N__35497),
            .I(\b2v_inst11.count_offZ0Z_13 ));
    Odrv4 I__8145 (
            .O(N__35494),
            .I(\b2v_inst11.count_offZ0Z_13 ));
    CascadeMux I__8144 (
            .O(N__35489),
            .I(N__35486));
    InMux I__8143 (
            .O(N__35486),
            .I(N__35483));
    LocalMux I__8142 (
            .O(N__35483),
            .I(N__35479));
    InMux I__8141 (
            .O(N__35482),
            .I(N__35476));
    Span4Mux_v I__8140 (
            .O(N__35479),
            .I(N__35471));
    LocalMux I__8139 (
            .O(N__35476),
            .I(N__35471));
    Odrv4 I__8138 (
            .O(N__35471),
            .I(\b2v_inst11.count_offZ0Z_14 ));
    InMux I__8137 (
            .O(N__35468),
            .I(N__35465));
    LocalMux I__8136 (
            .O(N__35465),
            .I(\b2v_inst11.un34_clk_100khz_10 ));
    InMux I__8135 (
            .O(N__35462),
            .I(N__35459));
    LocalMux I__8134 (
            .O(N__35459),
            .I(N__35455));
    InMux I__8133 (
            .O(N__35458),
            .I(N__35452));
    Span4Mux_v I__8132 (
            .O(N__35455),
            .I(N__35449));
    LocalMux I__8131 (
            .O(N__35452),
            .I(N__35446));
    Odrv4 I__8130 (
            .O(N__35449),
            .I(\b2v_inst11.count_offZ0Z_7 ));
    Odrv4 I__8129 (
            .O(N__35446),
            .I(\b2v_inst11.count_offZ0Z_7 ));
    InMux I__8128 (
            .O(N__35441),
            .I(N__35438));
    LocalMux I__8127 (
            .O(N__35438),
            .I(N__35434));
    InMux I__8126 (
            .O(N__35437),
            .I(N__35431));
    Span4Mux_s1_h I__8125 (
            .O(N__35434),
            .I(N__35428));
    LocalMux I__8124 (
            .O(N__35431),
            .I(N__35425));
    Odrv4 I__8123 (
            .O(N__35428),
            .I(\b2v_inst11.count_offZ0Z_8 ));
    Odrv12 I__8122 (
            .O(N__35425),
            .I(\b2v_inst11.count_offZ0Z_8 ));
    CascadeMux I__8121 (
            .O(N__35420),
            .I(N__35417));
    InMux I__8120 (
            .O(N__35417),
            .I(N__35413));
    InMux I__8119 (
            .O(N__35416),
            .I(N__35410));
    LocalMux I__8118 (
            .O(N__35413),
            .I(N__35407));
    LocalMux I__8117 (
            .O(N__35410),
            .I(N__35404));
    Span4Mux_v I__8116 (
            .O(N__35407),
            .I(N__35401));
    Span4Mux_s2_h I__8115 (
            .O(N__35404),
            .I(N__35398));
    Odrv4 I__8114 (
            .O(N__35401),
            .I(\b2v_inst11.count_offZ0Z_3 ));
    Odrv4 I__8113 (
            .O(N__35398),
            .I(\b2v_inst11.count_offZ0Z_3 ));
    InMux I__8112 (
            .O(N__35393),
            .I(N__35389));
    InMux I__8111 (
            .O(N__35392),
            .I(N__35386));
    LocalMux I__8110 (
            .O(N__35389),
            .I(N__35383));
    LocalMux I__8109 (
            .O(N__35386),
            .I(N__35380));
    Span4Mux_s3_h I__8108 (
            .O(N__35383),
            .I(N__35377));
    Span4Mux_s2_h I__8107 (
            .O(N__35380),
            .I(N__35374));
    Odrv4 I__8106 (
            .O(N__35377),
            .I(\b2v_inst11.count_offZ0Z_4 ));
    Odrv4 I__8105 (
            .O(N__35374),
            .I(\b2v_inst11.count_offZ0Z_4 ));
    InMux I__8104 (
            .O(N__35369),
            .I(N__35366));
    LocalMux I__8103 (
            .O(N__35366),
            .I(\b2v_inst11.un34_clk_100khz_8 ));
    CascadeMux I__8102 (
            .O(N__35363),
            .I(N__35359));
    InMux I__8101 (
            .O(N__35362),
            .I(N__35355));
    InMux I__8100 (
            .O(N__35359),
            .I(N__35352));
    InMux I__8099 (
            .O(N__35358),
            .I(N__35349));
    LocalMux I__8098 (
            .O(N__35355),
            .I(N__35344));
    LocalMux I__8097 (
            .O(N__35352),
            .I(N__35344));
    LocalMux I__8096 (
            .O(N__35349),
            .I(\b2v_inst11.count_offZ0Z_1 ));
    Odrv4 I__8095 (
            .O(N__35344),
            .I(\b2v_inst11.count_offZ0Z_1 ));
    InMux I__8094 (
            .O(N__35339),
            .I(N__35336));
    LocalMux I__8093 (
            .O(N__35336),
            .I(\b2v_inst11.count_off_0_1 ));
    CascadeMux I__8092 (
            .O(N__35333),
            .I(N__35329));
    InMux I__8091 (
            .O(N__35332),
            .I(N__35318));
    InMux I__8090 (
            .O(N__35329),
            .I(N__35318));
    InMux I__8089 (
            .O(N__35328),
            .I(N__35318));
    InMux I__8088 (
            .O(N__35327),
            .I(N__35315));
    InMux I__8087 (
            .O(N__35326),
            .I(N__35310));
    InMux I__8086 (
            .O(N__35325),
            .I(N__35310));
    LocalMux I__8085 (
            .O(N__35318),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    LocalMux I__8084 (
            .O(N__35315),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    LocalMux I__8083 (
            .O(N__35310),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    InMux I__8082 (
            .O(N__35303),
            .I(N__35288));
    InMux I__8081 (
            .O(N__35302),
            .I(N__35288));
    InMux I__8080 (
            .O(N__35301),
            .I(N__35288));
    InMux I__8079 (
            .O(N__35300),
            .I(N__35279));
    InMux I__8078 (
            .O(N__35299),
            .I(N__35279));
    InMux I__8077 (
            .O(N__35298),
            .I(N__35279));
    InMux I__8076 (
            .O(N__35297),
            .I(N__35279));
    InMux I__8075 (
            .O(N__35296),
            .I(N__35266));
    InMux I__8074 (
            .O(N__35295),
            .I(N__35266));
    LocalMux I__8073 (
            .O(N__35288),
            .I(N__35261));
    LocalMux I__8072 (
            .O(N__35279),
            .I(N__35261));
    InMux I__8071 (
            .O(N__35278),
            .I(N__35254));
    InMux I__8070 (
            .O(N__35277),
            .I(N__35254));
    InMux I__8069 (
            .O(N__35276),
            .I(N__35254));
    InMux I__8068 (
            .O(N__35275),
            .I(N__35245));
    InMux I__8067 (
            .O(N__35274),
            .I(N__35245));
    InMux I__8066 (
            .O(N__35273),
            .I(N__35245));
    InMux I__8065 (
            .O(N__35272),
            .I(N__35245));
    InMux I__8064 (
            .O(N__35271),
            .I(N__35242));
    LocalMux I__8063 (
            .O(N__35266),
            .I(\b2v_inst11.N_125 ));
    Odrv4 I__8062 (
            .O(N__35261),
            .I(\b2v_inst11.N_125 ));
    LocalMux I__8061 (
            .O(N__35254),
            .I(\b2v_inst11.N_125 ));
    LocalMux I__8060 (
            .O(N__35245),
            .I(\b2v_inst11.N_125 ));
    LocalMux I__8059 (
            .O(N__35242),
            .I(\b2v_inst11.N_125 ));
    InMux I__8058 (
            .O(N__35231),
            .I(N__35228));
    LocalMux I__8057 (
            .O(N__35228),
            .I(\b2v_inst11.count_off_0_0 ));
    InMux I__8056 (
            .O(N__35225),
            .I(N__35222));
    LocalMux I__8055 (
            .O(N__35222),
            .I(\b2v_inst11.count_off_0_9 ));
    InMux I__8054 (
            .O(N__35219),
            .I(N__35213));
    InMux I__8053 (
            .O(N__35218),
            .I(N__35213));
    LocalMux I__8052 (
            .O(N__35213),
            .I(\b2v_inst11.count_off_1_9 ));
    InMux I__8051 (
            .O(N__35210),
            .I(N__35207));
    LocalMux I__8050 (
            .O(N__35207),
            .I(\b2v_inst11.count_offZ0Z_9 ));
    CascadeMux I__8049 (
            .O(N__35204),
            .I(N__35201));
    InMux I__8048 (
            .O(N__35201),
            .I(N__35193));
    InMux I__8047 (
            .O(N__35200),
            .I(N__35193));
    InMux I__8046 (
            .O(N__35199),
            .I(N__35189));
    CascadeMux I__8045 (
            .O(N__35198),
            .I(N__35185));
    LocalMux I__8044 (
            .O(N__35193),
            .I(N__35179));
    InMux I__8043 (
            .O(N__35192),
            .I(N__35176));
    LocalMux I__8042 (
            .O(N__35189),
            .I(N__35172));
    InMux I__8041 (
            .O(N__35188),
            .I(N__35167));
    InMux I__8040 (
            .O(N__35185),
            .I(N__35167));
    InMux I__8039 (
            .O(N__35184),
            .I(N__35164));
    InMux I__8038 (
            .O(N__35183),
            .I(N__35161));
    InMux I__8037 (
            .O(N__35182),
            .I(N__35158));
    Span4Mux_v I__8036 (
            .O(N__35179),
            .I(N__35155));
    LocalMux I__8035 (
            .O(N__35176),
            .I(N__35152));
    InMux I__8034 (
            .O(N__35175),
            .I(N__35149));
    Span4Mux_s1_h I__8033 (
            .O(N__35172),
            .I(N__35146));
    LocalMux I__8032 (
            .O(N__35167),
            .I(N__35139));
    LocalMux I__8031 (
            .O(N__35164),
            .I(N__35139));
    LocalMux I__8030 (
            .O(N__35161),
            .I(N__35139));
    LocalMux I__8029 (
            .O(N__35158),
            .I(N__35136));
    Span4Mux_h I__8028 (
            .O(N__35155),
            .I(N__35128));
    Span4Mux_h I__8027 (
            .O(N__35152),
            .I(N__35128));
    LocalMux I__8026 (
            .O(N__35149),
            .I(N__35128));
    Span4Mux_h I__8025 (
            .O(N__35146),
            .I(N__35121));
    Span4Mux_v I__8024 (
            .O(N__35139),
            .I(N__35121));
    Span4Mux_h I__8023 (
            .O(N__35136),
            .I(N__35121));
    InMux I__8022 (
            .O(N__35135),
            .I(N__35118));
    Odrv4 I__8021 (
            .O(N__35128),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__8020 (
            .O(N__35121),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    LocalMux I__8019 (
            .O(N__35118),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    InMux I__8018 (
            .O(N__35111),
            .I(N__35097));
    InMux I__8017 (
            .O(N__35110),
            .I(N__35097));
    InMux I__8016 (
            .O(N__35109),
            .I(N__35097));
    CascadeMux I__8015 (
            .O(N__35108),
            .I(N__35085));
    InMux I__8014 (
            .O(N__35107),
            .I(N__35078));
    InMux I__8013 (
            .O(N__35106),
            .I(N__35078));
    InMux I__8012 (
            .O(N__35105),
            .I(N__35073));
    InMux I__8011 (
            .O(N__35104),
            .I(N__35073));
    LocalMux I__8010 (
            .O(N__35097),
            .I(N__35069));
    InMux I__8009 (
            .O(N__35096),
            .I(N__35066));
    CascadeMux I__8008 (
            .O(N__35095),
            .I(N__35063));
    InMux I__8007 (
            .O(N__35094),
            .I(N__35059));
    InMux I__8006 (
            .O(N__35093),
            .I(N__35052));
    InMux I__8005 (
            .O(N__35092),
            .I(N__35052));
    InMux I__8004 (
            .O(N__35091),
            .I(N__35052));
    InMux I__8003 (
            .O(N__35090),
            .I(N__35045));
    InMux I__8002 (
            .O(N__35089),
            .I(N__35045));
    InMux I__8001 (
            .O(N__35088),
            .I(N__35045));
    InMux I__8000 (
            .O(N__35085),
            .I(N__35040));
    InMux I__7999 (
            .O(N__35084),
            .I(N__35040));
    InMux I__7998 (
            .O(N__35083),
            .I(N__35037));
    LocalMux I__7997 (
            .O(N__35078),
            .I(N__35032));
    LocalMux I__7996 (
            .O(N__35073),
            .I(N__35032));
    CascadeMux I__7995 (
            .O(N__35072),
            .I(N__35027));
    Span4Mux_s2_h I__7994 (
            .O(N__35069),
            .I(N__35022));
    LocalMux I__7993 (
            .O(N__35066),
            .I(N__35019));
    InMux I__7992 (
            .O(N__35063),
            .I(N__35014));
    InMux I__7991 (
            .O(N__35062),
            .I(N__35014));
    LocalMux I__7990 (
            .O(N__35059),
            .I(N__35007));
    LocalMux I__7989 (
            .O(N__35052),
            .I(N__35007));
    LocalMux I__7988 (
            .O(N__35045),
            .I(N__35007));
    LocalMux I__7987 (
            .O(N__35040),
            .I(N__35004));
    LocalMux I__7986 (
            .O(N__35037),
            .I(N__34999));
    Span4Mux_v I__7985 (
            .O(N__35032),
            .I(N__34999));
    InMux I__7984 (
            .O(N__35031),
            .I(N__34996));
    InMux I__7983 (
            .O(N__35030),
            .I(N__34991));
    InMux I__7982 (
            .O(N__35027),
            .I(N__34991));
    InMux I__7981 (
            .O(N__35026),
            .I(N__34986));
    InMux I__7980 (
            .O(N__35025),
            .I(N__34986));
    Span4Mux_v I__7979 (
            .O(N__35022),
            .I(N__34983));
    Span4Mux_v I__7978 (
            .O(N__35019),
            .I(N__34976));
    LocalMux I__7977 (
            .O(N__35014),
            .I(N__34976));
    Span4Mux_s3_h I__7976 (
            .O(N__35007),
            .I(N__34976));
    Odrv12 I__7975 (
            .O(N__35004),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    Odrv4 I__7974 (
            .O(N__34999),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__7973 (
            .O(N__34996),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__7972 (
            .O(N__34991),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__7971 (
            .O(N__34986),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    Odrv4 I__7970 (
            .O(N__34983),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    Odrv4 I__7969 (
            .O(N__34976),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    InMux I__7968 (
            .O(N__34961),
            .I(N__34958));
    LocalMux I__7967 (
            .O(N__34958),
            .I(N__34955));
    Span4Mux_v I__7966 (
            .O(N__34955),
            .I(N__34952));
    Odrv4 I__7965 (
            .O(N__34952),
            .I(G_6_i_a3_1));
    CascadeMux I__7964 (
            .O(N__34949),
            .I(N_5_cascade_));
    IoInMux I__7963 (
            .O(N__34946),
            .I(N__34942));
    IoInMux I__7962 (
            .O(N__34945),
            .I(N__34939));
    LocalMux I__7961 (
            .O(N__34942),
            .I(N__34933));
    LocalMux I__7960 (
            .O(N__34939),
            .I(N__34933));
    CascadeMux I__7959 (
            .O(N__34938),
            .I(N__34923));
    IoSpan4Mux I__7958 (
            .O(N__34933),
            .I(N__34920));
    InMux I__7957 (
            .O(N__34932),
            .I(N__34916));
    InMux I__7956 (
            .O(N__34931),
            .I(N__34913));
    InMux I__7955 (
            .O(N__34930),
            .I(N__34910));
    InMux I__7954 (
            .O(N__34929),
            .I(N__34907));
    InMux I__7953 (
            .O(N__34928),
            .I(N__34904));
    InMux I__7952 (
            .O(N__34927),
            .I(N__34901));
    InMux I__7951 (
            .O(N__34926),
            .I(N__34898));
    InMux I__7950 (
            .O(N__34923),
            .I(N__34895));
    Span4Mux_s3_h I__7949 (
            .O(N__34920),
            .I(N__34891));
    InMux I__7948 (
            .O(N__34919),
            .I(N__34888));
    LocalMux I__7947 (
            .O(N__34916),
            .I(N__34885));
    LocalMux I__7946 (
            .O(N__34913),
            .I(N__34878));
    LocalMux I__7945 (
            .O(N__34910),
            .I(N__34878));
    LocalMux I__7944 (
            .O(N__34907),
            .I(N__34875));
    LocalMux I__7943 (
            .O(N__34904),
            .I(N__34870));
    LocalMux I__7942 (
            .O(N__34901),
            .I(N__34870));
    LocalMux I__7941 (
            .O(N__34898),
            .I(N__34865));
    LocalMux I__7940 (
            .O(N__34895),
            .I(N__34865));
    InMux I__7939 (
            .O(N__34894),
            .I(N__34862));
    Span4Mux_h I__7938 (
            .O(N__34891),
            .I(N__34857));
    LocalMux I__7937 (
            .O(N__34888),
            .I(N__34857));
    Span4Mux_v I__7936 (
            .O(N__34885),
            .I(N__34854));
    InMux I__7935 (
            .O(N__34884),
            .I(N__34849));
    InMux I__7934 (
            .O(N__34883),
            .I(N__34849));
    Span12Mux_s3_h I__7933 (
            .O(N__34878),
            .I(N__34846));
    Span4Mux_v I__7932 (
            .O(N__34875),
            .I(N__34837));
    Span4Mux_s3_h I__7931 (
            .O(N__34870),
            .I(N__34837));
    Span4Mux_s3_h I__7930 (
            .O(N__34865),
            .I(N__34837));
    LocalMux I__7929 (
            .O(N__34862),
            .I(N__34837));
    Odrv4 I__7928 (
            .O(N__34857),
            .I(v5s_enn));
    Odrv4 I__7927 (
            .O(N__34854),
            .I(v5s_enn));
    LocalMux I__7926 (
            .O(N__34849),
            .I(v5s_enn));
    Odrv12 I__7925 (
            .O(N__34846),
            .I(v5s_enn));
    Odrv4 I__7924 (
            .O(N__34837),
            .I(v5s_enn));
    InMux I__7923 (
            .O(N__34826),
            .I(N__34823));
    LocalMux I__7922 (
            .O(N__34823),
            .I(N__34820));
    Odrv12 I__7921 (
            .O(N__34820),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_rn_1 ));
    CascadeMux I__7920 (
            .O(N__34817),
            .I(b2v_inst11_un1_clk_100khz_52_and_i_0_cascade_));
    InMux I__7919 (
            .O(N__34814),
            .I(N__34801));
    InMux I__7918 (
            .O(N__34813),
            .I(N__34792));
    InMux I__7917 (
            .O(N__34812),
            .I(N__34787));
    InMux I__7916 (
            .O(N__34811),
            .I(N__34787));
    InMux I__7915 (
            .O(N__34810),
            .I(N__34784));
    InMux I__7914 (
            .O(N__34809),
            .I(N__34779));
    InMux I__7913 (
            .O(N__34808),
            .I(N__34779));
    InMux I__7912 (
            .O(N__34807),
            .I(N__34776));
    InMux I__7911 (
            .O(N__34806),
            .I(N__34773));
    InMux I__7910 (
            .O(N__34805),
            .I(N__34770));
    InMux I__7909 (
            .O(N__34804),
            .I(N__34767));
    LocalMux I__7908 (
            .O(N__34801),
            .I(N__34764));
    InMux I__7907 (
            .O(N__34800),
            .I(N__34757));
    InMux I__7906 (
            .O(N__34799),
            .I(N__34757));
    InMux I__7905 (
            .O(N__34798),
            .I(N__34757));
    InMux I__7904 (
            .O(N__34797),
            .I(N__34752));
    InMux I__7903 (
            .O(N__34796),
            .I(N__34752));
    InMux I__7902 (
            .O(N__34795),
            .I(N__34749));
    LocalMux I__7901 (
            .O(N__34792),
            .I(N__34744));
    LocalMux I__7900 (
            .O(N__34787),
            .I(N__34740));
    LocalMux I__7899 (
            .O(N__34784),
            .I(N__34732));
    LocalMux I__7898 (
            .O(N__34779),
            .I(N__34732));
    LocalMux I__7897 (
            .O(N__34776),
            .I(N__34717));
    LocalMux I__7896 (
            .O(N__34773),
            .I(N__34717));
    LocalMux I__7895 (
            .O(N__34770),
            .I(N__34717));
    LocalMux I__7894 (
            .O(N__34767),
            .I(N__34717));
    Span4Mux_h I__7893 (
            .O(N__34764),
            .I(N__34717));
    LocalMux I__7892 (
            .O(N__34757),
            .I(N__34717));
    LocalMux I__7891 (
            .O(N__34752),
            .I(N__34717));
    LocalMux I__7890 (
            .O(N__34749),
            .I(N__34714));
    InMux I__7889 (
            .O(N__34748),
            .I(N__34711));
    InMux I__7888 (
            .O(N__34747),
            .I(N__34708));
    Span4Mux_s3_h I__7887 (
            .O(N__34744),
            .I(N__34705));
    InMux I__7886 (
            .O(N__34743),
            .I(N__34702));
    Span4Mux_h I__7885 (
            .O(N__34740),
            .I(N__34699));
    InMux I__7884 (
            .O(N__34739),
            .I(N__34694));
    InMux I__7883 (
            .O(N__34738),
            .I(N__34694));
    InMux I__7882 (
            .O(N__34737),
            .I(N__34691));
    Span4Mux_v I__7881 (
            .O(N__34732),
            .I(N__34686));
    Span4Mux_v I__7880 (
            .O(N__34717),
            .I(N__34686));
    Span4Mux_s2_h I__7879 (
            .O(N__34714),
            .I(N__34683));
    LocalMux I__7878 (
            .O(N__34711),
            .I(N__34678));
    LocalMux I__7877 (
            .O(N__34708),
            .I(N__34678));
    Odrv4 I__7876 (
            .O(N__34705),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    LocalMux I__7875 (
            .O(N__34702),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv4 I__7874 (
            .O(N__34699),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    LocalMux I__7873 (
            .O(N__34694),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    LocalMux I__7872 (
            .O(N__34691),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv4 I__7871 (
            .O(N__34686),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv4 I__7870 (
            .O(N__34683),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv12 I__7869 (
            .O(N__34678),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    InMux I__7868 (
            .O(N__34661),
            .I(N__34658));
    LocalMux I__7867 (
            .O(N__34658),
            .I(N__34655));
    Odrv12 I__7866 (
            .O(N__34655),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_sn ));
    CascadeMux I__7865 (
            .O(N__34652),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_0_cascade_ ));
    InMux I__7864 (
            .O(N__34649),
            .I(N__34646));
    LocalMux I__7863 (
            .O(N__34646),
            .I(\b2v_inst11.N_6063_0_0 ));
    InMux I__7862 (
            .O(N__34643),
            .I(N__34637));
    InMux I__7861 (
            .O(N__34642),
            .I(N__34637));
    LocalMux I__7860 (
            .O(N__34637),
            .I(N__34634));
    Span4Mux_h I__7859 (
            .O(N__34634),
            .I(N__34631));
    Span4Mux_h I__7858 (
            .O(N__34631),
            .I(N__34628));
    Odrv4 I__7857 (
            .O(N__34628),
            .I(\b2v_inst11.dutycycle_eena_14_0_0 ));
    InMux I__7856 (
            .O(N__34625),
            .I(N__34616));
    InMux I__7855 (
            .O(N__34624),
            .I(N__34611));
    InMux I__7854 (
            .O(N__34623),
            .I(N__34608));
    CascadeMux I__7853 (
            .O(N__34622),
            .I(N__34605));
    InMux I__7852 (
            .O(N__34621),
            .I(N__34596));
    InMux I__7851 (
            .O(N__34620),
            .I(N__34593));
    InMux I__7850 (
            .O(N__34619),
            .I(N__34590));
    LocalMux I__7849 (
            .O(N__34616),
            .I(N__34587));
    InMux I__7848 (
            .O(N__34615),
            .I(N__34584));
    InMux I__7847 (
            .O(N__34614),
            .I(N__34581));
    LocalMux I__7846 (
            .O(N__34611),
            .I(N__34578));
    LocalMux I__7845 (
            .O(N__34608),
            .I(N__34575));
    InMux I__7844 (
            .O(N__34605),
            .I(N__34572));
    InMux I__7843 (
            .O(N__34604),
            .I(N__34569));
    InMux I__7842 (
            .O(N__34603),
            .I(N__34566));
    InMux I__7841 (
            .O(N__34602),
            .I(N__34563));
    InMux I__7840 (
            .O(N__34601),
            .I(N__34556));
    InMux I__7839 (
            .O(N__34600),
            .I(N__34556));
    InMux I__7838 (
            .O(N__34599),
            .I(N__34556));
    LocalMux I__7837 (
            .O(N__34596),
            .I(N__34550));
    LocalMux I__7836 (
            .O(N__34593),
            .I(N__34550));
    LocalMux I__7835 (
            .O(N__34590),
            .I(N__34547));
    Span4Mux_v I__7834 (
            .O(N__34587),
            .I(N__34544));
    LocalMux I__7833 (
            .O(N__34584),
            .I(N__34539));
    LocalMux I__7832 (
            .O(N__34581),
            .I(N__34539));
    Span4Mux_v I__7831 (
            .O(N__34578),
            .I(N__34536));
    Span4Mux_v I__7830 (
            .O(N__34575),
            .I(N__34531));
    LocalMux I__7829 (
            .O(N__34572),
            .I(N__34531));
    LocalMux I__7828 (
            .O(N__34569),
            .I(N__34526));
    LocalMux I__7827 (
            .O(N__34566),
            .I(N__34526));
    LocalMux I__7826 (
            .O(N__34563),
            .I(N__34521));
    LocalMux I__7825 (
            .O(N__34556),
            .I(N__34521));
    InMux I__7824 (
            .O(N__34555),
            .I(N__34518));
    Span4Mux_v I__7823 (
            .O(N__34550),
            .I(N__34515));
    Span4Mux_v I__7822 (
            .O(N__34547),
            .I(N__34508));
    Span4Mux_s2_h I__7821 (
            .O(N__34544),
            .I(N__34508));
    Span4Mux_v I__7820 (
            .O(N__34539),
            .I(N__34508));
    Span4Mux_s2_v I__7819 (
            .O(N__34536),
            .I(N__34503));
    Span4Mux_v I__7818 (
            .O(N__34531),
            .I(N__34503));
    Span4Mux_v I__7817 (
            .O(N__34526),
            .I(N__34496));
    Span4Mux_h I__7816 (
            .O(N__34521),
            .I(N__34496));
    LocalMux I__7815 (
            .O(N__34518),
            .I(N__34496));
    Span4Mux_h I__7814 (
            .O(N__34515),
            .I(N__34488));
    Span4Mux_v I__7813 (
            .O(N__34508),
            .I(N__34488));
    Span4Mux_h I__7812 (
            .O(N__34503),
            .I(N__34483));
    Span4Mux_v I__7811 (
            .O(N__34496),
            .I(N__34483));
    InMux I__7810 (
            .O(N__34495),
            .I(N__34480));
    InMux I__7809 (
            .O(N__34494),
            .I(N__34477));
    InMux I__7808 (
            .O(N__34493),
            .I(N__34474));
    IoSpan4Mux I__7807 (
            .O(N__34488),
            .I(N__34469));
    IoSpan4Mux I__7806 (
            .O(N__34483),
            .I(N__34469));
    LocalMux I__7805 (
            .O(N__34480),
            .I(N__34462));
    LocalMux I__7804 (
            .O(N__34477),
            .I(N__34462));
    LocalMux I__7803 (
            .O(N__34474),
            .I(N__34462));
    Odrv4 I__7802 (
            .O(N__34469),
            .I(slp_s3n));
    Odrv12 I__7801 (
            .O(N__34462),
            .I(slp_s3n));
    InMux I__7800 (
            .O(N__34457),
            .I(N__34449));
    CascadeMux I__7799 (
            .O(N__34456),
            .I(N__34446));
    InMux I__7798 (
            .O(N__34455),
            .I(N__34442));
    CascadeMux I__7797 (
            .O(N__34454),
            .I(N__34439));
    InMux I__7796 (
            .O(N__34453),
            .I(N__34434));
    InMux I__7795 (
            .O(N__34452),
            .I(N__34434));
    LocalMux I__7794 (
            .O(N__34449),
            .I(N__34429));
    InMux I__7793 (
            .O(N__34446),
            .I(N__34426));
    CascadeMux I__7792 (
            .O(N__34445),
            .I(N__34423));
    LocalMux I__7791 (
            .O(N__34442),
            .I(N__34418));
    InMux I__7790 (
            .O(N__34439),
            .I(N__34415));
    LocalMux I__7789 (
            .O(N__34434),
            .I(N__34412));
    InMux I__7788 (
            .O(N__34433),
            .I(N__34409));
    InMux I__7787 (
            .O(N__34432),
            .I(N__34406));
    Span4Mux_v I__7786 (
            .O(N__34429),
            .I(N__34400));
    LocalMux I__7785 (
            .O(N__34426),
            .I(N__34400));
    InMux I__7784 (
            .O(N__34423),
            .I(N__34397));
    InMux I__7783 (
            .O(N__34422),
            .I(N__34392));
    InMux I__7782 (
            .O(N__34421),
            .I(N__34389));
    Span4Mux_v I__7781 (
            .O(N__34418),
            .I(N__34385));
    LocalMux I__7780 (
            .O(N__34415),
            .I(N__34382));
    Span4Mux_h I__7779 (
            .O(N__34412),
            .I(N__34375));
    LocalMux I__7778 (
            .O(N__34409),
            .I(N__34375));
    LocalMux I__7777 (
            .O(N__34406),
            .I(N__34375));
    InMux I__7776 (
            .O(N__34405),
            .I(N__34372));
    Span4Mux_h I__7775 (
            .O(N__34400),
            .I(N__34369));
    LocalMux I__7774 (
            .O(N__34397),
            .I(N__34366));
    InMux I__7773 (
            .O(N__34396),
            .I(N__34363));
    InMux I__7772 (
            .O(N__34395),
            .I(N__34360));
    LocalMux I__7771 (
            .O(N__34392),
            .I(N__34355));
    LocalMux I__7770 (
            .O(N__34389),
            .I(N__34355));
    InMux I__7769 (
            .O(N__34388),
            .I(N__34352));
    Span4Mux_h I__7768 (
            .O(N__34385),
            .I(N__34343));
    Span4Mux_v I__7767 (
            .O(N__34382),
            .I(N__34343));
    Span4Mux_v I__7766 (
            .O(N__34375),
            .I(N__34343));
    LocalMux I__7765 (
            .O(N__34372),
            .I(N__34343));
    Sp12to4 I__7764 (
            .O(N__34369),
            .I(N__34330));
    Sp12to4 I__7763 (
            .O(N__34366),
            .I(N__34330));
    LocalMux I__7762 (
            .O(N__34363),
            .I(N__34330));
    LocalMux I__7761 (
            .O(N__34360),
            .I(N__34330));
    Sp12to4 I__7760 (
            .O(N__34355),
            .I(N__34330));
    LocalMux I__7759 (
            .O(N__34352),
            .I(N__34330));
    Span4Mux_v I__7758 (
            .O(N__34343),
            .I(N__34327));
    Span12Mux_v I__7757 (
            .O(N__34330),
            .I(N__34324));
    Odrv4 I__7756 (
            .O(N__34327),
            .I(gpio_fpga_soc_4));
    Odrv12 I__7755 (
            .O(N__34324),
            .I(gpio_fpga_soc_4));
    IoInMux I__7754 (
            .O(N__34319),
            .I(N__34316));
    LocalMux I__7753 (
            .O(N__34316),
            .I(N__34313));
    IoSpan4Mux I__7752 (
            .O(N__34313),
            .I(N__34308));
    CascadeMux I__7751 (
            .O(N__34312),
            .I(N__34305));
    CascadeMux I__7750 (
            .O(N__34311),
            .I(N__34302));
    IoSpan4Mux I__7749 (
            .O(N__34308),
            .I(N__34297));
    InMux I__7748 (
            .O(N__34305),
            .I(N__34294));
    InMux I__7747 (
            .O(N__34302),
            .I(N__34291));
    InMux I__7746 (
            .O(N__34301),
            .I(N__34281));
    CascadeMux I__7745 (
            .O(N__34300),
            .I(N__34278));
    Span4Mux_s3_v I__7744 (
            .O(N__34297),
            .I(N__34270));
    LocalMux I__7743 (
            .O(N__34294),
            .I(N__34270));
    LocalMux I__7742 (
            .O(N__34291),
            .I(N__34270));
    InMux I__7741 (
            .O(N__34290),
            .I(N__34265));
    InMux I__7740 (
            .O(N__34289),
            .I(N__34265));
    CascadeMux I__7739 (
            .O(N__34288),
            .I(N__34262));
    CascadeMux I__7738 (
            .O(N__34287),
            .I(N__34259));
    CascadeMux I__7737 (
            .O(N__34286),
            .I(N__34256));
    CascadeMux I__7736 (
            .O(N__34285),
            .I(N__34253));
    InMux I__7735 (
            .O(N__34284),
            .I(N__34245));
    LocalMux I__7734 (
            .O(N__34281),
            .I(N__34242));
    InMux I__7733 (
            .O(N__34278),
            .I(N__34238));
    InMux I__7732 (
            .O(N__34277),
            .I(N__34235));
    Span4Mux_v I__7731 (
            .O(N__34270),
            .I(N__34230));
    LocalMux I__7730 (
            .O(N__34265),
            .I(N__34230));
    InMux I__7729 (
            .O(N__34262),
            .I(N__34225));
    InMux I__7728 (
            .O(N__34259),
            .I(N__34225));
    InMux I__7727 (
            .O(N__34256),
            .I(N__34222));
    InMux I__7726 (
            .O(N__34253),
            .I(N__34216));
    InMux I__7725 (
            .O(N__34252),
            .I(N__34211));
    InMux I__7724 (
            .O(N__34251),
            .I(N__34211));
    InMux I__7723 (
            .O(N__34250),
            .I(N__34208));
    InMux I__7722 (
            .O(N__34249),
            .I(N__34205));
    InMux I__7721 (
            .O(N__34248),
            .I(N__34202));
    LocalMux I__7720 (
            .O(N__34245),
            .I(N__34197));
    Span4Mux_v I__7719 (
            .O(N__34242),
            .I(N__34194));
    InMux I__7718 (
            .O(N__34241),
            .I(N__34191));
    LocalMux I__7717 (
            .O(N__34238),
            .I(N__34186));
    LocalMux I__7716 (
            .O(N__34235),
            .I(N__34186));
    Sp12to4 I__7715 (
            .O(N__34230),
            .I(N__34183));
    LocalMux I__7714 (
            .O(N__34225),
            .I(N__34178));
    LocalMux I__7713 (
            .O(N__34222),
            .I(N__34175));
    InMux I__7712 (
            .O(N__34221),
            .I(N__34172));
    InMux I__7711 (
            .O(N__34220),
            .I(N__34169));
    InMux I__7710 (
            .O(N__34219),
            .I(N__34166));
    LocalMux I__7709 (
            .O(N__34216),
            .I(N__34163));
    LocalMux I__7708 (
            .O(N__34211),
            .I(N__34160));
    LocalMux I__7707 (
            .O(N__34208),
            .I(N__34155));
    LocalMux I__7706 (
            .O(N__34205),
            .I(N__34155));
    LocalMux I__7705 (
            .O(N__34202),
            .I(N__34152));
    InMux I__7704 (
            .O(N__34201),
            .I(N__34149));
    InMux I__7703 (
            .O(N__34200),
            .I(N__34146));
    Span12Mux_s8_v I__7702 (
            .O(N__34197),
            .I(N__34143));
    Sp12to4 I__7701 (
            .O(N__34194),
            .I(N__34134));
    LocalMux I__7700 (
            .O(N__34191),
            .I(N__34134));
    Span12Mux_s8_v I__7699 (
            .O(N__34186),
            .I(N__34134));
    Span12Mux_s7_v I__7698 (
            .O(N__34183),
            .I(N__34134));
    InMux I__7697 (
            .O(N__34182),
            .I(N__34131));
    InMux I__7696 (
            .O(N__34181),
            .I(N__34128));
    Span4Mux_h I__7695 (
            .O(N__34178),
            .I(N__34117));
    Span4Mux_h I__7694 (
            .O(N__34175),
            .I(N__34117));
    LocalMux I__7693 (
            .O(N__34172),
            .I(N__34117));
    LocalMux I__7692 (
            .O(N__34169),
            .I(N__34117));
    LocalMux I__7691 (
            .O(N__34166),
            .I(N__34117));
    Span4Mux_h I__7690 (
            .O(N__34163),
            .I(N__34110));
    Span4Mux_h I__7689 (
            .O(N__34160),
            .I(N__34110));
    Span4Mux_s3_h I__7688 (
            .O(N__34155),
            .I(N__34110));
    Span4Mux_s2_h I__7687 (
            .O(N__34152),
            .I(N__34107));
    LocalMux I__7686 (
            .O(N__34149),
            .I(N__34102));
    LocalMux I__7685 (
            .O(N__34146),
            .I(N__34102));
    Odrv12 I__7684 (
            .O(N__34143),
            .I(rsmrstn));
    Odrv12 I__7683 (
            .O(N__34134),
            .I(rsmrstn));
    LocalMux I__7682 (
            .O(N__34131),
            .I(rsmrstn));
    LocalMux I__7681 (
            .O(N__34128),
            .I(rsmrstn));
    Odrv4 I__7680 (
            .O(N__34117),
            .I(rsmrstn));
    Odrv4 I__7679 (
            .O(N__34110),
            .I(rsmrstn));
    Odrv4 I__7678 (
            .O(N__34107),
            .I(rsmrstn));
    Odrv12 I__7677 (
            .O(N__34102),
            .I(rsmrstn));
    InMux I__7676 (
            .O(N__34085),
            .I(N__34082));
    LocalMux I__7675 (
            .O(N__34082),
            .I(N__34079));
    Span4Mux_v I__7674 (
            .O(N__34079),
            .I(N__34075));
    InMux I__7673 (
            .O(N__34078),
            .I(N__34072));
    Odrv4 I__7672 (
            .O(N__34075),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0 ));
    LocalMux I__7671 (
            .O(N__34072),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0 ));
    InMux I__7670 (
            .O(N__34067),
            .I(N__34053));
    InMux I__7669 (
            .O(N__34066),
            .I(N__34049));
    InMux I__7668 (
            .O(N__34065),
            .I(N__34045));
    InMux I__7667 (
            .O(N__34064),
            .I(N__34042));
    InMux I__7666 (
            .O(N__34063),
            .I(N__34035));
    InMux I__7665 (
            .O(N__34062),
            .I(N__34035));
    InMux I__7664 (
            .O(N__34061),
            .I(N__34032));
    InMux I__7663 (
            .O(N__34060),
            .I(N__34027));
    InMux I__7662 (
            .O(N__34059),
            .I(N__34027));
    InMux I__7661 (
            .O(N__34058),
            .I(N__34020));
    InMux I__7660 (
            .O(N__34057),
            .I(N__34020));
    InMux I__7659 (
            .O(N__34056),
            .I(N__34020));
    LocalMux I__7658 (
            .O(N__34053),
            .I(N__34017));
    InMux I__7657 (
            .O(N__34052),
            .I(N__34011));
    LocalMux I__7656 (
            .O(N__34049),
            .I(N__34008));
    InMux I__7655 (
            .O(N__34048),
            .I(N__34005));
    LocalMux I__7654 (
            .O(N__34045),
            .I(N__34000));
    LocalMux I__7653 (
            .O(N__34042),
            .I(N__34000));
    InMux I__7652 (
            .O(N__34041),
            .I(N__33995));
    InMux I__7651 (
            .O(N__34040),
            .I(N__33995));
    LocalMux I__7650 (
            .O(N__34035),
            .I(N__33990));
    LocalMux I__7649 (
            .O(N__34032),
            .I(N__33990));
    LocalMux I__7648 (
            .O(N__34027),
            .I(N__33985));
    LocalMux I__7647 (
            .O(N__34020),
            .I(N__33985));
    Span12Mux_s2_h I__7646 (
            .O(N__34017),
            .I(N__33982));
    InMux I__7645 (
            .O(N__34016),
            .I(N__33979));
    InMux I__7644 (
            .O(N__34015),
            .I(N__33976));
    InMux I__7643 (
            .O(N__34014),
            .I(N__33973));
    LocalMux I__7642 (
            .O(N__34011),
            .I(N__33970));
    Span4Mux_h I__7641 (
            .O(N__34008),
            .I(N__33961));
    LocalMux I__7640 (
            .O(N__34005),
            .I(N__33961));
    Span4Mux_s3_h I__7639 (
            .O(N__34000),
            .I(N__33961));
    LocalMux I__7638 (
            .O(N__33995),
            .I(N__33961));
    Span4Mux_s2_h I__7637 (
            .O(N__33990),
            .I(N__33958));
    Span4Mux_s2_h I__7636 (
            .O(N__33985),
            .I(N__33955));
    Odrv12 I__7635 (
            .O(N__33982),
            .I(\b2v_inst11.N_2946_i ));
    LocalMux I__7634 (
            .O(N__33979),
            .I(\b2v_inst11.N_2946_i ));
    LocalMux I__7633 (
            .O(N__33976),
            .I(\b2v_inst11.N_2946_i ));
    LocalMux I__7632 (
            .O(N__33973),
            .I(\b2v_inst11.N_2946_i ));
    Odrv12 I__7631 (
            .O(N__33970),
            .I(\b2v_inst11.N_2946_i ));
    Odrv4 I__7630 (
            .O(N__33961),
            .I(\b2v_inst11.N_2946_i ));
    Odrv4 I__7629 (
            .O(N__33958),
            .I(\b2v_inst11.N_2946_i ));
    Odrv4 I__7628 (
            .O(N__33955),
            .I(\b2v_inst11.N_2946_i ));
    CascadeMux I__7627 (
            .O(N__33938),
            .I(N__33934));
    InMux I__7626 (
            .O(N__33937),
            .I(N__33930));
    InMux I__7625 (
            .O(N__33934),
            .I(N__33925));
    InMux I__7624 (
            .O(N__33933),
            .I(N__33922));
    LocalMux I__7623 (
            .O(N__33930),
            .I(N__33914));
    InMux I__7622 (
            .O(N__33929),
            .I(N__33909));
    InMux I__7621 (
            .O(N__33928),
            .I(N__33909));
    LocalMux I__7620 (
            .O(N__33925),
            .I(N__33904));
    LocalMux I__7619 (
            .O(N__33922),
            .I(N__33904));
    InMux I__7618 (
            .O(N__33921),
            .I(N__33899));
    InMux I__7617 (
            .O(N__33920),
            .I(N__33899));
    InMux I__7616 (
            .O(N__33919),
            .I(N__33895));
    InMux I__7615 (
            .O(N__33918),
            .I(N__33892));
    InMux I__7614 (
            .O(N__33917),
            .I(N__33888));
    Span4Mux_h I__7613 (
            .O(N__33914),
            .I(N__33874));
    LocalMux I__7612 (
            .O(N__33909),
            .I(N__33874));
    Span4Mux_h I__7611 (
            .O(N__33904),
            .I(N__33874));
    LocalMux I__7610 (
            .O(N__33899),
            .I(N__33871));
    InMux I__7609 (
            .O(N__33898),
            .I(N__33868));
    LocalMux I__7608 (
            .O(N__33895),
            .I(N__33861));
    LocalMux I__7607 (
            .O(N__33892),
            .I(N__33861));
    InMux I__7606 (
            .O(N__33891),
            .I(N__33858));
    LocalMux I__7605 (
            .O(N__33888),
            .I(N__33855));
    CascadeMux I__7604 (
            .O(N__33887),
            .I(N__33851));
    InMux I__7603 (
            .O(N__33886),
            .I(N__33837));
    InMux I__7602 (
            .O(N__33885),
            .I(N__33837));
    InMux I__7601 (
            .O(N__33884),
            .I(N__33832));
    InMux I__7600 (
            .O(N__33883),
            .I(N__33832));
    InMux I__7599 (
            .O(N__33882),
            .I(N__33827));
    InMux I__7598 (
            .O(N__33881),
            .I(N__33827));
    Span4Mux_v I__7597 (
            .O(N__33874),
            .I(N__33824));
    Span4Mux_v I__7596 (
            .O(N__33871),
            .I(N__33819));
    LocalMux I__7595 (
            .O(N__33868),
            .I(N__33819));
    InMux I__7594 (
            .O(N__33867),
            .I(N__33814));
    InMux I__7593 (
            .O(N__33866),
            .I(N__33814));
    Span4Mux_v I__7592 (
            .O(N__33861),
            .I(N__33811));
    LocalMux I__7591 (
            .O(N__33858),
            .I(N__33808));
    Span4Mux_v I__7590 (
            .O(N__33855),
            .I(N__33805));
    InMux I__7589 (
            .O(N__33854),
            .I(N__33796));
    InMux I__7588 (
            .O(N__33851),
            .I(N__33796));
    InMux I__7587 (
            .O(N__33850),
            .I(N__33796));
    InMux I__7586 (
            .O(N__33849),
            .I(N__33796));
    InMux I__7585 (
            .O(N__33848),
            .I(N__33793));
    InMux I__7584 (
            .O(N__33847),
            .I(N__33786));
    InMux I__7583 (
            .O(N__33846),
            .I(N__33786));
    InMux I__7582 (
            .O(N__33845),
            .I(N__33786));
    InMux I__7581 (
            .O(N__33844),
            .I(N__33779));
    InMux I__7580 (
            .O(N__33843),
            .I(N__33779));
    InMux I__7579 (
            .O(N__33842),
            .I(N__33779));
    LocalMux I__7578 (
            .O(N__33837),
            .I(N__33776));
    LocalMux I__7577 (
            .O(N__33832),
            .I(N__33773));
    LocalMux I__7576 (
            .O(N__33827),
            .I(N__33764));
    Span4Mux_h I__7575 (
            .O(N__33824),
            .I(N__33764));
    Span4Mux_h I__7574 (
            .O(N__33819),
            .I(N__33764));
    LocalMux I__7573 (
            .O(N__33814),
            .I(N__33764));
    Span4Mux_h I__7572 (
            .O(N__33811),
            .I(N__33759));
    Span4Mux_v I__7571 (
            .O(N__33808),
            .I(N__33759));
    Span4Mux_h I__7570 (
            .O(N__33805),
            .I(N__33754));
    LocalMux I__7569 (
            .O(N__33796),
            .I(N__33754));
    LocalMux I__7568 (
            .O(N__33793),
            .I(N__33745));
    LocalMux I__7567 (
            .O(N__33786),
            .I(N__33745));
    LocalMux I__7566 (
            .O(N__33779),
            .I(N__33745));
    Span12Mux_s5_v I__7565 (
            .O(N__33776),
            .I(N__33745));
    Span4Mux_v I__7564 (
            .O(N__33773),
            .I(N__33740));
    Span4Mux_v I__7563 (
            .O(N__33764),
            .I(N__33740));
    Odrv4 I__7562 (
            .O(N__33759),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ));
    Odrv4 I__7561 (
            .O(N__33754),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ));
    Odrv12 I__7560 (
            .O(N__33745),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ));
    Odrv4 I__7559 (
            .O(N__33740),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ));
    CascadeMux I__7558 (
            .O(N__33731),
            .I(N__33727));
    InMux I__7557 (
            .O(N__33730),
            .I(N__33723));
    InMux I__7556 (
            .O(N__33727),
            .I(N__33720));
    InMux I__7555 (
            .O(N__33726),
            .I(N__33717));
    LocalMux I__7554 (
            .O(N__33723),
            .I(N__33711));
    LocalMux I__7553 (
            .O(N__33720),
            .I(N__33711));
    LocalMux I__7552 (
            .O(N__33717),
            .I(N__33708));
    InMux I__7551 (
            .O(N__33716),
            .I(N__33704));
    Span4Mux_s0_h I__7550 (
            .O(N__33711),
            .I(N__33699));
    Span4Mux_v I__7549 (
            .O(N__33708),
            .I(N__33699));
    InMux I__7548 (
            .O(N__33707),
            .I(N__33696));
    LocalMux I__7547 (
            .O(N__33704),
            .I(N__33693));
    Span4Mux_h I__7546 (
            .O(N__33699),
            .I(N__33688));
    LocalMux I__7545 (
            .O(N__33696),
            .I(N__33688));
    Span4Mux_v I__7544 (
            .O(N__33693),
            .I(N__33685));
    Span4Mux_h I__7543 (
            .O(N__33688),
            .I(N__33682));
    Span4Mux_h I__7542 (
            .O(N__33685),
            .I(N__33679));
    Odrv4 I__7541 (
            .O(N__33682),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_5 ));
    Odrv4 I__7540 (
            .O(N__33679),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_5 ));
    InMux I__7539 (
            .O(N__33674),
            .I(N__33671));
    LocalMux I__7538 (
            .O(N__33671),
            .I(N__33668));
    Odrv4 I__7537 (
            .O(N__33668),
            .I(\b2v_inst11.g0_1_1 ));
    InMux I__7536 (
            .O(N__33665),
            .I(N__33662));
    LocalMux I__7535 (
            .O(N__33662),
            .I(N__33659));
    Span4Mux_v I__7534 (
            .O(N__33659),
            .I(N__33656));
    Odrv4 I__7533 (
            .O(N__33656),
            .I(vddq_ok));
    InMux I__7532 (
            .O(N__33653),
            .I(N__33650));
    LocalMux I__7531 (
            .O(N__33650),
            .I(N__33647));
    Span4Mux_h I__7530 (
            .O(N__33647),
            .I(N__33643));
    InMux I__7529 (
            .O(N__33646),
            .I(N__33640));
    Span4Mux_v I__7528 (
            .O(N__33643),
            .I(N__33634));
    LocalMux I__7527 (
            .O(N__33640),
            .I(N__33634));
    InMux I__7526 (
            .O(N__33639),
            .I(N__33629));
    Span4Mux_v I__7525 (
            .O(N__33634),
            .I(N__33626));
    InMux I__7524 (
            .O(N__33633),
            .I(N__33623));
    CascadeMux I__7523 (
            .O(N__33632),
            .I(N__33619));
    LocalMux I__7522 (
            .O(N__33629),
            .I(N__33614));
    Span4Mux_h I__7521 (
            .O(N__33626),
            .I(N__33609));
    LocalMux I__7520 (
            .O(N__33623),
            .I(N__33609));
    InMux I__7519 (
            .O(N__33622),
            .I(N__33606));
    InMux I__7518 (
            .O(N__33619),
            .I(N__33603));
    InMux I__7517 (
            .O(N__33618),
            .I(N__33600));
    InMux I__7516 (
            .O(N__33617),
            .I(N__33597));
    Span12Mux_s3_h I__7515 (
            .O(N__33614),
            .I(N__33594));
    Sp12to4 I__7514 (
            .O(N__33609),
            .I(N__33583));
    LocalMux I__7513 (
            .O(N__33606),
            .I(N__33583));
    LocalMux I__7512 (
            .O(N__33603),
            .I(N__33583));
    LocalMux I__7511 (
            .O(N__33600),
            .I(N__33583));
    LocalMux I__7510 (
            .O(N__33597),
            .I(N__33583));
    Odrv12 I__7509 (
            .O(N__33594),
            .I(VCCST_EN_i_0_o3_0));
    Odrv12 I__7508 (
            .O(N__33583),
            .I(VCCST_EN_i_0_o3_0));
    InMux I__7507 (
            .O(N__33578),
            .I(N__33573));
    InMux I__7506 (
            .O(N__33577),
            .I(N__33570));
    InMux I__7505 (
            .O(N__33576),
            .I(N__33567));
    LocalMux I__7504 (
            .O(N__33573),
            .I(N__33562));
    LocalMux I__7503 (
            .O(N__33570),
            .I(N__33562));
    LocalMux I__7502 (
            .O(N__33567),
            .I(N__33559));
    Span4Mux_h I__7501 (
            .O(N__33562),
            .I(N__33556));
    Sp12to4 I__7500 (
            .O(N__33559),
            .I(N__33553));
    Span4Mux_h I__7499 (
            .O(N__33556),
            .I(N__33550));
    Span12Mux_s10_v I__7498 (
            .O(N__33553),
            .I(N__33547));
    Span4Mux_v I__7497 (
            .O(N__33550),
            .I(N__33544));
    Odrv12 I__7496 (
            .O(N__33547),
            .I(\b2v_inst16.N_208_0 ));
    Odrv4 I__7495 (
            .O(N__33544),
            .I(\b2v_inst16.N_208_0 ));
    InMux I__7494 (
            .O(N__33539),
            .I(N__33536));
    LocalMux I__7493 (
            .O(N__33536),
            .I(\b2v_inst11.count_off_1_1 ));
    CascadeMux I__7492 (
            .O(N__33533),
            .I(\b2v_inst11.g0_13_1_cascade_ ));
    CascadeMux I__7491 (
            .O(N__33530),
            .I(\b2v_inst11.N_4690_0_0_cascade_ ));
    InMux I__7490 (
            .O(N__33527),
            .I(N__33524));
    LocalMux I__7489 (
            .O(N__33524),
            .I(\b2v_inst11.N_19_0 ));
    InMux I__7488 (
            .O(N__33521),
            .I(N__33518));
    LocalMux I__7487 (
            .O(N__33518),
            .I(\b2v_inst11.N_19_1 ));
    CascadeMux I__7486 (
            .O(N__33515),
            .I(N__33510));
    CascadeMux I__7485 (
            .O(N__33514),
            .I(N__33505));
    CascadeMux I__7484 (
            .O(N__33513),
            .I(N__33502));
    InMux I__7483 (
            .O(N__33510),
            .I(N__33495));
    InMux I__7482 (
            .O(N__33509),
            .I(N__33495));
    InMux I__7481 (
            .O(N__33508),
            .I(N__33492));
    InMux I__7480 (
            .O(N__33505),
            .I(N__33489));
    InMux I__7479 (
            .O(N__33502),
            .I(N__33484));
    InMux I__7478 (
            .O(N__33501),
            .I(N__33484));
    InMux I__7477 (
            .O(N__33500),
            .I(N__33481));
    LocalMux I__7476 (
            .O(N__33495),
            .I(N__33478));
    LocalMux I__7475 (
            .O(N__33492),
            .I(N__33474));
    LocalMux I__7474 (
            .O(N__33489),
            .I(N__33471));
    LocalMux I__7473 (
            .O(N__33484),
            .I(N__33468));
    LocalMux I__7472 (
            .O(N__33481),
            .I(N__33464));
    Span4Mux_s2_h I__7471 (
            .O(N__33478),
            .I(N__33461));
    InMux I__7470 (
            .O(N__33477),
            .I(N__33458));
    Span4Mux_s3_h I__7469 (
            .O(N__33474),
            .I(N__33451));
    Span4Mux_s3_h I__7468 (
            .O(N__33471),
            .I(N__33451));
    Span4Mux_v I__7467 (
            .O(N__33468),
            .I(N__33451));
    InMux I__7466 (
            .O(N__33467),
            .I(N__33448));
    Odrv12 I__7465 (
            .O(N__33464),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__7464 (
            .O(N__33461),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    LocalMux I__7463 (
            .O(N__33458),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__7462 (
            .O(N__33451),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    LocalMux I__7461 (
            .O(N__33448),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    InMux I__7460 (
            .O(N__33437),
            .I(N__33434));
    LocalMux I__7459 (
            .O(N__33434),
            .I(\b2v_inst11.un1_dutycycle_172_m0 ));
    InMux I__7458 (
            .O(N__33431),
            .I(N__33428));
    LocalMux I__7457 (
            .O(N__33428),
            .I(N__33425));
    Span12Mux_s10_v I__7456 (
            .O(N__33425),
            .I(N__33422));
    Odrv12 I__7455 (
            .O(N__33422),
            .I(\b2v_inst11.g3_3 ));
    InMux I__7454 (
            .O(N__33419),
            .I(N__33412));
    InMux I__7453 (
            .O(N__33418),
            .I(N__33408));
    InMux I__7452 (
            .O(N__33417),
            .I(N__33403));
    InMux I__7451 (
            .O(N__33416),
            .I(N__33398));
    InMux I__7450 (
            .O(N__33415),
            .I(N__33398));
    LocalMux I__7449 (
            .O(N__33412),
            .I(N__33395));
    InMux I__7448 (
            .O(N__33411),
            .I(N__33392));
    LocalMux I__7447 (
            .O(N__33408),
            .I(N__33389));
    InMux I__7446 (
            .O(N__33407),
            .I(N__33386));
    InMux I__7445 (
            .O(N__33406),
            .I(N__33381));
    LocalMux I__7444 (
            .O(N__33403),
            .I(N__33372));
    LocalMux I__7443 (
            .O(N__33398),
            .I(N__33372));
    Span4Mux_v I__7442 (
            .O(N__33395),
            .I(N__33369));
    LocalMux I__7441 (
            .O(N__33392),
            .I(N__33366));
    Span4Mux_v I__7440 (
            .O(N__33389),
            .I(N__33361));
    LocalMux I__7439 (
            .O(N__33386),
            .I(N__33361));
    InMux I__7438 (
            .O(N__33385),
            .I(N__33356));
    InMux I__7437 (
            .O(N__33384),
            .I(N__33356));
    LocalMux I__7436 (
            .O(N__33381),
            .I(N__33353));
    InMux I__7435 (
            .O(N__33380),
            .I(N__33348));
    InMux I__7434 (
            .O(N__33379),
            .I(N__33348));
    InMux I__7433 (
            .O(N__33378),
            .I(N__33345));
    InMux I__7432 (
            .O(N__33377),
            .I(N__33342));
    Span12Mux_s8_v I__7431 (
            .O(N__33372),
            .I(N__33339));
    Span4Mux_v I__7430 (
            .O(N__33369),
            .I(N__33330));
    Span4Mux_h I__7429 (
            .O(N__33366),
            .I(N__33330));
    Span4Mux_v I__7428 (
            .O(N__33361),
            .I(N__33330));
    LocalMux I__7427 (
            .O(N__33356),
            .I(N__33330));
    Span4Mux_h I__7426 (
            .O(N__33353),
            .I(N__33327));
    LocalMux I__7425 (
            .O(N__33348),
            .I(\b2v_inst11.N_172 ));
    LocalMux I__7424 (
            .O(N__33345),
            .I(\b2v_inst11.N_172 ));
    LocalMux I__7423 (
            .O(N__33342),
            .I(\b2v_inst11.N_172 ));
    Odrv12 I__7422 (
            .O(N__33339),
            .I(\b2v_inst11.N_172 ));
    Odrv4 I__7421 (
            .O(N__33330),
            .I(\b2v_inst11.N_172 ));
    Odrv4 I__7420 (
            .O(N__33327),
            .I(\b2v_inst11.N_172 ));
    CascadeMux I__7419 (
            .O(N__33314),
            .I(N__33308));
    InMux I__7418 (
            .O(N__33313),
            .I(N__33299));
    InMux I__7417 (
            .O(N__33312),
            .I(N__33299));
    InMux I__7416 (
            .O(N__33311),
            .I(N__33294));
    InMux I__7415 (
            .O(N__33308),
            .I(N__33294));
    InMux I__7414 (
            .O(N__33307),
            .I(N__33288));
    InMux I__7413 (
            .O(N__33306),
            .I(N__33288));
    InMux I__7412 (
            .O(N__33305),
            .I(N__33285));
    InMux I__7411 (
            .O(N__33304),
            .I(N__33282));
    LocalMux I__7410 (
            .O(N__33299),
            .I(N__33276));
    LocalMux I__7409 (
            .O(N__33294),
            .I(N__33273));
    InMux I__7408 (
            .O(N__33293),
            .I(N__33270));
    LocalMux I__7407 (
            .O(N__33288),
            .I(N__33267));
    LocalMux I__7406 (
            .O(N__33285),
            .I(N__33264));
    LocalMux I__7405 (
            .O(N__33282),
            .I(N__33261));
    InMux I__7404 (
            .O(N__33281),
            .I(N__33253));
    InMux I__7403 (
            .O(N__33280),
            .I(N__33253));
    CascadeMux I__7402 (
            .O(N__33279),
            .I(N__33250));
    Span4Mux_s1_h I__7401 (
            .O(N__33276),
            .I(N__33243));
    Span4Mux_s1_h I__7400 (
            .O(N__33273),
            .I(N__33243));
    LocalMux I__7399 (
            .O(N__33270),
            .I(N__33243));
    Span12Mux_s5_h I__7398 (
            .O(N__33267),
            .I(N__33240));
    Span4Mux_v I__7397 (
            .O(N__33264),
            .I(N__33235));
    Span4Mux_v I__7396 (
            .O(N__33261),
            .I(N__33235));
    InMux I__7395 (
            .O(N__33260),
            .I(N__33228));
    InMux I__7394 (
            .O(N__33259),
            .I(N__33228));
    InMux I__7393 (
            .O(N__33258),
            .I(N__33228));
    LocalMux I__7392 (
            .O(N__33253),
            .I(N__33225));
    InMux I__7391 (
            .O(N__33250),
            .I(N__33222));
    Span4Mux_h I__7390 (
            .O(N__33243),
            .I(N__33219));
    Odrv12 I__7389 (
            .O(N__33240),
            .I(\b2v_inst11.N_200_i ));
    Odrv4 I__7388 (
            .O(N__33235),
            .I(\b2v_inst11.N_200_i ));
    LocalMux I__7387 (
            .O(N__33228),
            .I(\b2v_inst11.N_200_i ));
    Odrv4 I__7386 (
            .O(N__33225),
            .I(\b2v_inst11.N_200_i ));
    LocalMux I__7385 (
            .O(N__33222),
            .I(\b2v_inst11.N_200_i ));
    Odrv4 I__7384 (
            .O(N__33219),
            .I(\b2v_inst11.N_200_i ));
    InMux I__7383 (
            .O(N__33206),
            .I(N__33200));
    InMux I__7382 (
            .O(N__33205),
            .I(N__33200));
    LocalMux I__7381 (
            .O(N__33200),
            .I(\b2v_inst11.N_3099_0_0 ));
    InMux I__7380 (
            .O(N__33197),
            .I(N__33193));
    CascadeMux I__7379 (
            .O(N__33196),
            .I(N__33188));
    LocalMux I__7378 (
            .O(N__33193),
            .I(N__33183));
    InMux I__7377 (
            .O(N__33192),
            .I(N__33178));
    InMux I__7376 (
            .O(N__33191),
            .I(N__33178));
    InMux I__7375 (
            .O(N__33188),
            .I(N__33175));
    InMux I__7374 (
            .O(N__33187),
            .I(N__33171));
    CascadeMux I__7373 (
            .O(N__33186),
            .I(N__33167));
    Span4Mux_s2_v I__7372 (
            .O(N__33183),
            .I(N__33162));
    LocalMux I__7371 (
            .O(N__33178),
            .I(N__33157));
    LocalMux I__7370 (
            .O(N__33175),
            .I(N__33157));
    InMux I__7369 (
            .O(N__33174),
            .I(N__33154));
    LocalMux I__7368 (
            .O(N__33171),
            .I(N__33151));
    InMux I__7367 (
            .O(N__33170),
            .I(N__33147));
    InMux I__7366 (
            .O(N__33167),
            .I(N__33141));
    InMux I__7365 (
            .O(N__33166),
            .I(N__33141));
    InMux I__7364 (
            .O(N__33165),
            .I(N__33138));
    Span4Mux_v I__7363 (
            .O(N__33162),
            .I(N__33131));
    Span4Mux_v I__7362 (
            .O(N__33157),
            .I(N__33131));
    LocalMux I__7361 (
            .O(N__33154),
            .I(N__33131));
    Span4Mux_h I__7360 (
            .O(N__33151),
            .I(N__33128));
    InMux I__7359 (
            .O(N__33150),
            .I(N__33125));
    LocalMux I__7358 (
            .O(N__33147),
            .I(N__33122));
    InMux I__7357 (
            .O(N__33146),
            .I(N__33119));
    LocalMux I__7356 (
            .O(N__33141),
            .I(N__33114));
    LocalMux I__7355 (
            .O(N__33138),
            .I(N__33114));
    Span4Mux_h I__7354 (
            .O(N__33131),
            .I(N__33111));
    Odrv4 I__7353 (
            .O(N__33128),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    LocalMux I__7352 (
            .O(N__33125),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    Odrv4 I__7351 (
            .O(N__33122),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    LocalMux I__7350 (
            .O(N__33119),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    Odrv12 I__7349 (
            .O(N__33114),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    Odrv4 I__7348 (
            .O(N__33111),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    InMux I__7347 (
            .O(N__33098),
            .I(N__33095));
    LocalMux I__7346 (
            .O(N__33095),
            .I(N__33092));
    Span4Mux_v I__7345 (
            .O(N__33092),
            .I(N__33089));
    Odrv4 I__7344 (
            .O(N__33089),
            .I(\b2v_inst11.N_237 ));
    InMux I__7343 (
            .O(N__33086),
            .I(N__33083));
    LocalMux I__7342 (
            .O(N__33083),
            .I(\b2v_inst11.N_293_0_0 ));
    CascadeMux I__7341 (
            .O(N__33080),
            .I(N__33075));
    InMux I__7340 (
            .O(N__33079),
            .I(N__33071));
    InMux I__7339 (
            .O(N__33078),
            .I(N__33068));
    InMux I__7338 (
            .O(N__33075),
            .I(N__33065));
    CascadeMux I__7337 (
            .O(N__33074),
            .I(N__33062));
    LocalMux I__7336 (
            .O(N__33071),
            .I(N__33059));
    LocalMux I__7335 (
            .O(N__33068),
            .I(N__33056));
    LocalMux I__7334 (
            .O(N__33065),
            .I(N__33053));
    InMux I__7333 (
            .O(N__33062),
            .I(N__33050));
    Span4Mux_h I__7332 (
            .O(N__33059),
            .I(N__33046));
    Span4Mux_v I__7331 (
            .O(N__33056),
            .I(N__33039));
    Span4Mux_s1_h I__7330 (
            .O(N__33053),
            .I(N__33039));
    LocalMux I__7329 (
            .O(N__33050),
            .I(N__33039));
    InMux I__7328 (
            .O(N__33049),
            .I(N__33036));
    Span4Mux_v I__7327 (
            .O(N__33046),
            .I(N__33033));
    Span4Mux_h I__7326 (
            .O(N__33039),
            .I(N__33028));
    LocalMux I__7325 (
            .O(N__33036),
            .I(N__33028));
    Odrv4 I__7324 (
            .O(N__33033),
            .I(\b2v_inst11.count_clk_RNIZ0Z_6 ));
    Odrv4 I__7323 (
            .O(N__33028),
            .I(\b2v_inst11.count_clk_RNIZ0Z_6 ));
    CascadeMux I__7322 (
            .O(N__33023),
            .I(N__33020));
    InMux I__7321 (
            .O(N__33020),
            .I(N__33014));
    InMux I__7320 (
            .O(N__33019),
            .I(N__33014));
    LocalMux I__7319 (
            .O(N__33014),
            .I(\b2v_inst11.g2_1_0 ));
    InMux I__7318 (
            .O(N__33011),
            .I(N__33008));
    LocalMux I__7317 (
            .O(N__33008),
            .I(v5s_ok));
    CascadeMux I__7316 (
            .O(N__33005),
            .I(N__33002));
    InMux I__7315 (
            .O(N__33002),
            .I(N__32999));
    LocalMux I__7314 (
            .O(N__32999),
            .I(N__32996));
    Span12Mux_v I__7313 (
            .O(N__32996),
            .I(N__32993));
    Odrv12 I__7312 (
            .O(N__32993),
            .I(v33s_ok));
    InMux I__7311 (
            .O(N__32990),
            .I(N__32983));
    InMux I__7310 (
            .O(N__32989),
            .I(N__32976));
    InMux I__7309 (
            .O(N__32988),
            .I(N__32976));
    InMux I__7308 (
            .O(N__32987),
            .I(N__32976));
    InMux I__7307 (
            .O(N__32986),
            .I(N__32973));
    LocalMux I__7306 (
            .O(N__32983),
            .I(N__32965));
    LocalMux I__7305 (
            .O(N__32976),
            .I(N__32965));
    LocalMux I__7304 (
            .O(N__32973),
            .I(N__32965));
    InMux I__7303 (
            .O(N__32972),
            .I(N__32962));
    Span4Mux_v I__7302 (
            .O(N__32965),
            .I(N__32959));
    LocalMux I__7301 (
            .O(N__32962),
            .I(N__32956));
    Odrv4 I__7300 (
            .O(N__32959),
            .I(SYNTHESIZED_WIRE_8));
    Odrv4 I__7299 (
            .O(N__32956),
            .I(SYNTHESIZED_WIRE_8));
    IoInMux I__7298 (
            .O(N__32951),
            .I(N__32948));
    LocalMux I__7297 (
            .O(N__32948),
            .I(N__32945));
    Span4Mux_s2_v I__7296 (
            .O(N__32945),
            .I(N__32942));
    Sp12to4 I__7295 (
            .O(N__32942),
            .I(N__32939));
    Span12Mux_s11_h I__7294 (
            .O(N__32939),
            .I(N__32935));
    IoInMux I__7293 (
            .O(N__32938),
            .I(N__32932));
    Odrv12 I__7292 (
            .O(N__32935),
            .I(vccinaux_en));
    LocalMux I__7291 (
            .O(N__32932),
            .I(vccinaux_en));
    InMux I__7290 (
            .O(N__32927),
            .I(N__32924));
    LocalMux I__7289 (
            .O(N__32924),
            .I(N__32921));
    Odrv4 I__7288 (
            .O(N__32921),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_0 ));
    CascadeMux I__7287 (
            .O(N__32918),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_0_cascade_ ));
    InMux I__7286 (
            .O(N__32915),
            .I(N__32912));
    LocalMux I__7285 (
            .O(N__32912),
            .I(N__32901));
    CascadeMux I__7284 (
            .O(N__32911),
            .I(N__32898));
    InMux I__7283 (
            .O(N__32910),
            .I(N__32891));
    InMux I__7282 (
            .O(N__32909),
            .I(N__32888));
    InMux I__7281 (
            .O(N__32908),
            .I(N__32881));
    InMux I__7280 (
            .O(N__32907),
            .I(N__32881));
    InMux I__7279 (
            .O(N__32906),
            .I(N__32881));
    InMux I__7278 (
            .O(N__32905),
            .I(N__32876));
    InMux I__7277 (
            .O(N__32904),
            .I(N__32876));
    Span4Mux_v I__7276 (
            .O(N__32901),
            .I(N__32870));
    InMux I__7275 (
            .O(N__32898),
            .I(N__32865));
    InMux I__7274 (
            .O(N__32897),
            .I(N__32865));
    InMux I__7273 (
            .O(N__32896),
            .I(N__32862));
    InMux I__7272 (
            .O(N__32895),
            .I(N__32859));
    InMux I__7271 (
            .O(N__32894),
            .I(N__32856));
    LocalMux I__7270 (
            .O(N__32891),
            .I(N__32847));
    LocalMux I__7269 (
            .O(N__32888),
            .I(N__32847));
    LocalMux I__7268 (
            .O(N__32881),
            .I(N__32847));
    LocalMux I__7267 (
            .O(N__32876),
            .I(N__32847));
    InMux I__7266 (
            .O(N__32875),
            .I(N__32842));
    InMux I__7265 (
            .O(N__32874),
            .I(N__32842));
    InMux I__7264 (
            .O(N__32873),
            .I(N__32839));
    Span4Mux_v I__7263 (
            .O(N__32870),
            .I(N__32836));
    LocalMux I__7262 (
            .O(N__32865),
            .I(N__32833));
    LocalMux I__7261 (
            .O(N__32862),
            .I(N__32828));
    LocalMux I__7260 (
            .O(N__32859),
            .I(N__32828));
    LocalMux I__7259 (
            .O(N__32856),
            .I(N__32825));
    Span4Mux_v I__7258 (
            .O(N__32847),
            .I(N__32820));
    LocalMux I__7257 (
            .O(N__32842),
            .I(N__32817));
    LocalMux I__7256 (
            .O(N__32839),
            .I(N__32814));
    Span4Mux_h I__7255 (
            .O(N__32836),
            .I(N__32808));
    Span4Mux_v I__7254 (
            .O(N__32833),
            .I(N__32808));
    Span4Mux_v I__7253 (
            .O(N__32828),
            .I(N__32803));
    Span4Mux_v I__7252 (
            .O(N__32825),
            .I(N__32803));
    InMux I__7251 (
            .O(N__32824),
            .I(N__32800));
    InMux I__7250 (
            .O(N__32823),
            .I(N__32797));
    Span4Mux_v I__7249 (
            .O(N__32820),
            .I(N__32792));
    Span4Mux_v I__7248 (
            .O(N__32817),
            .I(N__32792));
    Span4Mux_v I__7247 (
            .O(N__32814),
            .I(N__32789));
    InMux I__7246 (
            .O(N__32813),
            .I(N__32786));
    Span4Mux_h I__7245 (
            .O(N__32808),
            .I(N__32783));
    Sp12to4 I__7244 (
            .O(N__32803),
            .I(N__32770));
    LocalMux I__7243 (
            .O(N__32800),
            .I(N__32770));
    LocalMux I__7242 (
            .O(N__32797),
            .I(N__32770));
    Sp12to4 I__7241 (
            .O(N__32792),
            .I(N__32770));
    Sp12to4 I__7240 (
            .O(N__32789),
            .I(N__32770));
    LocalMux I__7239 (
            .O(N__32786),
            .I(N__32770));
    Sp12to4 I__7238 (
            .O(N__32783),
            .I(N__32765));
    Span12Mux_s8_h I__7237 (
            .O(N__32770),
            .I(N__32765));
    Odrv12 I__7236 (
            .O(N__32765),
            .I(slp_s4n));
    InMux I__7235 (
            .O(N__32762),
            .I(N__32756));
    InMux I__7234 (
            .O(N__32761),
            .I(N__32756));
    LocalMux I__7233 (
            .O(N__32756),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_0 ));
    CascadeMux I__7232 (
            .O(N__32753),
            .I(\b2v_inst11.un1_dutycycle_172_m1_ns_1_cascade_ ));
    InMux I__7231 (
            .O(N__32750),
            .I(N__32747));
    LocalMux I__7230 (
            .O(N__32747),
            .I(\b2v_inst11.un1_dutycycle_172_m1 ));
    InMux I__7229 (
            .O(N__32744),
            .I(N__32741));
    LocalMux I__7228 (
            .O(N__32741),
            .I(\b2v_inst11.g0_i_2 ));
    CascadeMux I__7227 (
            .O(N__32738),
            .I(\b2v_inst11.g0_0_0Z0Z_0_cascade_ ));
    InMux I__7226 (
            .O(N__32735),
            .I(N__32732));
    LocalMux I__7225 (
            .O(N__32732),
            .I(\b2v_inst6.count_1_i_a3_7_0 ));
    InMux I__7224 (
            .O(N__32729),
            .I(N__32726));
    LocalMux I__7223 (
            .O(N__32726),
            .I(N__32723));
    Odrv12 I__7222 (
            .O(N__32723),
            .I(\b2v_inst6.count_1_i_a3_1_0 ));
    CascadeMux I__7221 (
            .O(N__32720),
            .I(\b2v_inst6.count_1_i_a3_12_0_cascade_ ));
    InMux I__7220 (
            .O(N__32717),
            .I(N__32714));
    LocalMux I__7219 (
            .O(N__32714),
            .I(\b2v_inst6.count_1_i_a3_2_0 ));
    InMux I__7218 (
            .O(N__32711),
            .I(N__32705));
    InMux I__7217 (
            .O(N__32710),
            .I(N__32705));
    LocalMux I__7216 (
            .O(N__32705),
            .I(\b2v_inst6.N_389 ));
    CascadeMux I__7215 (
            .O(N__32702),
            .I(\b2v_inst6.N_389_cascade_ ));
    InMux I__7214 (
            .O(N__32699),
            .I(N__32696));
    LocalMux I__7213 (
            .O(N__32696),
            .I(\b2v_inst6.count_0_0 ));
    InMux I__7212 (
            .O(N__32693),
            .I(N__32690));
    LocalMux I__7211 (
            .O(N__32690),
            .I(\b2v_inst6.count_rst_13 ));
    CascadeMux I__7210 (
            .O(N__32687),
            .I(N__32684));
    InMux I__7209 (
            .O(N__32684),
            .I(N__32681));
    LocalMux I__7208 (
            .O(N__32681),
            .I(N__32677));
    InMux I__7207 (
            .O(N__32680),
            .I(N__32674));
    Span4Mux_s0_v I__7206 (
            .O(N__32677),
            .I(N__32671));
    LocalMux I__7205 (
            .O(N__32674),
            .I(\b2v_inst6.un2_count_1_axb_1 ));
    Odrv4 I__7204 (
            .O(N__32671),
            .I(\b2v_inst6.un2_count_1_axb_1 ));
    CascadeMux I__7203 (
            .O(N__32666),
            .I(\b2v_inst6.un2_count_1_axb_1_cascade_ ));
    InMux I__7202 (
            .O(N__32663),
            .I(N__32659));
    InMux I__7201 (
            .O(N__32662),
            .I(N__32656));
    LocalMux I__7200 (
            .O(N__32659),
            .I(\b2v_inst6.count_0_1 ));
    LocalMux I__7199 (
            .O(N__32656),
            .I(\b2v_inst6.count_0_1 ));
    SRMux I__7198 (
            .O(N__32651),
            .I(N__32645));
    SRMux I__7197 (
            .O(N__32650),
            .I(N__32642));
    InMux I__7196 (
            .O(N__32649),
            .I(N__32636));
    SRMux I__7195 (
            .O(N__32648),
            .I(N__32636));
    LocalMux I__7194 (
            .O(N__32645),
            .I(N__32630));
    LocalMux I__7193 (
            .O(N__32642),
            .I(N__32630));
    SRMux I__7192 (
            .O(N__32641),
            .I(N__32627));
    LocalMux I__7191 (
            .O(N__32636),
            .I(N__32604));
    SRMux I__7190 (
            .O(N__32635),
            .I(N__32601));
    Span4Mux_s2_v I__7189 (
            .O(N__32630),
            .I(N__32596));
    LocalMux I__7188 (
            .O(N__32627),
            .I(N__32596));
    InMux I__7187 (
            .O(N__32626),
            .I(N__32585));
    InMux I__7186 (
            .O(N__32625),
            .I(N__32585));
    InMux I__7185 (
            .O(N__32624),
            .I(N__32585));
    InMux I__7184 (
            .O(N__32623),
            .I(N__32585));
    InMux I__7183 (
            .O(N__32622),
            .I(N__32585));
    InMux I__7182 (
            .O(N__32621),
            .I(N__32577));
    InMux I__7181 (
            .O(N__32620),
            .I(N__32577));
    InMux I__7180 (
            .O(N__32619),
            .I(N__32570));
    InMux I__7179 (
            .O(N__32618),
            .I(N__32570));
    InMux I__7178 (
            .O(N__32617),
            .I(N__32570));
    InMux I__7177 (
            .O(N__32616),
            .I(N__32567));
    InMux I__7176 (
            .O(N__32615),
            .I(N__32562));
    InMux I__7175 (
            .O(N__32614),
            .I(N__32562));
    SRMux I__7174 (
            .O(N__32613),
            .I(N__32549));
    InMux I__7173 (
            .O(N__32612),
            .I(N__32549));
    InMux I__7172 (
            .O(N__32611),
            .I(N__32549));
    InMux I__7171 (
            .O(N__32610),
            .I(N__32549));
    InMux I__7170 (
            .O(N__32609),
            .I(N__32549));
    InMux I__7169 (
            .O(N__32608),
            .I(N__32549));
    SRMux I__7168 (
            .O(N__32607),
            .I(N__32544));
    Span4Mux_v I__7167 (
            .O(N__32604),
            .I(N__32536));
    LocalMux I__7166 (
            .O(N__32601),
            .I(N__32536));
    Span4Mux_v I__7165 (
            .O(N__32596),
            .I(N__32531));
    LocalMux I__7164 (
            .O(N__32585),
            .I(N__32531));
    InMux I__7163 (
            .O(N__32584),
            .I(N__32524));
    InMux I__7162 (
            .O(N__32583),
            .I(N__32524));
    InMux I__7161 (
            .O(N__32582),
            .I(N__32524));
    LocalMux I__7160 (
            .O(N__32577),
            .I(N__32517));
    LocalMux I__7159 (
            .O(N__32570),
            .I(N__32517));
    LocalMux I__7158 (
            .O(N__32567),
            .I(N__32517));
    LocalMux I__7157 (
            .O(N__32562),
            .I(N__32512));
    LocalMux I__7156 (
            .O(N__32549),
            .I(N__32512));
    InMux I__7155 (
            .O(N__32548),
            .I(N__32507));
    InMux I__7154 (
            .O(N__32547),
            .I(N__32507));
    LocalMux I__7153 (
            .O(N__32544),
            .I(N__32504));
    InMux I__7152 (
            .O(N__32543),
            .I(N__32497));
    InMux I__7151 (
            .O(N__32542),
            .I(N__32497));
    InMux I__7150 (
            .O(N__32541),
            .I(N__32497));
    Span4Mux_s2_v I__7149 (
            .O(N__32536),
            .I(N__32490));
    Span4Mux_s2_v I__7148 (
            .O(N__32531),
            .I(N__32490));
    LocalMux I__7147 (
            .O(N__32524),
            .I(N__32490));
    Span4Mux_s2_v I__7146 (
            .O(N__32517),
            .I(N__32483));
    Span4Mux_s1_h I__7145 (
            .O(N__32512),
            .I(N__32483));
    LocalMux I__7144 (
            .O(N__32507),
            .I(N__32483));
    Odrv12 I__7143 (
            .O(N__32504),
            .I(\b2v_inst6.curr_state_RNIM6FE1Z0Z_1 ));
    LocalMux I__7142 (
            .O(N__32497),
            .I(\b2v_inst6.curr_state_RNIM6FE1Z0Z_1 ));
    Odrv4 I__7141 (
            .O(N__32490),
            .I(\b2v_inst6.curr_state_RNIM6FE1Z0Z_1 ));
    Odrv4 I__7140 (
            .O(N__32483),
            .I(\b2v_inst6.curr_state_RNIM6FE1Z0Z_1 ));
    InMux I__7139 (
            .O(N__32474),
            .I(N__32471));
    LocalMux I__7138 (
            .O(N__32471),
            .I(\b2v_inst6.count_rst_5 ));
    InMux I__7137 (
            .O(N__32468),
            .I(N__32464));
    InMux I__7136 (
            .O(N__32467),
            .I(N__32461));
    LocalMux I__7135 (
            .O(N__32464),
            .I(\b2v_inst6.count_0_9 ));
    LocalMux I__7134 (
            .O(N__32461),
            .I(\b2v_inst6.count_0_9 ));
    CascadeMux I__7133 (
            .O(N__32456),
            .I(N__32452));
    InMux I__7132 (
            .O(N__32455),
            .I(N__32448));
    InMux I__7131 (
            .O(N__32452),
            .I(N__32445));
    InMux I__7130 (
            .O(N__32451),
            .I(N__32442));
    LocalMux I__7129 (
            .O(N__32448),
            .I(N__32439));
    LocalMux I__7128 (
            .O(N__32445),
            .I(\b2v_inst6.countZ0Z_8 ));
    LocalMux I__7127 (
            .O(N__32442),
            .I(\b2v_inst6.countZ0Z_8 ));
    Odrv12 I__7126 (
            .O(N__32439),
            .I(\b2v_inst6.countZ0Z_8 ));
    CEMux I__7125 (
            .O(N__32432),
            .I(N__32424));
    CascadeMux I__7124 (
            .O(N__32431),
            .I(N__32419));
    CEMux I__7123 (
            .O(N__32430),
            .I(N__32416));
    CEMux I__7122 (
            .O(N__32429),
            .I(N__32413));
    CEMux I__7121 (
            .O(N__32428),
            .I(N__32410));
    CEMux I__7120 (
            .O(N__32427),
            .I(N__32407));
    LocalMux I__7119 (
            .O(N__32424),
            .I(N__32404));
    CEMux I__7118 (
            .O(N__32423),
            .I(N__32401));
    CEMux I__7117 (
            .O(N__32422),
            .I(N__32398));
    InMux I__7116 (
            .O(N__32419),
            .I(N__32393));
    LocalMux I__7115 (
            .O(N__32416),
            .I(N__32390));
    LocalMux I__7114 (
            .O(N__32413),
            .I(N__32383));
    LocalMux I__7113 (
            .O(N__32410),
            .I(N__32383));
    LocalMux I__7112 (
            .O(N__32407),
            .I(N__32383));
    Span4Mux_s0_v I__7111 (
            .O(N__32404),
            .I(N__32378));
    LocalMux I__7110 (
            .O(N__32401),
            .I(N__32378));
    LocalMux I__7109 (
            .O(N__32398),
            .I(N__32369));
    InMux I__7108 (
            .O(N__32397),
            .I(N__32353));
    InMux I__7107 (
            .O(N__32396),
            .I(N__32353));
    LocalMux I__7106 (
            .O(N__32393),
            .I(N__32344));
    IoSpan4Mux I__7105 (
            .O(N__32390),
            .I(N__32344));
    Span4Mux_v I__7104 (
            .O(N__32383),
            .I(N__32344));
    Span4Mux_v I__7103 (
            .O(N__32378),
            .I(N__32344));
    InMux I__7102 (
            .O(N__32377),
            .I(N__32333));
    InMux I__7101 (
            .O(N__32376),
            .I(N__32333));
    InMux I__7100 (
            .O(N__32375),
            .I(N__32333));
    InMux I__7099 (
            .O(N__32374),
            .I(N__32333));
    InMux I__7098 (
            .O(N__32373),
            .I(N__32333));
    InMux I__7097 (
            .O(N__32372),
            .I(N__32327));
    Span4Mux_s1_v I__7096 (
            .O(N__32369),
            .I(N__32324));
    InMux I__7095 (
            .O(N__32368),
            .I(N__32317));
    InMux I__7094 (
            .O(N__32367),
            .I(N__32317));
    InMux I__7093 (
            .O(N__32366),
            .I(N__32317));
    InMux I__7092 (
            .O(N__32365),
            .I(N__32312));
    InMux I__7091 (
            .O(N__32364),
            .I(N__32312));
    InMux I__7090 (
            .O(N__32363),
            .I(N__32303));
    InMux I__7089 (
            .O(N__32362),
            .I(N__32303));
    InMux I__7088 (
            .O(N__32361),
            .I(N__32303));
    InMux I__7087 (
            .O(N__32360),
            .I(N__32303));
    InMux I__7086 (
            .O(N__32359),
            .I(N__32298));
    InMux I__7085 (
            .O(N__32358),
            .I(N__32298));
    LocalMux I__7084 (
            .O(N__32353),
            .I(N__32295));
    Span4Mux_s0_v I__7083 (
            .O(N__32344),
            .I(N__32290));
    LocalMux I__7082 (
            .O(N__32333),
            .I(N__32290));
    InMux I__7081 (
            .O(N__32332),
            .I(N__32283));
    InMux I__7080 (
            .O(N__32331),
            .I(N__32283));
    InMux I__7079 (
            .O(N__32330),
            .I(N__32283));
    LocalMux I__7078 (
            .O(N__32327),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7077 (
            .O(N__32324),
            .I(\b2v_inst6.count_en ));
    LocalMux I__7076 (
            .O(N__32317),
            .I(\b2v_inst6.count_en ));
    LocalMux I__7075 (
            .O(N__32312),
            .I(\b2v_inst6.count_en ));
    LocalMux I__7074 (
            .O(N__32303),
            .I(\b2v_inst6.count_en ));
    LocalMux I__7073 (
            .O(N__32298),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7072 (
            .O(N__32295),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7071 (
            .O(N__32290),
            .I(\b2v_inst6.count_en ));
    LocalMux I__7070 (
            .O(N__32283),
            .I(\b2v_inst6.count_en ));
    InMux I__7069 (
            .O(N__32264),
            .I(N__32261));
    LocalMux I__7068 (
            .O(N__32261),
            .I(N__32258));
    Odrv4 I__7067 (
            .O(N__32258),
            .I(\b2v_inst6.count_1_i_a3_4_0 ));
    InMux I__7066 (
            .O(N__32255),
            .I(N__32252));
    LocalMux I__7065 (
            .O(N__32252),
            .I(N__32249));
    Span4Mux_v I__7064 (
            .O(N__32249),
            .I(N__32245));
    InMux I__7063 (
            .O(N__32248),
            .I(N__32242));
    Odrv4 I__7062 (
            .O(N__32245),
            .I(\b2v_inst5.N_51 ));
    LocalMux I__7061 (
            .O(N__32242),
            .I(\b2v_inst5.N_51 ));
    CascadeMux I__7060 (
            .O(N__32237),
            .I(N__32234));
    InMux I__7059 (
            .O(N__32234),
            .I(N__32231));
    LocalMux I__7058 (
            .O(N__32231),
            .I(N__32228));
    Odrv12 I__7057 (
            .O(N__32228),
            .I(\b2v_inst5.curr_state_0_1 ));
    CascadeMux I__7056 (
            .O(N__32225),
            .I(N__32216));
    CascadeMux I__7055 (
            .O(N__32224),
            .I(N__32211));
    InMux I__7054 (
            .O(N__32223),
            .I(N__32208));
    InMux I__7053 (
            .O(N__32222),
            .I(N__32205));
    InMux I__7052 (
            .O(N__32221),
            .I(N__32202));
    InMux I__7051 (
            .O(N__32220),
            .I(N__32199));
    InMux I__7050 (
            .O(N__32219),
            .I(N__32196));
    InMux I__7049 (
            .O(N__32216),
            .I(N__32191));
    InMux I__7048 (
            .O(N__32215),
            .I(N__32191));
    InMux I__7047 (
            .O(N__32214),
            .I(N__32188));
    InMux I__7046 (
            .O(N__32211),
            .I(N__32185));
    LocalMux I__7045 (
            .O(N__32208),
            .I(N__32170));
    LocalMux I__7044 (
            .O(N__32205),
            .I(N__32167));
    LocalMux I__7043 (
            .O(N__32202),
            .I(N__32164));
    LocalMux I__7042 (
            .O(N__32199),
            .I(N__32161));
    LocalMux I__7041 (
            .O(N__32196),
            .I(N__32158));
    LocalMux I__7040 (
            .O(N__32191),
            .I(N__32155));
    LocalMux I__7039 (
            .O(N__32188),
            .I(N__32152));
    LocalMux I__7038 (
            .O(N__32185),
            .I(N__32149));
    CEMux I__7037 (
            .O(N__32184),
            .I(N__32108));
    CEMux I__7036 (
            .O(N__32183),
            .I(N__32108));
    CEMux I__7035 (
            .O(N__32182),
            .I(N__32108));
    CEMux I__7034 (
            .O(N__32181),
            .I(N__32108));
    CEMux I__7033 (
            .O(N__32180),
            .I(N__32108));
    CEMux I__7032 (
            .O(N__32179),
            .I(N__32108));
    CEMux I__7031 (
            .O(N__32178),
            .I(N__32108));
    CEMux I__7030 (
            .O(N__32177),
            .I(N__32108));
    CEMux I__7029 (
            .O(N__32176),
            .I(N__32108));
    CEMux I__7028 (
            .O(N__32175),
            .I(N__32108));
    CEMux I__7027 (
            .O(N__32174),
            .I(N__32108));
    CEMux I__7026 (
            .O(N__32173),
            .I(N__32108));
    Glb2LocalMux I__7025 (
            .O(N__32170),
            .I(N__32108));
    Glb2LocalMux I__7024 (
            .O(N__32167),
            .I(N__32108));
    Glb2LocalMux I__7023 (
            .O(N__32164),
            .I(N__32108));
    Glb2LocalMux I__7022 (
            .O(N__32161),
            .I(N__32108));
    Glb2LocalMux I__7021 (
            .O(N__32158),
            .I(N__32108));
    Glb2LocalMux I__7020 (
            .O(N__32155),
            .I(N__32108));
    Glb2LocalMux I__7019 (
            .O(N__32152),
            .I(N__32108));
    Glb2LocalMux I__7018 (
            .O(N__32149),
            .I(N__32108));
    GlobalMux I__7017 (
            .O(N__32108),
            .I(N__32105));
    gio2CtrlBuf I__7016 (
            .O(N__32105),
            .I(N_606_g));
    InMux I__7015 (
            .O(N__32102),
            .I(N__32097));
    InMux I__7014 (
            .O(N__32101),
            .I(N__32094));
    InMux I__7013 (
            .O(N__32100),
            .I(N__32091));
    LocalMux I__7012 (
            .O(N__32097),
            .I(N__32088));
    LocalMux I__7011 (
            .O(N__32094),
            .I(N__32085));
    LocalMux I__7010 (
            .O(N__32091),
            .I(\b2v_inst6.countZ0Z_0 ));
    Odrv4 I__7009 (
            .O(N__32088),
            .I(\b2v_inst6.countZ0Z_0 ));
    Odrv4 I__7008 (
            .O(N__32085),
            .I(\b2v_inst6.countZ0Z_0 ));
    InMux I__7007 (
            .O(N__32078),
            .I(N__32073));
    InMux I__7006 (
            .O(N__32077),
            .I(N__32068));
    InMux I__7005 (
            .O(N__32076),
            .I(N__32068));
    LocalMux I__7004 (
            .O(N__32073),
            .I(N__32063));
    LocalMux I__7003 (
            .O(N__32068),
            .I(N__32063));
    Odrv4 I__7002 (
            .O(N__32063),
            .I(\b2v_inst6.N_3036_i ));
    IoInMux I__7001 (
            .O(N__32060),
            .I(N__32056));
    CascadeMux I__7000 (
            .O(N__32059),
            .I(N__32053));
    LocalMux I__6999 (
            .O(N__32056),
            .I(N__32049));
    InMux I__6998 (
            .O(N__32053),
            .I(N__32043));
    InMux I__6997 (
            .O(N__32052),
            .I(N__32043));
    Span4Mux_s3_h I__6996 (
            .O(N__32049),
            .I(N__32040));
    InMux I__6995 (
            .O(N__32048),
            .I(N__32037));
    LocalMux I__6994 (
            .O(N__32043),
            .I(N__32034));
    Span4Mux_v I__6993 (
            .O(N__32040),
            .I(N__32029));
    LocalMux I__6992 (
            .O(N__32037),
            .I(N__32029));
    Span4Mux_h I__6991 (
            .O(N__32034),
            .I(N__32024));
    Span4Mux_h I__6990 (
            .O(N__32029),
            .I(N__32024));
    Span4Mux_h I__6989 (
            .O(N__32024),
            .I(N__32021));
    Odrv4 I__6988 (
            .O(N__32021),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__6987 (
            .O(N__32018),
            .I(\b2v_inst6.count_rst_9_cascade_ ));
    InMux I__6986 (
            .O(N__32015),
            .I(N__32010));
    InMux I__6985 (
            .O(N__32014),
            .I(N__32007));
    InMux I__6984 (
            .O(N__32013),
            .I(N__32004));
    LocalMux I__6983 (
            .O(N__32010),
            .I(N__32001));
    LocalMux I__6982 (
            .O(N__32007),
            .I(\b2v_inst6.countZ0Z_5 ));
    LocalMux I__6981 (
            .O(N__32004),
            .I(\b2v_inst6.countZ0Z_5 ));
    Odrv4 I__6980 (
            .O(N__32001),
            .I(\b2v_inst6.countZ0Z_5 ));
    InMux I__6979 (
            .O(N__31994),
            .I(N__31988));
    InMux I__6978 (
            .O(N__31993),
            .I(N__31988));
    LocalMux I__6977 (
            .O(N__31988),
            .I(N__31985));
    Odrv4 I__6976 (
            .O(N__31985),
            .I(\b2v_inst6.un2_count_1_cry_4_THRU_CO ));
    CascadeMux I__6975 (
            .O(N__31982),
            .I(\b2v_inst6.countZ0Z_5_cascade_ ));
    InMux I__6974 (
            .O(N__31979),
            .I(N__31976));
    LocalMux I__6973 (
            .O(N__31976),
            .I(\b2v_inst6.count_0_5 ));
    CascadeMux I__6972 (
            .O(N__31973),
            .I(N__31970));
    InMux I__6971 (
            .O(N__31970),
            .I(N__31967));
    LocalMux I__6970 (
            .O(N__31967),
            .I(N__31963));
    InMux I__6969 (
            .O(N__31966),
            .I(N__31960));
    Odrv4 I__6968 (
            .O(N__31963),
            .I(\b2v_inst6.un2_count_1_cry_10_THRU_CO ));
    LocalMux I__6967 (
            .O(N__31960),
            .I(\b2v_inst6.un2_count_1_cry_10_THRU_CO ));
    InMux I__6966 (
            .O(N__31955),
            .I(N__31936));
    InMux I__6965 (
            .O(N__31954),
            .I(N__31936));
    InMux I__6964 (
            .O(N__31953),
            .I(N__31931));
    InMux I__6963 (
            .O(N__31952),
            .I(N__31931));
    InMux I__6962 (
            .O(N__31951),
            .I(N__31924));
    InMux I__6961 (
            .O(N__31950),
            .I(N__31924));
    InMux I__6960 (
            .O(N__31949),
            .I(N__31924));
    InMux I__6959 (
            .O(N__31948),
            .I(N__31912));
    InMux I__6958 (
            .O(N__31947),
            .I(N__31912));
    InMux I__6957 (
            .O(N__31946),
            .I(N__31912));
    InMux I__6956 (
            .O(N__31945),
            .I(N__31912));
    InMux I__6955 (
            .O(N__31944),
            .I(N__31912));
    InMux I__6954 (
            .O(N__31943),
            .I(N__31909));
    InMux I__6953 (
            .O(N__31942),
            .I(N__31904));
    InMux I__6952 (
            .O(N__31941),
            .I(N__31904));
    LocalMux I__6951 (
            .O(N__31936),
            .I(N__31897));
    LocalMux I__6950 (
            .O(N__31931),
            .I(N__31897));
    LocalMux I__6949 (
            .O(N__31924),
            .I(N__31897));
    InMux I__6948 (
            .O(N__31923),
            .I(N__31894));
    LocalMux I__6947 (
            .O(N__31912),
            .I(N__31891));
    LocalMux I__6946 (
            .O(N__31909),
            .I(N__31884));
    LocalMux I__6945 (
            .O(N__31904),
            .I(N__31884));
    Span4Mux_v I__6944 (
            .O(N__31897),
            .I(N__31884));
    LocalMux I__6943 (
            .O(N__31894),
            .I(\b2v_inst6.N_394 ));
    Odrv4 I__6942 (
            .O(N__31891),
            .I(\b2v_inst6.N_394 ));
    Odrv4 I__6941 (
            .O(N__31884),
            .I(\b2v_inst6.N_394 ));
    CascadeMux I__6940 (
            .O(N__31877),
            .I(\b2v_inst6.count_rst_3_cascade_ ));
    InMux I__6939 (
            .O(N__31874),
            .I(N__31871));
    LocalMux I__6938 (
            .O(N__31871),
            .I(N__31868));
    Odrv4 I__6937 (
            .O(N__31868),
            .I(\b2v_inst6.count_0_11 ));
    InMux I__6936 (
            .O(N__31865),
            .I(N__31862));
    LocalMux I__6935 (
            .O(N__31862),
            .I(\b2v_inst6.count_RNIM6FE1Z0Z_0 ));
    CascadeMux I__6934 (
            .O(N__31859),
            .I(\b2v_inst6.countZ0Z_0_cascade_ ));
    CascadeMux I__6933 (
            .O(N__31856),
            .I(N__31851));
    InMux I__6932 (
            .O(N__31855),
            .I(N__31848));
    InMux I__6931 (
            .O(N__31854),
            .I(N__31844));
    InMux I__6930 (
            .O(N__31851),
            .I(N__31841));
    LocalMux I__6929 (
            .O(N__31848),
            .I(N__31838));
    InMux I__6928 (
            .O(N__31847),
            .I(N__31835));
    LocalMux I__6927 (
            .O(N__31844),
            .I(\b2v_inst6.countZ0Z_11 ));
    LocalMux I__6926 (
            .O(N__31841),
            .I(\b2v_inst6.countZ0Z_11 ));
    Odrv12 I__6925 (
            .O(N__31838),
            .I(\b2v_inst6.countZ0Z_11 ));
    LocalMux I__6924 (
            .O(N__31835),
            .I(\b2v_inst6.countZ0Z_11 ));
    CascadeMux I__6923 (
            .O(N__31826),
            .I(\b2v_inst6.count_rst_13_cascade_ ));
    InMux I__6922 (
            .O(N__31823),
            .I(N__31820));
    LocalMux I__6921 (
            .O(N__31820),
            .I(N__31817));
    Odrv4 I__6920 (
            .O(N__31817),
            .I(\b2v_inst6.count_1_i_a3_5_0 ));
    InMux I__6919 (
            .O(N__31814),
            .I(N__31811));
    LocalMux I__6918 (
            .O(N__31811),
            .I(N__31808));
    Odrv12 I__6917 (
            .O(N__31808),
            .I(\b2v_inst6.count_1_i_a3_6_0 ));
    CascadeMux I__6916 (
            .O(N__31805),
            .I(\b2v_inst6.count_1_i_a3_3_0_cascade_ ));
    InMux I__6915 (
            .O(N__31802),
            .I(N__31799));
    LocalMux I__6914 (
            .O(N__31799),
            .I(\b2v_inst6.count_0_14 ));
    InMux I__6913 (
            .O(N__31796),
            .I(N__31790));
    InMux I__6912 (
            .O(N__31795),
            .I(N__31790));
    LocalMux I__6911 (
            .O(N__31790),
            .I(\b2v_inst6.un2_count_1_cry_13_c_RNI06SPZ0Z1 ));
    InMux I__6910 (
            .O(N__31787),
            .I(N__31784));
    LocalMux I__6909 (
            .O(N__31784),
            .I(\b2v_inst6.countZ0Z_14 ));
    InMux I__6908 (
            .O(N__31781),
            .I(N__31777));
    InMux I__6907 (
            .O(N__31780),
            .I(N__31774));
    LocalMux I__6906 (
            .O(N__31777),
            .I(\b2v_inst6.count_0_2 ));
    LocalMux I__6905 (
            .O(N__31774),
            .I(\b2v_inst6.count_0_2 ));
    CascadeMux I__6904 (
            .O(N__31769),
            .I(\b2v_inst6.countZ0Z_14_cascade_ ));
    InMux I__6903 (
            .O(N__31766),
            .I(N__31757));
    InMux I__6902 (
            .O(N__31765),
            .I(N__31757));
    InMux I__6901 (
            .O(N__31764),
            .I(N__31757));
    LocalMux I__6900 (
            .O(N__31757),
            .I(\b2v_inst6.count_rst_12 ));
    InMux I__6899 (
            .O(N__31754),
            .I(N__31751));
    LocalMux I__6898 (
            .O(N__31751),
            .I(\b2v_inst6.un2_count_1_axb_12 ));
    InMux I__6897 (
            .O(N__31748),
            .I(N__31745));
    LocalMux I__6896 (
            .O(N__31745),
            .I(N__31740));
    InMux I__6895 (
            .O(N__31744),
            .I(N__31735));
    InMux I__6894 (
            .O(N__31743),
            .I(N__31735));
    Odrv4 I__6893 (
            .O(N__31740),
            .I(\b2v_inst6.count_rst_2 ));
    LocalMux I__6892 (
            .O(N__31735),
            .I(\b2v_inst6.count_rst_2 ));
    InMux I__6891 (
            .O(N__31730),
            .I(N__31727));
    LocalMux I__6890 (
            .O(N__31727),
            .I(N__31724));
    Span4Mux_v I__6889 (
            .O(N__31724),
            .I(N__31720));
    InMux I__6888 (
            .O(N__31723),
            .I(N__31717));
    Odrv4 I__6887 (
            .O(N__31720),
            .I(\b2v_inst6.count_0_12 ));
    LocalMux I__6886 (
            .O(N__31717),
            .I(\b2v_inst6.count_0_12 ));
    InMux I__6885 (
            .O(N__31712),
            .I(N__31705));
    InMux I__6884 (
            .O(N__31711),
            .I(N__31705));
    InMux I__6883 (
            .O(N__31710),
            .I(N__31702));
    LocalMux I__6882 (
            .O(N__31705),
            .I(\b2v_inst6.count_rst_1 ));
    LocalMux I__6881 (
            .O(N__31702),
            .I(\b2v_inst6.count_rst_1 ));
    InMux I__6880 (
            .O(N__31697),
            .I(N__31693));
    InMux I__6879 (
            .O(N__31696),
            .I(N__31690));
    LocalMux I__6878 (
            .O(N__31693),
            .I(N__31687));
    LocalMux I__6877 (
            .O(N__31690),
            .I(\b2v_inst6.count_0_13 ));
    Odrv4 I__6876 (
            .O(N__31687),
            .I(\b2v_inst6.count_0_13 ));
    InMux I__6875 (
            .O(N__31682),
            .I(N__31679));
    LocalMux I__6874 (
            .O(N__31679),
            .I(\b2v_inst6.un2_count_1_axb_13 ));
    InMux I__6873 (
            .O(N__31676),
            .I(N__31673));
    LocalMux I__6872 (
            .O(N__31673),
            .I(N__31669));
    InMux I__6871 (
            .O(N__31672),
            .I(N__31666));
    Span4Mux_s1_h I__6870 (
            .O(N__31669),
            .I(N__31663));
    LocalMux I__6869 (
            .O(N__31666),
            .I(N__31660));
    Odrv4 I__6868 (
            .O(N__31663),
            .I(\b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ));
    Odrv4 I__6867 (
            .O(N__31660),
            .I(\b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ));
    InMux I__6866 (
            .O(N__31655),
            .I(N__31652));
    LocalMux I__6865 (
            .O(N__31652),
            .I(\b2v_inst6.count_0_6 ));
    CascadeMux I__6864 (
            .O(N__31649),
            .I(\b2v_inst6.N_394_cascade_ ));
    InMux I__6863 (
            .O(N__31646),
            .I(N__31640));
    InMux I__6862 (
            .O(N__31645),
            .I(N__31640));
    LocalMux I__6861 (
            .O(N__31640),
            .I(\b2v_inst6.un2_count_1_cry_3_THRU_CO ));
    CascadeMux I__6860 (
            .O(N__31637),
            .I(\b2v_inst6.un2_count_1_axb_4_cascade_ ));
    InMux I__6859 (
            .O(N__31634),
            .I(N__31631));
    LocalMux I__6858 (
            .O(N__31631),
            .I(\b2v_inst6.count_rst_10 ));
    InMux I__6857 (
            .O(N__31628),
            .I(N__31622));
    InMux I__6856 (
            .O(N__31627),
            .I(N__31622));
    LocalMux I__6855 (
            .O(N__31622),
            .I(\b2v_inst6.count_0_4 ));
    CascadeMux I__6854 (
            .O(N__31619),
            .I(\b2v_inst6.count_rst_11_cascade_ ));
    CascadeMux I__6853 (
            .O(N__31616),
            .I(N__31612));
    CascadeMux I__6852 (
            .O(N__31615),
            .I(N__31608));
    InMux I__6851 (
            .O(N__31612),
            .I(N__31605));
    InMux I__6850 (
            .O(N__31611),
            .I(N__31602));
    InMux I__6849 (
            .O(N__31608),
            .I(N__31599));
    LocalMux I__6848 (
            .O(N__31605),
            .I(\b2v_inst6.countZ0Z_3 ));
    LocalMux I__6847 (
            .O(N__31602),
            .I(\b2v_inst6.countZ0Z_3 ));
    LocalMux I__6846 (
            .O(N__31599),
            .I(\b2v_inst6.countZ0Z_3 ));
    InMux I__6845 (
            .O(N__31592),
            .I(N__31586));
    InMux I__6844 (
            .O(N__31591),
            .I(N__31586));
    LocalMux I__6843 (
            .O(N__31586),
            .I(\b2v_inst6.un2_count_1_cry_2_THRU_CO ));
    CascadeMux I__6842 (
            .O(N__31583),
            .I(\b2v_inst6.countZ0Z_3_cascade_ ));
    InMux I__6841 (
            .O(N__31580),
            .I(N__31577));
    LocalMux I__6840 (
            .O(N__31577),
            .I(\b2v_inst6.count_0_3 ));
    InMux I__6839 (
            .O(N__31574),
            .I(N__31571));
    LocalMux I__6838 (
            .O(N__31571),
            .I(\b2v_inst6.un2_count_1_axb_2 ));
    InMux I__6837 (
            .O(N__31568),
            .I(N__31562));
    InMux I__6836 (
            .O(N__31567),
            .I(N__31562));
    LocalMux I__6835 (
            .O(N__31562),
            .I(\b2v_inst11.un3_count_off_1_cry_14_c_RNI7DTZ0Z63 ));
    InMux I__6834 (
            .O(N__31559),
            .I(N__31556));
    LocalMux I__6833 (
            .O(N__31556),
            .I(\b2v_inst11.count_off_0_15 ));
    InMux I__6832 (
            .O(N__31553),
            .I(N__31547));
    InMux I__6831 (
            .O(N__31552),
            .I(N__31547));
    LocalMux I__6830 (
            .O(N__31547),
            .I(N__31544));
    Odrv4 I__6829 (
            .O(N__31544),
            .I(\b2v_inst11.count_off_1_6 ));
    InMux I__6828 (
            .O(N__31541),
            .I(N__31538));
    LocalMux I__6827 (
            .O(N__31538),
            .I(\b2v_inst11.count_off_0_6 ));
    InMux I__6826 (
            .O(N__31535),
            .I(N__31529));
    InMux I__6825 (
            .O(N__31534),
            .I(N__31529));
    LocalMux I__6824 (
            .O(N__31529),
            .I(N__31526));
    Odrv4 I__6823 (
            .O(N__31526),
            .I(\b2v_inst11.count_off_1_7 ));
    InMux I__6822 (
            .O(N__31523),
            .I(N__31520));
    LocalMux I__6821 (
            .O(N__31520),
            .I(\b2v_inst11.count_off_0_7 ));
    InMux I__6820 (
            .O(N__31517),
            .I(N__31511));
    InMux I__6819 (
            .O(N__31516),
            .I(N__31511));
    LocalMux I__6818 (
            .O(N__31511),
            .I(N__31508));
    Odrv4 I__6817 (
            .O(N__31508),
            .I(\b2v_inst11.count_off_1_8 ));
    InMux I__6816 (
            .O(N__31505),
            .I(N__31502));
    LocalMux I__6815 (
            .O(N__31502),
            .I(\b2v_inst11.count_off_0_8 ));
    CascadeMux I__6814 (
            .O(N__31499),
            .I(\b2v_inst6.count_rst_10_cascade_ ));
    CascadeMux I__6813 (
            .O(N__31496),
            .I(N__31492));
    CascadeMux I__6812 (
            .O(N__31495),
            .I(N__31489));
    InMux I__6811 (
            .O(N__31492),
            .I(N__31486));
    InMux I__6810 (
            .O(N__31489),
            .I(N__31483));
    LocalMux I__6809 (
            .O(N__31486),
            .I(\b2v_inst6.un2_count_1_axb_4 ));
    LocalMux I__6808 (
            .O(N__31483),
            .I(\b2v_inst6.un2_count_1_axb_4 ));
    InMux I__6807 (
            .O(N__31478),
            .I(\b2v_inst11.un3_count_off_1_cry_7 ));
    InMux I__6806 (
            .O(N__31475),
            .I(bfn_11_14_0_));
    InMux I__6805 (
            .O(N__31472),
            .I(\b2v_inst11.un3_count_off_1_cry_9 ));
    InMux I__6804 (
            .O(N__31469),
            .I(\b2v_inst11.un3_count_off_1_cry_10 ));
    InMux I__6803 (
            .O(N__31466),
            .I(\b2v_inst11.un3_count_off_1_cry_11 ));
    InMux I__6802 (
            .O(N__31463),
            .I(\b2v_inst11.un3_count_off_1_cry_12 ));
    InMux I__6801 (
            .O(N__31460),
            .I(\b2v_inst11.un3_count_off_1_cry_13 ));
    InMux I__6800 (
            .O(N__31457),
            .I(\b2v_inst11.un3_count_off_1_cry_14 ));
    InMux I__6799 (
            .O(N__31454),
            .I(N__31450));
    InMux I__6798 (
            .O(N__31453),
            .I(N__31447));
    LocalMux I__6797 (
            .O(N__31450),
            .I(N__31444));
    LocalMux I__6796 (
            .O(N__31447),
            .I(\b2v_inst11.count_off_1_14 ));
    Odrv4 I__6795 (
            .O(N__31444),
            .I(\b2v_inst11.count_off_1_14 ));
    InMux I__6794 (
            .O(N__31439),
            .I(N__31436));
    LocalMux I__6793 (
            .O(N__31436),
            .I(N__31433));
    Odrv4 I__6792 (
            .O(N__31433),
            .I(\b2v_inst11.count_off_0_14 ));
    CascadeMux I__6791 (
            .O(N__31430),
            .I(\b2v_inst11.N_125_cascade_ ));
    InMux I__6790 (
            .O(N__31427),
            .I(N__31424));
    LocalMux I__6789 (
            .O(N__31424),
            .I(N__31421));
    Span4Mux_v I__6788 (
            .O(N__31421),
            .I(N__31417));
    InMux I__6787 (
            .O(N__31420),
            .I(N__31414));
    Odrv4 I__6786 (
            .O(N__31417),
            .I(\b2v_inst11.N_382_N ));
    LocalMux I__6785 (
            .O(N__31414),
            .I(\b2v_inst11.N_382_N ));
    InMux I__6784 (
            .O(N__31409),
            .I(\b2v_inst11.un3_count_off_1_cry_1 ));
    InMux I__6783 (
            .O(N__31406),
            .I(\b2v_inst11.un3_count_off_1_cry_2 ));
    InMux I__6782 (
            .O(N__31403),
            .I(\b2v_inst11.un3_count_off_1_cry_3 ));
    InMux I__6781 (
            .O(N__31400),
            .I(\b2v_inst11.un3_count_off_1_cry_4 ));
    InMux I__6780 (
            .O(N__31397),
            .I(\b2v_inst11.un3_count_off_1_cry_5 ));
    InMux I__6779 (
            .O(N__31394),
            .I(\b2v_inst11.un3_count_off_1_cry_6 ));
    CascadeMux I__6778 (
            .O(N__31391),
            .I(N__31388));
    InMux I__6777 (
            .O(N__31388),
            .I(N__31382));
    InMux I__6776 (
            .O(N__31387),
            .I(N__31382));
    LocalMux I__6775 (
            .O(N__31382),
            .I(\b2v_inst11.N_119_f0_1 ));
    InMux I__6774 (
            .O(N__31379),
            .I(N__31370));
    CascadeMux I__6773 (
            .O(N__31378),
            .I(N__31366));
    CascadeMux I__6772 (
            .O(N__31377),
            .I(N__31361));
    InMux I__6771 (
            .O(N__31376),
            .I(N__31358));
    InMux I__6770 (
            .O(N__31375),
            .I(N__31351));
    InMux I__6769 (
            .O(N__31374),
            .I(N__31351));
    InMux I__6768 (
            .O(N__31373),
            .I(N__31351));
    LocalMux I__6767 (
            .O(N__31370),
            .I(N__31347));
    InMux I__6766 (
            .O(N__31369),
            .I(N__31344));
    InMux I__6765 (
            .O(N__31366),
            .I(N__31339));
    InMux I__6764 (
            .O(N__31365),
            .I(N__31339));
    CascadeMux I__6763 (
            .O(N__31364),
            .I(N__31336));
    InMux I__6762 (
            .O(N__31361),
            .I(N__31333));
    LocalMux I__6761 (
            .O(N__31358),
            .I(N__31327));
    LocalMux I__6760 (
            .O(N__31351),
            .I(N__31327));
    InMux I__6759 (
            .O(N__31350),
            .I(N__31324));
    Span4Mux_s1_v I__6758 (
            .O(N__31347),
            .I(N__31319));
    LocalMux I__6757 (
            .O(N__31344),
            .I(N__31319));
    LocalMux I__6756 (
            .O(N__31339),
            .I(N__31316));
    InMux I__6755 (
            .O(N__31336),
            .I(N__31313));
    LocalMux I__6754 (
            .O(N__31333),
            .I(N__31306));
    InMux I__6753 (
            .O(N__31332),
            .I(N__31303));
    Span4Mux_v I__6752 (
            .O(N__31327),
            .I(N__31298));
    LocalMux I__6751 (
            .O(N__31324),
            .I(N__31298));
    Span4Mux_v I__6750 (
            .O(N__31319),
            .I(N__31291));
    Span4Mux_v I__6749 (
            .O(N__31316),
            .I(N__31291));
    LocalMux I__6748 (
            .O(N__31313),
            .I(N__31291));
    InMux I__6747 (
            .O(N__31312),
            .I(N__31288));
    InMux I__6746 (
            .O(N__31311),
            .I(N__31283));
    InMux I__6745 (
            .O(N__31310),
            .I(N__31283));
    InMux I__6744 (
            .O(N__31309),
            .I(N__31280));
    Span4Mux_h I__6743 (
            .O(N__31306),
            .I(N__31277));
    LocalMux I__6742 (
            .O(N__31303),
            .I(N__31272));
    Span4Mux_h I__6741 (
            .O(N__31298),
            .I(N__31272));
    Span4Mux_h I__6740 (
            .O(N__31291),
            .I(N__31267));
    LocalMux I__6739 (
            .O(N__31288),
            .I(N__31267));
    LocalMux I__6738 (
            .O(N__31283),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__6737 (
            .O(N__31280),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__6736 (
            .O(N__31277),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__6735 (
            .O(N__31272),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__6734 (
            .O(N__31267),
            .I(\b2v_inst11.dutycycle ));
    InMux I__6733 (
            .O(N__31256),
            .I(N__31253));
    LocalMux I__6732 (
            .O(N__31253),
            .I(\b2v_inst11.dutycycle_eena_0 ));
    IoInMux I__6731 (
            .O(N__31250),
            .I(N__31245));
    InMux I__6730 (
            .O(N__31249),
            .I(N__31241));
    CascadeMux I__6729 (
            .O(N__31248),
            .I(N__31232));
    LocalMux I__6728 (
            .O(N__31245),
            .I(N__31229));
    CascadeMux I__6727 (
            .O(N__31244),
            .I(N__31222));
    LocalMux I__6726 (
            .O(N__31241),
            .I(N__31218));
    InMux I__6725 (
            .O(N__31240),
            .I(N__31215));
    InMux I__6724 (
            .O(N__31239),
            .I(N__31212));
    InMux I__6723 (
            .O(N__31238),
            .I(N__31200));
    InMux I__6722 (
            .O(N__31237),
            .I(N__31200));
    InMux I__6721 (
            .O(N__31236),
            .I(N__31200));
    InMux I__6720 (
            .O(N__31235),
            .I(N__31200));
    InMux I__6719 (
            .O(N__31232),
            .I(N__31197));
    IoSpan4Mux I__6718 (
            .O(N__31229),
            .I(N__31186));
    InMux I__6717 (
            .O(N__31228),
            .I(N__31177));
    InMux I__6716 (
            .O(N__31227),
            .I(N__31177));
    InMux I__6715 (
            .O(N__31226),
            .I(N__31177));
    InMux I__6714 (
            .O(N__31225),
            .I(N__31177));
    InMux I__6713 (
            .O(N__31222),
            .I(N__31172));
    InMux I__6712 (
            .O(N__31221),
            .I(N__31172));
    Span4Mux_h I__6711 (
            .O(N__31218),
            .I(N__31165));
    LocalMux I__6710 (
            .O(N__31215),
            .I(N__31165));
    LocalMux I__6709 (
            .O(N__31212),
            .I(N__31165));
    InMux I__6708 (
            .O(N__31211),
            .I(N__31162));
    InMux I__6707 (
            .O(N__31210),
            .I(N__31157));
    InMux I__6706 (
            .O(N__31209),
            .I(N__31157));
    LocalMux I__6705 (
            .O(N__31200),
            .I(N__31154));
    LocalMux I__6704 (
            .O(N__31197),
            .I(N__31148));
    InMux I__6703 (
            .O(N__31196),
            .I(N__31145));
    InMux I__6702 (
            .O(N__31195),
            .I(N__31140));
    InMux I__6701 (
            .O(N__31194),
            .I(N__31140));
    InMux I__6700 (
            .O(N__31193),
            .I(N__31135));
    InMux I__6699 (
            .O(N__31192),
            .I(N__31135));
    InMux I__6698 (
            .O(N__31191),
            .I(N__31128));
    InMux I__6697 (
            .O(N__31190),
            .I(N__31128));
    InMux I__6696 (
            .O(N__31189),
            .I(N__31128));
    Span4Mux_s0_v I__6695 (
            .O(N__31186),
            .I(N__31125));
    LocalMux I__6694 (
            .O(N__31177),
            .I(N__31119));
    LocalMux I__6693 (
            .O(N__31172),
            .I(N__31119));
    Span4Mux_v I__6692 (
            .O(N__31165),
            .I(N__31114));
    LocalMux I__6691 (
            .O(N__31162),
            .I(N__31114));
    LocalMux I__6690 (
            .O(N__31157),
            .I(N__31111));
    Span4Mux_v I__6689 (
            .O(N__31154),
            .I(N__31108));
    InMux I__6688 (
            .O(N__31153),
            .I(N__31101));
    InMux I__6687 (
            .O(N__31152),
            .I(N__31101));
    InMux I__6686 (
            .O(N__31151),
            .I(N__31101));
    Span4Mux_h I__6685 (
            .O(N__31148),
            .I(N__31088));
    LocalMux I__6684 (
            .O(N__31145),
            .I(N__31088));
    LocalMux I__6683 (
            .O(N__31140),
            .I(N__31088));
    LocalMux I__6682 (
            .O(N__31135),
            .I(N__31088));
    LocalMux I__6681 (
            .O(N__31128),
            .I(N__31088));
    Span4Mux_v I__6680 (
            .O(N__31125),
            .I(N__31088));
    InMux I__6679 (
            .O(N__31124),
            .I(N__31085));
    Span4Mux_v I__6678 (
            .O(N__31119),
            .I(N__31082));
    Span4Mux_v I__6677 (
            .O(N__31114),
            .I(N__31079));
    Span4Mux_h I__6676 (
            .O(N__31111),
            .I(N__31070));
    Span4Mux_h I__6675 (
            .O(N__31108),
            .I(N__31070));
    LocalMux I__6674 (
            .O(N__31101),
            .I(N__31070));
    Span4Mux_v I__6673 (
            .O(N__31088),
            .I(N__31070));
    LocalMux I__6672 (
            .O(N__31085),
            .I(G_146));
    Odrv4 I__6671 (
            .O(N__31082),
            .I(G_146));
    Odrv4 I__6670 (
            .O(N__31079),
            .I(G_146));
    Odrv4 I__6669 (
            .O(N__31070),
            .I(G_146));
    InMux I__6668 (
            .O(N__31061),
            .I(N__31058));
    LocalMux I__6667 (
            .O(N__31058),
            .I(\b2v_inst11.dutycycle_1_0_1 ));
    CascadeMux I__6666 (
            .O(N__31055),
            .I(\b2v_inst11.dutycycle_eena_0_cascade_ ));
    InMux I__6665 (
            .O(N__31052),
            .I(N__31046));
    InMux I__6664 (
            .O(N__31051),
            .I(N__31046));
    LocalMux I__6663 (
            .O(N__31046),
            .I(\b2v_inst11.dutycycleZ1Z_1 ));
    SRMux I__6662 (
            .O(N__31043),
            .I(N__31040));
    LocalMux I__6661 (
            .O(N__31040),
            .I(N__31033));
    SRMux I__6660 (
            .O(N__31039),
            .I(N__31028));
    SRMux I__6659 (
            .O(N__31038),
            .I(N__31025));
    SRMux I__6658 (
            .O(N__31037),
            .I(N__31022));
    SRMux I__6657 (
            .O(N__31036),
            .I(N__31017));
    Span4Mux_h I__6656 (
            .O(N__31033),
            .I(N__31014));
    SRMux I__6655 (
            .O(N__31032),
            .I(N__31011));
    SRMux I__6654 (
            .O(N__31031),
            .I(N__31008));
    LocalMux I__6653 (
            .O(N__31028),
            .I(N__31005));
    LocalMux I__6652 (
            .O(N__31025),
            .I(N__31002));
    LocalMux I__6651 (
            .O(N__31022),
            .I(N__30999));
    SRMux I__6650 (
            .O(N__31021),
            .I(N__30996));
    SRMux I__6649 (
            .O(N__31020),
            .I(N__30993));
    LocalMux I__6648 (
            .O(N__31017),
            .I(N__30990));
    Span4Mux_s2_h I__6647 (
            .O(N__31014),
            .I(N__30985));
    LocalMux I__6646 (
            .O(N__31011),
            .I(N__30985));
    LocalMux I__6645 (
            .O(N__31008),
            .I(N__30981));
    Span4Mux_v I__6644 (
            .O(N__31005),
            .I(N__30978));
    Span4Mux_v I__6643 (
            .O(N__31002),
            .I(N__30975));
    Span4Mux_v I__6642 (
            .O(N__30999),
            .I(N__30970));
    LocalMux I__6641 (
            .O(N__30996),
            .I(N__30970));
    LocalMux I__6640 (
            .O(N__30993),
            .I(N__30967));
    Span4Mux_v I__6639 (
            .O(N__30990),
            .I(N__30964));
    Span4Mux_h I__6638 (
            .O(N__30985),
            .I(N__30961));
    SRMux I__6637 (
            .O(N__30984),
            .I(N__30958));
    Span4Mux_h I__6636 (
            .O(N__30981),
            .I(N__30955));
    Span4Mux_h I__6635 (
            .O(N__30978),
            .I(N__30952));
    Span4Mux_h I__6634 (
            .O(N__30975),
            .I(N__30947));
    Span4Mux_v I__6633 (
            .O(N__30970),
            .I(N__30947));
    Span4Mux_h I__6632 (
            .O(N__30967),
            .I(N__30944));
    Span4Mux_s1_h I__6631 (
            .O(N__30964),
            .I(N__30939));
    Span4Mux_h I__6630 (
            .O(N__30961),
            .I(N__30939));
    LocalMux I__6629 (
            .O(N__30958),
            .I(N__30936));
    Span4Mux_h I__6628 (
            .O(N__30955),
            .I(N__30931));
    Span4Mux_s1_h I__6627 (
            .O(N__30952),
            .I(N__30931));
    Span4Mux_h I__6626 (
            .O(N__30947),
            .I(N__30928));
    Odrv4 I__6625 (
            .O(N__30944),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv4 I__6624 (
            .O(N__30939),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv12 I__6623 (
            .O(N__30936),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv4 I__6622 (
            .O(N__30931),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv4 I__6621 (
            .O(N__30928),
            .I(\b2v_inst11.N_224_iZ0 ));
    CascadeMux I__6620 (
            .O(N__30917),
            .I(\b2v_inst11.count_off_1_0_cascade_ ));
    InMux I__6619 (
            .O(N__30914),
            .I(N__30911));
    LocalMux I__6618 (
            .O(N__30911),
            .I(N__30908));
    Span4Mux_h I__6617 (
            .O(N__30908),
            .I(N__30905));
    Odrv4 I__6616 (
            .O(N__30905),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_330_N ));
    InMux I__6615 (
            .O(N__30902),
            .I(N__30899));
    LocalMux I__6614 (
            .O(N__30899),
            .I(N__30890));
    InMux I__6613 (
            .O(N__30898),
            .I(N__30885));
    InMux I__6612 (
            .O(N__30897),
            .I(N__30885));
    InMux I__6611 (
            .O(N__30896),
            .I(N__30879));
    InMux I__6610 (
            .O(N__30895),
            .I(N__30876));
    InMux I__6609 (
            .O(N__30894),
            .I(N__30871));
    InMux I__6608 (
            .O(N__30893),
            .I(N__30871));
    Span4Mux_v I__6607 (
            .O(N__30890),
            .I(N__30866));
    LocalMux I__6606 (
            .O(N__30885),
            .I(N__30866));
    InMux I__6605 (
            .O(N__30884),
            .I(N__30859));
    InMux I__6604 (
            .O(N__30883),
            .I(N__30859));
    InMux I__6603 (
            .O(N__30882),
            .I(N__30859));
    LocalMux I__6602 (
            .O(N__30879),
            .I(\b2v_inst11.func_state ));
    LocalMux I__6601 (
            .O(N__30876),
            .I(\b2v_inst11.func_state ));
    LocalMux I__6600 (
            .O(N__30871),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__6599 (
            .O(N__30866),
            .I(\b2v_inst11.func_state ));
    LocalMux I__6598 (
            .O(N__30859),
            .I(\b2v_inst11.func_state ));
    InMux I__6597 (
            .O(N__30848),
            .I(N__30845));
    LocalMux I__6596 (
            .O(N__30845),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0 ));
    InMux I__6595 (
            .O(N__30842),
            .I(N__30838));
    InMux I__6594 (
            .O(N__30841),
            .I(N__30835));
    LocalMux I__6593 (
            .O(N__30838),
            .I(N__30832));
    LocalMux I__6592 (
            .O(N__30835),
            .I(\b2v_inst11.N_382 ));
    Odrv12 I__6591 (
            .O(N__30832),
            .I(\b2v_inst11.N_382 ));
    InMux I__6590 (
            .O(N__30827),
            .I(N__30821));
    InMux I__6589 (
            .O(N__30826),
            .I(N__30821));
    LocalMux I__6588 (
            .O(N__30821),
            .I(N__30817));
    InMux I__6587 (
            .O(N__30820),
            .I(N__30814));
    Span4Mux_h I__6586 (
            .O(N__30817),
            .I(N__30811));
    LocalMux I__6585 (
            .O(N__30814),
            .I(N__30808));
    Odrv4 I__6584 (
            .O(N__30811),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_1 ));
    Odrv4 I__6583 (
            .O(N__30808),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_1 ));
    CascadeMux I__6582 (
            .O(N__30803),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ));
    CascadeMux I__6581 (
            .O(N__30800),
            .I(\b2v_inst11.N_315_cascade_ ));
    InMux I__6580 (
            .O(N__30797),
            .I(N__30794));
    LocalMux I__6579 (
            .O(N__30794),
            .I(N__30791));
    Span4Mux_s3_h I__6578 (
            .O(N__30791),
            .I(N__30788));
    Odrv4 I__6577 (
            .O(N__30788),
            .I(\b2v_inst11.count_clk_RNIDQ4A1Z0Z_7 ));
    CascadeMux I__6576 (
            .O(N__30785),
            .I(N__30782));
    InMux I__6575 (
            .O(N__30782),
            .I(N__30779));
    LocalMux I__6574 (
            .O(N__30779),
            .I(N__30774));
    InMux I__6573 (
            .O(N__30778),
            .I(N__30769));
    InMux I__6572 (
            .O(N__30777),
            .I(N__30769));
    Odrv4 I__6571 (
            .O(N__30774),
            .I(\b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2 ));
    LocalMux I__6570 (
            .O(N__30769),
            .I(\b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2 ));
    CascadeMux I__6569 (
            .O(N__30764),
            .I(\b2v_inst11.func_state_1_ss0_i_0_o3_0_cascade_ ));
    InMux I__6568 (
            .O(N__30761),
            .I(N__30758));
    LocalMux I__6567 (
            .O(N__30758),
            .I(N__30754));
    InMux I__6566 (
            .O(N__30757),
            .I(N__30751));
    Span4Mux_v I__6565 (
            .O(N__30754),
            .I(N__30748));
    LocalMux I__6564 (
            .O(N__30751),
            .I(N__30745));
    Span4Mux_h I__6563 (
            .O(N__30748),
            .I(N__30742));
    Span4Mux_h I__6562 (
            .O(N__30745),
            .I(N__30739));
    Odrv4 I__6561 (
            .O(N__30742),
            .I(\b2v_inst11.N_430 ));
    Odrv4 I__6560 (
            .O(N__30739),
            .I(\b2v_inst11.N_430 ));
    InMux I__6559 (
            .O(N__30734),
            .I(N__30719));
    InMux I__6558 (
            .O(N__30733),
            .I(N__30719));
    InMux I__6557 (
            .O(N__30732),
            .I(N__30714));
    InMux I__6556 (
            .O(N__30731),
            .I(N__30714));
    InMux I__6555 (
            .O(N__30730),
            .I(N__30707));
    InMux I__6554 (
            .O(N__30729),
            .I(N__30707));
    InMux I__6553 (
            .O(N__30728),
            .I(N__30707));
    CascadeMux I__6552 (
            .O(N__30727),
            .I(N__30702));
    CascadeMux I__6551 (
            .O(N__30726),
            .I(N__30695));
    CascadeMux I__6550 (
            .O(N__30725),
            .I(N__30685));
    CascadeMux I__6549 (
            .O(N__30724),
            .I(N__30682));
    LocalMux I__6548 (
            .O(N__30719),
            .I(N__30673));
    LocalMux I__6547 (
            .O(N__30714),
            .I(N__30673));
    LocalMux I__6546 (
            .O(N__30707),
            .I(N__30673));
    CascadeMux I__6545 (
            .O(N__30706),
            .I(N__30670));
    CascadeMux I__6544 (
            .O(N__30705),
            .I(N__30667));
    InMux I__6543 (
            .O(N__30702),
            .I(N__30664));
    InMux I__6542 (
            .O(N__30701),
            .I(N__30661));
    InMux I__6541 (
            .O(N__30700),
            .I(N__30658));
    InMux I__6540 (
            .O(N__30699),
            .I(N__30653));
    InMux I__6539 (
            .O(N__30698),
            .I(N__30653));
    InMux I__6538 (
            .O(N__30695),
            .I(N__30644));
    InMux I__6537 (
            .O(N__30694),
            .I(N__30644));
    InMux I__6536 (
            .O(N__30693),
            .I(N__30644));
    InMux I__6535 (
            .O(N__30692),
            .I(N__30644));
    InMux I__6534 (
            .O(N__30691),
            .I(N__30639));
    InMux I__6533 (
            .O(N__30690),
            .I(N__30639));
    CascadeMux I__6532 (
            .O(N__30689),
            .I(N__30628));
    CascadeMux I__6531 (
            .O(N__30688),
            .I(N__30624));
    InMux I__6530 (
            .O(N__30685),
            .I(N__30614));
    InMux I__6529 (
            .O(N__30682),
            .I(N__30614));
    InMux I__6528 (
            .O(N__30681),
            .I(N__30614));
    InMux I__6527 (
            .O(N__30680),
            .I(N__30614));
    Span4Mux_v I__6526 (
            .O(N__30673),
            .I(N__30608));
    InMux I__6525 (
            .O(N__30670),
            .I(N__30605));
    InMux I__6524 (
            .O(N__30667),
            .I(N__30599));
    LocalMux I__6523 (
            .O(N__30664),
            .I(N__30592));
    LocalMux I__6522 (
            .O(N__30661),
            .I(N__30583));
    LocalMux I__6521 (
            .O(N__30658),
            .I(N__30583));
    LocalMux I__6520 (
            .O(N__30653),
            .I(N__30583));
    LocalMux I__6519 (
            .O(N__30644),
            .I(N__30583));
    LocalMux I__6518 (
            .O(N__30639),
            .I(N__30580));
    CascadeMux I__6517 (
            .O(N__30638),
            .I(N__30571));
    InMux I__6516 (
            .O(N__30637),
            .I(N__30568));
    InMux I__6515 (
            .O(N__30636),
            .I(N__30563));
    InMux I__6514 (
            .O(N__30635),
            .I(N__30563));
    InMux I__6513 (
            .O(N__30634),
            .I(N__30560));
    InMux I__6512 (
            .O(N__30633),
            .I(N__30552));
    InMux I__6511 (
            .O(N__30632),
            .I(N__30552));
    InMux I__6510 (
            .O(N__30631),
            .I(N__30549));
    InMux I__6509 (
            .O(N__30628),
            .I(N__30544));
    InMux I__6508 (
            .O(N__30627),
            .I(N__30544));
    InMux I__6507 (
            .O(N__30624),
            .I(N__30540));
    InMux I__6506 (
            .O(N__30623),
            .I(N__30537));
    LocalMux I__6505 (
            .O(N__30614),
            .I(N__30534));
    InMux I__6504 (
            .O(N__30613),
            .I(N__30527));
    InMux I__6503 (
            .O(N__30612),
            .I(N__30527));
    InMux I__6502 (
            .O(N__30611),
            .I(N__30527));
    Span4Mux_h I__6501 (
            .O(N__30608),
            .I(N__30522));
    LocalMux I__6500 (
            .O(N__30605),
            .I(N__30522));
    InMux I__6499 (
            .O(N__30604),
            .I(N__30519));
    InMux I__6498 (
            .O(N__30603),
            .I(N__30516));
    CascadeMux I__6497 (
            .O(N__30602),
            .I(N__30511));
    LocalMux I__6496 (
            .O(N__30599),
            .I(N__30506));
    InMux I__6495 (
            .O(N__30598),
            .I(N__30503));
    InMux I__6494 (
            .O(N__30597),
            .I(N__30496));
    InMux I__6493 (
            .O(N__30596),
            .I(N__30496));
    InMux I__6492 (
            .O(N__30595),
            .I(N__30496));
    Span4Mux_s3_v I__6491 (
            .O(N__30592),
            .I(N__30489));
    Span4Mux_s3_v I__6490 (
            .O(N__30583),
            .I(N__30489));
    Span4Mux_s3_v I__6489 (
            .O(N__30580),
            .I(N__30489));
    InMux I__6488 (
            .O(N__30579),
            .I(N__30482));
    InMux I__6487 (
            .O(N__30578),
            .I(N__30482));
    InMux I__6486 (
            .O(N__30577),
            .I(N__30482));
    InMux I__6485 (
            .O(N__30576),
            .I(N__30477));
    InMux I__6484 (
            .O(N__30575),
            .I(N__30477));
    InMux I__6483 (
            .O(N__30574),
            .I(N__30474));
    InMux I__6482 (
            .O(N__30571),
            .I(N__30471));
    LocalMux I__6481 (
            .O(N__30568),
            .I(N__30464));
    LocalMux I__6480 (
            .O(N__30563),
            .I(N__30464));
    LocalMux I__6479 (
            .O(N__30560),
            .I(N__30464));
    InMux I__6478 (
            .O(N__30559),
            .I(N__30457));
    InMux I__6477 (
            .O(N__30558),
            .I(N__30457));
    InMux I__6476 (
            .O(N__30557),
            .I(N__30457));
    LocalMux I__6475 (
            .O(N__30552),
            .I(N__30454));
    LocalMux I__6474 (
            .O(N__30549),
            .I(N__30451));
    LocalMux I__6473 (
            .O(N__30544),
            .I(N__30448));
    InMux I__6472 (
            .O(N__30543),
            .I(N__30445));
    LocalMux I__6471 (
            .O(N__30540),
            .I(N__30442));
    LocalMux I__6470 (
            .O(N__30537),
            .I(N__30429));
    Span4Mux_s1_v I__6469 (
            .O(N__30534),
            .I(N__30429));
    LocalMux I__6468 (
            .O(N__30527),
            .I(N__30429));
    Span4Mux_h I__6467 (
            .O(N__30522),
            .I(N__30429));
    LocalMux I__6466 (
            .O(N__30519),
            .I(N__30429));
    LocalMux I__6465 (
            .O(N__30516),
            .I(N__30429));
    InMux I__6464 (
            .O(N__30515),
            .I(N__30424));
    InMux I__6463 (
            .O(N__30514),
            .I(N__30424));
    InMux I__6462 (
            .O(N__30511),
            .I(N__30421));
    InMux I__6461 (
            .O(N__30510),
            .I(N__30415));
    InMux I__6460 (
            .O(N__30509),
            .I(N__30415));
    Span4Mux_v I__6459 (
            .O(N__30506),
            .I(N__30410));
    LocalMux I__6458 (
            .O(N__30503),
            .I(N__30410));
    LocalMux I__6457 (
            .O(N__30496),
            .I(N__30407));
    Sp12to4 I__6456 (
            .O(N__30489),
            .I(N__30402));
    LocalMux I__6455 (
            .O(N__30482),
            .I(N__30402));
    LocalMux I__6454 (
            .O(N__30477),
            .I(N__30399));
    LocalMux I__6453 (
            .O(N__30474),
            .I(N__30392));
    LocalMux I__6452 (
            .O(N__30471),
            .I(N__30392));
    Sp12to4 I__6451 (
            .O(N__30464),
            .I(N__30392));
    LocalMux I__6450 (
            .O(N__30457),
            .I(N__30388));
    Span4Mux_s2_v I__6449 (
            .O(N__30454),
            .I(N__30379));
    Span4Mux_v I__6448 (
            .O(N__30451),
            .I(N__30379));
    Span4Mux_h I__6447 (
            .O(N__30448),
            .I(N__30379));
    LocalMux I__6446 (
            .O(N__30445),
            .I(N__30379));
    Span4Mux_h I__6445 (
            .O(N__30442),
            .I(N__30372));
    Span4Mux_v I__6444 (
            .O(N__30429),
            .I(N__30372));
    LocalMux I__6443 (
            .O(N__30424),
            .I(N__30372));
    LocalMux I__6442 (
            .O(N__30421),
            .I(N__30369));
    InMux I__6441 (
            .O(N__30420),
            .I(N__30366));
    LocalMux I__6440 (
            .O(N__30415),
            .I(N__30361));
    Span4Mux_v I__6439 (
            .O(N__30410),
            .I(N__30361));
    Span4Mux_s3_h I__6438 (
            .O(N__30407),
            .I(N__30358));
    Span12Mux_s7_h I__6437 (
            .O(N__30402),
            .I(N__30351));
    Span12Mux_s7_h I__6436 (
            .O(N__30399),
            .I(N__30351));
    Span12Mux_s3_v I__6435 (
            .O(N__30392),
            .I(N__30351));
    InMux I__6434 (
            .O(N__30391),
            .I(N__30348));
    Span4Mux_s2_v I__6433 (
            .O(N__30388),
            .I(N__30337));
    Span4Mux_h I__6432 (
            .O(N__30379),
            .I(N__30337));
    Span4Mux_v I__6431 (
            .O(N__30372),
            .I(N__30337));
    Span4Mux_s3_h I__6430 (
            .O(N__30369),
            .I(N__30337));
    LocalMux I__6429 (
            .O(N__30366),
            .I(N__30337));
    Odrv4 I__6428 (
            .O(N__30361),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__6427 (
            .O(N__30358),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv12 I__6426 (
            .O(N__30351),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__6425 (
            .O(N__30348),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__6424 (
            .O(N__30337),
            .I(SYNTHESIZED_WIRE_1keep_3));
    CascadeMux I__6423 (
            .O(N__30326),
            .I(N__30321));
    CascadeMux I__6422 (
            .O(N__30325),
            .I(N__30318));
    InMux I__6421 (
            .O(N__30324),
            .I(N__30315));
    InMux I__6420 (
            .O(N__30321),
            .I(N__30310));
    InMux I__6419 (
            .O(N__30318),
            .I(N__30310));
    LocalMux I__6418 (
            .O(N__30315),
            .I(N__30303));
    LocalMux I__6417 (
            .O(N__30310),
            .I(N__30300));
    InMux I__6416 (
            .O(N__30309),
            .I(N__30297));
    InMux I__6415 (
            .O(N__30308),
            .I(N__30294));
    CascadeMux I__6414 (
            .O(N__30307),
            .I(N__30291));
    CascadeMux I__6413 (
            .O(N__30306),
            .I(N__30287));
    Span4Mux_v I__6412 (
            .O(N__30303),
            .I(N__30283));
    Span4Mux_s2_h I__6411 (
            .O(N__30300),
            .I(N__30278));
    LocalMux I__6410 (
            .O(N__30297),
            .I(N__30278));
    LocalMux I__6409 (
            .O(N__30294),
            .I(N__30272));
    InMux I__6408 (
            .O(N__30291),
            .I(N__30265));
    InMux I__6407 (
            .O(N__30290),
            .I(N__30265));
    InMux I__6406 (
            .O(N__30287),
            .I(N__30265));
    InMux I__6405 (
            .O(N__30286),
            .I(N__30262));
    Sp12to4 I__6404 (
            .O(N__30283),
            .I(N__30259));
    Span4Mux_h I__6403 (
            .O(N__30278),
            .I(N__30256));
    InMux I__6402 (
            .O(N__30277),
            .I(N__30251));
    InMux I__6401 (
            .O(N__30276),
            .I(N__30251));
    InMux I__6400 (
            .O(N__30275),
            .I(N__30248));
    Span4Mux_v I__6399 (
            .O(N__30272),
            .I(N__30241));
    LocalMux I__6398 (
            .O(N__30265),
            .I(N__30241));
    LocalMux I__6397 (
            .O(N__30262),
            .I(N__30241));
    Odrv12 I__6396 (
            .O(N__30259),
            .I(\b2v_inst11.N_161 ));
    Odrv4 I__6395 (
            .O(N__30256),
            .I(\b2v_inst11.N_161 ));
    LocalMux I__6394 (
            .O(N__30251),
            .I(\b2v_inst11.N_161 ));
    LocalMux I__6393 (
            .O(N__30248),
            .I(\b2v_inst11.N_161 ));
    Odrv4 I__6392 (
            .O(N__30241),
            .I(\b2v_inst11.N_161 ));
    InMux I__6391 (
            .O(N__30230),
            .I(N__30227));
    LocalMux I__6390 (
            .O(N__30227),
            .I(\b2v_inst11.N_339 ));
    InMux I__6389 (
            .O(N__30224),
            .I(N__30221));
    LocalMux I__6388 (
            .O(N__30221),
            .I(N__30218));
    Span4Mux_s2_h I__6387 (
            .O(N__30218),
            .I(N__30215));
    Span4Mux_v I__6386 (
            .O(N__30215),
            .I(N__30212));
    Odrv4 I__6385 (
            .O(N__30212),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ));
    CascadeMux I__6384 (
            .O(N__30209),
            .I(\b2v_inst11.dutycycle_1_0_1_cascade_ ));
    InMux I__6383 (
            .O(N__30206),
            .I(N__30203));
    LocalMux I__6382 (
            .O(N__30203),
            .I(\b2v_inst11.dutycycle_eena ));
    CascadeMux I__6381 (
            .O(N__30200),
            .I(N__30197));
    InMux I__6380 (
            .O(N__30197),
            .I(N__30191));
    InMux I__6379 (
            .O(N__30196),
            .I(N__30191));
    LocalMux I__6378 (
            .O(N__30191),
            .I(\b2v_inst11.dutycycleZ1Z_0 ));
    CascadeMux I__6377 (
            .O(N__30188),
            .I(\b2v_inst11.dutycycle_eena_cascade_ ));
    CascadeMux I__6376 (
            .O(N__30185),
            .I(N__30180));
    CascadeMux I__6375 (
            .O(N__30184),
            .I(N__30177));
    InMux I__6374 (
            .O(N__30183),
            .I(N__30172));
    InMux I__6373 (
            .O(N__30180),
            .I(N__30169));
    InMux I__6372 (
            .O(N__30177),
            .I(N__30161));
    InMux I__6371 (
            .O(N__30176),
            .I(N__30161));
    CascadeMux I__6370 (
            .O(N__30175),
            .I(N__30158));
    LocalMux I__6369 (
            .O(N__30172),
            .I(N__30155));
    LocalMux I__6368 (
            .O(N__30169),
            .I(N__30151));
    InMux I__6367 (
            .O(N__30168),
            .I(N__30148));
    InMux I__6366 (
            .O(N__30167),
            .I(N__30145));
    CascadeMux I__6365 (
            .O(N__30166),
            .I(N__30139));
    LocalMux I__6364 (
            .O(N__30161),
            .I(N__30136));
    InMux I__6363 (
            .O(N__30158),
            .I(N__30133));
    Span4Mux_s1_v I__6362 (
            .O(N__30155),
            .I(N__30130));
    InMux I__6361 (
            .O(N__30154),
            .I(N__30127));
    Span4Mux_v I__6360 (
            .O(N__30151),
            .I(N__30119));
    LocalMux I__6359 (
            .O(N__30148),
            .I(N__30119));
    LocalMux I__6358 (
            .O(N__30145),
            .I(N__30119));
    CascadeMux I__6357 (
            .O(N__30144),
            .I(N__30116));
    InMux I__6356 (
            .O(N__30143),
            .I(N__30112));
    InMux I__6355 (
            .O(N__30142),
            .I(N__30107));
    InMux I__6354 (
            .O(N__30139),
            .I(N__30107));
    Span4Mux_v I__6353 (
            .O(N__30136),
            .I(N__30102));
    LocalMux I__6352 (
            .O(N__30133),
            .I(N__30102));
    Span4Mux_h I__6351 (
            .O(N__30130),
            .I(N__30097));
    LocalMux I__6350 (
            .O(N__30127),
            .I(N__30097));
    InMux I__6349 (
            .O(N__30126),
            .I(N__30094));
    Span4Mux_v I__6348 (
            .O(N__30119),
            .I(N__30091));
    InMux I__6347 (
            .O(N__30116),
            .I(N__30088));
    InMux I__6346 (
            .O(N__30115),
            .I(N__30085));
    LocalMux I__6345 (
            .O(N__30112),
            .I(N__30078));
    LocalMux I__6344 (
            .O(N__30107),
            .I(N__30078));
    Span4Mux_h I__6343 (
            .O(N__30102),
            .I(N__30078));
    Span4Mux_v I__6342 (
            .O(N__30097),
            .I(N__30073));
    LocalMux I__6341 (
            .O(N__30094),
            .I(N__30073));
    Span4Mux_h I__6340 (
            .O(N__30091),
            .I(N__30068));
    LocalMux I__6339 (
            .O(N__30088),
            .I(N__30068));
    LocalMux I__6338 (
            .O(N__30085),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__6337 (
            .O(N__30078),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__6336 (
            .O(N__30073),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__6335 (
            .O(N__30068),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    CascadeMux I__6334 (
            .O(N__30059),
            .I(\b2v_inst11.dutycycleZ0Z_0_cascade_ ));
    InMux I__6333 (
            .O(N__30056),
            .I(N__30050));
    InMux I__6332 (
            .O(N__30055),
            .I(N__30050));
    LocalMux I__6331 (
            .O(N__30050),
            .I(\b2v_inst11.dutycycle_1_0_0 ));
    InMux I__6330 (
            .O(N__30047),
            .I(N__30044));
    LocalMux I__6329 (
            .O(N__30044),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2 ));
    CascadeMux I__6328 (
            .O(N__30041),
            .I(\b2v_inst11.dutycycleZ0Z_2_cascade_ ));
    InMux I__6327 (
            .O(N__30038),
            .I(N__30035));
    LocalMux I__6326 (
            .O(N__30035),
            .I(N__30032));
    Span4Mux_h I__6325 (
            .O(N__30032),
            .I(N__30029));
    Span4Mux_h I__6324 (
            .O(N__30029),
            .I(N__30026));
    Span4Mux_v I__6323 (
            .O(N__30026),
            .I(N__30023));
    Odrv4 I__6322 (
            .O(N__30023),
            .I(\b2v_inst11.mult1_un152_sum_i ));
    CascadeMux I__6321 (
            .O(N__30020),
            .I(N__30016));
    InMux I__6320 (
            .O(N__30019),
            .I(N__30011));
    InMux I__6319 (
            .O(N__30016),
            .I(N__30011));
    LocalMux I__6318 (
            .O(N__30011),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_0_2 ));
    InMux I__6317 (
            .O(N__30008),
            .I(N__30002));
    InMux I__6316 (
            .O(N__30007),
            .I(N__30002));
    LocalMux I__6315 (
            .O(N__30002),
            .I(N__29999));
    Odrv4 I__6314 (
            .O(N__29999),
            .I(\b2v_inst11.N_168 ));
    InMux I__6313 (
            .O(N__29996),
            .I(N__29990));
    InMux I__6312 (
            .O(N__29995),
            .I(N__29990));
    LocalMux I__6311 (
            .O(N__29990),
            .I(N__29987));
    Odrv4 I__6310 (
            .O(N__29987),
            .I(\b2v_inst11.dutycycle_RNIAEUL3Z0Z_2 ));
    CascadeMux I__6309 (
            .O(N__29984),
            .I(N__29981));
    InMux I__6308 (
            .O(N__29981),
            .I(N__29975));
    InMux I__6307 (
            .O(N__29980),
            .I(N__29975));
    LocalMux I__6306 (
            .O(N__29975),
            .I(\b2v_inst11.dutycycleZ1Z_2 ));
    InMux I__6305 (
            .O(N__29972),
            .I(N__29958));
    CascadeMux I__6304 (
            .O(N__29971),
            .I(N__29954));
    InMux I__6303 (
            .O(N__29970),
            .I(N__29948));
    InMux I__6302 (
            .O(N__29969),
            .I(N__29948));
    InMux I__6301 (
            .O(N__29968),
            .I(N__29943));
    InMux I__6300 (
            .O(N__29967),
            .I(N__29943));
    InMux I__6299 (
            .O(N__29966),
            .I(N__29938));
    InMux I__6298 (
            .O(N__29965),
            .I(N__29935));
    InMux I__6297 (
            .O(N__29964),
            .I(N__29932));
    InMux I__6296 (
            .O(N__29963),
            .I(N__29927));
    InMux I__6295 (
            .O(N__29962),
            .I(N__29927));
    InMux I__6294 (
            .O(N__29961),
            .I(N__29923));
    LocalMux I__6293 (
            .O(N__29958),
            .I(N__29920));
    InMux I__6292 (
            .O(N__29957),
            .I(N__29917));
    InMux I__6291 (
            .O(N__29954),
            .I(N__29912));
    InMux I__6290 (
            .O(N__29953),
            .I(N__29912));
    LocalMux I__6289 (
            .O(N__29948),
            .I(N__29907));
    LocalMux I__6288 (
            .O(N__29943),
            .I(N__29907));
    InMux I__6287 (
            .O(N__29942),
            .I(N__29903));
    InMux I__6286 (
            .O(N__29941),
            .I(N__29900));
    LocalMux I__6285 (
            .O(N__29938),
            .I(N__29897));
    LocalMux I__6284 (
            .O(N__29935),
            .I(N__29892));
    LocalMux I__6283 (
            .O(N__29932),
            .I(N__29892));
    LocalMux I__6282 (
            .O(N__29927),
            .I(N__29887));
    InMux I__6281 (
            .O(N__29926),
            .I(N__29883));
    LocalMux I__6280 (
            .O(N__29923),
            .I(N__29878));
    Span4Mux_v I__6279 (
            .O(N__29920),
            .I(N__29878));
    LocalMux I__6278 (
            .O(N__29917),
            .I(N__29871));
    LocalMux I__6277 (
            .O(N__29912),
            .I(N__29871));
    Span4Mux_h I__6276 (
            .O(N__29907),
            .I(N__29871));
    InMux I__6275 (
            .O(N__29906),
            .I(N__29868));
    LocalMux I__6274 (
            .O(N__29903),
            .I(N__29865));
    LocalMux I__6273 (
            .O(N__29900),
            .I(N__29858));
    Span4Mux_v I__6272 (
            .O(N__29897),
            .I(N__29858));
    Span4Mux_h I__6271 (
            .O(N__29892),
            .I(N__29858));
    InMux I__6270 (
            .O(N__29891),
            .I(N__29855));
    InMux I__6269 (
            .O(N__29890),
            .I(N__29852));
    Span4Mux_v I__6268 (
            .O(N__29887),
            .I(N__29849));
    InMux I__6267 (
            .O(N__29886),
            .I(N__29846));
    LocalMux I__6266 (
            .O(N__29883),
            .I(N__29841));
    Span4Mux_h I__6265 (
            .O(N__29878),
            .I(N__29841));
    Span4Mux_v I__6264 (
            .O(N__29871),
            .I(N__29838));
    LocalMux I__6263 (
            .O(N__29868),
            .I(N__29835));
    Span4Mux_v I__6262 (
            .O(N__29865),
            .I(N__29826));
    Span4Mux_v I__6261 (
            .O(N__29858),
            .I(N__29826));
    LocalMux I__6260 (
            .O(N__29855),
            .I(N__29826));
    LocalMux I__6259 (
            .O(N__29852),
            .I(N__29826));
    Odrv4 I__6258 (
            .O(N__29849),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    LocalMux I__6257 (
            .O(N__29846),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__6256 (
            .O(N__29841),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__6255 (
            .O(N__29838),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv12 I__6254 (
            .O(N__29835),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__6253 (
            .O(N__29826),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    CascadeMux I__6252 (
            .O(N__29813),
            .I(N__29810));
    InMux I__6251 (
            .O(N__29810),
            .I(N__29804));
    InMux I__6250 (
            .O(N__29809),
            .I(N__29804));
    LocalMux I__6249 (
            .O(N__29804),
            .I(N__29801));
    Span4Mux_v I__6248 (
            .O(N__29801),
            .I(N__29798));
    Sp12to4 I__6247 (
            .O(N__29798),
            .I(N__29794));
    InMux I__6246 (
            .O(N__29797),
            .I(N__29791));
    Odrv12 I__6245 (
            .O(N__29794),
            .I(\b2v_inst11.N_365 ));
    LocalMux I__6244 (
            .O(N__29791),
            .I(\b2v_inst11.N_365 ));
    InMux I__6243 (
            .O(N__29786),
            .I(N__29783));
    LocalMux I__6242 (
            .O(N__29783),
            .I(N__29780));
    Span4Mux_v I__6241 (
            .O(N__29780),
            .I(N__29777));
    Span4Mux_h I__6240 (
            .O(N__29777),
            .I(N__29774));
    Odrv4 I__6239 (
            .O(N__29774),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1 ));
    CascadeMux I__6238 (
            .O(N__29771),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1_cascade_ ));
    InMux I__6237 (
            .O(N__29768),
            .I(N__29765));
    LocalMux I__6236 (
            .O(N__29765),
            .I(N__29762));
    Span4Mux_v I__6235 (
            .O(N__29762),
            .I(N__29759));
    Odrv4 I__6234 (
            .O(N__29759),
            .I(\b2v_inst11.N_186_i ));
    InMux I__6233 (
            .O(N__29756),
            .I(N__29750));
    InMux I__6232 (
            .O(N__29755),
            .I(N__29743));
    InMux I__6231 (
            .O(N__29754),
            .I(N__29743));
    InMux I__6230 (
            .O(N__29753),
            .I(N__29743));
    LocalMux I__6229 (
            .O(N__29750),
            .I(N__29738));
    LocalMux I__6228 (
            .O(N__29743),
            .I(N__29738));
    Span4Mux_v I__6227 (
            .O(N__29738),
            .I(N__29735));
    Span4Mux_h I__6226 (
            .O(N__29735),
            .I(N__29732));
    Odrv4 I__6225 (
            .O(N__29732),
            .I(\b2v_inst6.N_192 ));
    InMux I__6224 (
            .O(N__29729),
            .I(N__29726));
    LocalMux I__6223 (
            .O(N__29726),
            .I(N__29722));
    InMux I__6222 (
            .O(N__29725),
            .I(N__29719));
    Odrv12 I__6221 (
            .O(N__29722),
            .I(N_241));
    LocalMux I__6220 (
            .O(N__29719),
            .I(N_241));
    InMux I__6219 (
            .O(N__29714),
            .I(N__29708));
    InMux I__6218 (
            .O(N__29713),
            .I(N__29708));
    LocalMux I__6217 (
            .O(N__29708),
            .I(\b2v_inst6.N_276_0 ));
    CascadeMux I__6216 (
            .O(N__29705),
            .I(N__29701));
    CascadeMux I__6215 (
            .O(N__29704),
            .I(N__29698));
    InMux I__6214 (
            .O(N__29701),
            .I(N__29694));
    InMux I__6213 (
            .O(N__29698),
            .I(N__29691));
    InMux I__6212 (
            .O(N__29697),
            .I(N__29688));
    LocalMux I__6211 (
            .O(N__29694),
            .I(\b2v_inst6.curr_state_RNIUP4B1Z0Z_0 ));
    LocalMux I__6210 (
            .O(N__29691),
            .I(\b2v_inst6.curr_state_RNIUP4B1Z0Z_0 ));
    LocalMux I__6209 (
            .O(N__29688),
            .I(\b2v_inst6.curr_state_RNIUP4B1Z0Z_0 ));
    InMux I__6208 (
            .O(N__29681),
            .I(N__29675));
    InMux I__6207 (
            .O(N__29680),
            .I(N__29675));
    LocalMux I__6206 (
            .O(N__29675),
            .I(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ));
    InMux I__6205 (
            .O(N__29672),
            .I(N__29669));
    LocalMux I__6204 (
            .O(N__29669),
            .I(N__29666));
    Span4Mux_v I__6203 (
            .O(N__29666),
            .I(N__29663));
    Span4Mux_h I__6202 (
            .O(N__29663),
            .I(N__29660));
    Odrv4 I__6201 (
            .O(N__29660),
            .I(\b2v_inst11.N_9 ));
    CascadeMux I__6200 (
            .O(N__29657),
            .I(\b2v_inst11.N_172_cascade_ ));
    InMux I__6199 (
            .O(N__29654),
            .I(N__29651));
    LocalMux I__6198 (
            .O(N__29651),
            .I(N__29648));
    Span4Mux_v I__6197 (
            .O(N__29648),
            .I(N__29645));
    Odrv4 I__6196 (
            .O(N__29645),
            .I(\b2v_inst11.g0_i_a7_1_3 ));
    CascadeMux I__6195 (
            .O(N__29642),
            .I(\b2v_inst11.g0_i_0_cascade_ ));
    InMux I__6194 (
            .O(N__29639),
            .I(N__29631));
    InMux I__6193 (
            .O(N__29638),
            .I(N__29631));
    CascadeMux I__6192 (
            .O(N__29637),
            .I(N__29628));
    InMux I__6191 (
            .O(N__29636),
            .I(N__29625));
    LocalMux I__6190 (
            .O(N__29631),
            .I(N__29620));
    InMux I__6189 (
            .O(N__29628),
            .I(N__29617));
    LocalMux I__6188 (
            .O(N__29625),
            .I(N__29614));
    InMux I__6187 (
            .O(N__29624),
            .I(N__29609));
    InMux I__6186 (
            .O(N__29623),
            .I(N__29609));
    Sp12to4 I__6185 (
            .O(N__29620),
            .I(N__29602));
    LocalMux I__6184 (
            .O(N__29617),
            .I(N__29602));
    Span4Mux_s3_h I__6183 (
            .O(N__29614),
            .I(N__29597));
    LocalMux I__6182 (
            .O(N__29609),
            .I(N__29597));
    InMux I__6181 (
            .O(N__29608),
            .I(N__29592));
    InMux I__6180 (
            .O(N__29607),
            .I(N__29592));
    Odrv12 I__6179 (
            .O(N__29602),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    Odrv4 I__6178 (
            .O(N__29597),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    LocalMux I__6177 (
            .O(N__29592),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    InMux I__6176 (
            .O(N__29585),
            .I(N__29582));
    LocalMux I__6175 (
            .O(N__29582),
            .I(N__29579));
    Span4Mux_h I__6174 (
            .O(N__29579),
            .I(N__29576));
    Odrv4 I__6173 (
            .O(N__29576),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8 ));
    CascadeMux I__6172 (
            .O(N__29573),
            .I(\b2v_inst11.N_295_cascade_ ));
    InMux I__6171 (
            .O(N__29570),
            .I(N__29567));
    LocalMux I__6170 (
            .O(N__29567),
            .I(N__29564));
    Odrv12 I__6169 (
            .O(N__29564),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3_out ));
    InMux I__6168 (
            .O(N__29561),
            .I(N__29558));
    LocalMux I__6167 (
            .O(N__29558),
            .I(N__29555));
    Span4Mux_v I__6166 (
            .O(N__29555),
            .I(N__29552));
    Span4Mux_h I__6165 (
            .O(N__29552),
            .I(N__29549));
    Odrv4 I__6164 (
            .O(N__29549),
            .I(\b2v_inst11.N_355 ));
    InMux I__6163 (
            .O(N__29546),
            .I(N__29543));
    LocalMux I__6162 (
            .O(N__29543),
            .I(\b2v_inst6.curr_state_1_1 ));
    CascadeMux I__6161 (
            .O(N__29540),
            .I(\b2v_inst6.N_42_cascade_ ));
    InMux I__6160 (
            .O(N__29537),
            .I(N__29530));
    InMux I__6159 (
            .O(N__29536),
            .I(N__29530));
    InMux I__6158 (
            .O(N__29535),
            .I(N__29527));
    LocalMux I__6157 (
            .O(N__29530),
            .I(\b2v_inst6.curr_stateZ0Z_1 ));
    LocalMux I__6156 (
            .O(N__29527),
            .I(\b2v_inst6.curr_stateZ0Z_1 ));
    CascadeMux I__6155 (
            .O(N__29522),
            .I(\b2v_inst6.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__6154 (
            .O(N__29519),
            .I(\b2v_inst6.N_3053_i_cascade_ ));
    InMux I__6153 (
            .O(N__29516),
            .I(N__29511));
    InMux I__6152 (
            .O(N__29515),
            .I(N__29506));
    InMux I__6151 (
            .O(N__29514),
            .I(N__29506));
    LocalMux I__6150 (
            .O(N__29511),
            .I(\b2v_inst6.N_3034_i ));
    LocalMux I__6149 (
            .O(N__29506),
            .I(\b2v_inst6.N_3034_i ));
    CascadeMux I__6148 (
            .O(N__29501),
            .I(\b2v_inst6.N_3034_i_cascade_ ));
    CascadeMux I__6147 (
            .O(N__29498),
            .I(\b2v_inst6.curr_state_RNIUP4B1Z0Z_0_cascade_ ));
    CascadeMux I__6146 (
            .O(N__29495),
            .I(\b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ));
    InMux I__6145 (
            .O(N__29492),
            .I(N__29484));
    InMux I__6144 (
            .O(N__29491),
            .I(N__29477));
    InMux I__6143 (
            .O(N__29490),
            .I(N__29477));
    InMux I__6142 (
            .O(N__29489),
            .I(N__29477));
    InMux I__6141 (
            .O(N__29488),
            .I(N__29472));
    InMux I__6140 (
            .O(N__29487),
            .I(N__29472));
    LocalMux I__6139 (
            .O(N__29484),
            .I(N__29465));
    LocalMux I__6138 (
            .O(N__29477),
            .I(N__29465));
    LocalMux I__6137 (
            .O(N__29472),
            .I(N__29465));
    Span4Mux_s2_v I__6136 (
            .O(N__29465),
            .I(N__29462));
    Span4Mux_v I__6135 (
            .O(N__29462),
            .I(N__29459));
    Span4Mux_h I__6134 (
            .O(N__29459),
            .I(N__29456));
    Odrv4 I__6133 (
            .O(N__29456),
            .I(N_222));
    InMux I__6132 (
            .O(N__29453),
            .I(N__29444));
    InMux I__6131 (
            .O(N__29452),
            .I(N__29444));
    InMux I__6130 (
            .O(N__29451),
            .I(N__29444));
    LocalMux I__6129 (
            .O(N__29444),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    CascadeMux I__6128 (
            .O(N__29441),
            .I(N__29437));
    InMux I__6127 (
            .O(N__29440),
            .I(N__29429));
    InMux I__6126 (
            .O(N__29437),
            .I(N__29429));
    InMux I__6125 (
            .O(N__29436),
            .I(N__29429));
    LocalMux I__6124 (
            .O(N__29429),
            .I(\b2v_inst6.N_3053_i ));
    CascadeMux I__6123 (
            .O(N__29426),
            .I(N__29422));
    InMux I__6122 (
            .O(N__29425),
            .I(N__29419));
    InMux I__6121 (
            .O(N__29422),
            .I(N__29416));
    LocalMux I__6120 (
            .O(N__29419),
            .I(N__29413));
    LocalMux I__6119 (
            .O(N__29416),
            .I(\b2v_inst6.un2_count_1_axb_9 ));
    Odrv4 I__6118 (
            .O(N__29413),
            .I(\b2v_inst6.un2_count_1_axb_9 ));
    InMux I__6117 (
            .O(N__29408),
            .I(N__29402));
    InMux I__6116 (
            .O(N__29407),
            .I(N__29402));
    LocalMux I__6115 (
            .O(N__29402),
            .I(N__29399));
    Odrv12 I__6114 (
            .O(N__29399),
            .I(\b2v_inst6.un2_count_1_cry_8_THRU_CO ));
    CascadeMux I__6113 (
            .O(N__29396),
            .I(\b2v_inst6.un2_count_1_axb_9_cascade_ ));
    CascadeMux I__6112 (
            .O(N__29393),
            .I(\b2v_inst6.count_rst_6_cascade_ ));
    CascadeMux I__6111 (
            .O(N__29390),
            .I(N__29386));
    InMux I__6110 (
            .O(N__29389),
            .I(N__29381));
    InMux I__6109 (
            .O(N__29386),
            .I(N__29381));
    LocalMux I__6108 (
            .O(N__29381),
            .I(N__29378));
    Odrv12 I__6107 (
            .O(N__29378),
            .I(\b2v_inst6.un2_count_1_cry_7_THRU_CO ));
    CascadeMux I__6106 (
            .O(N__29375),
            .I(\b2v_inst6.countZ0Z_8_cascade_ ));
    InMux I__6105 (
            .O(N__29372),
            .I(N__29369));
    LocalMux I__6104 (
            .O(N__29369),
            .I(N__29366));
    Odrv4 I__6103 (
            .O(N__29366),
            .I(\b2v_inst6.count_0_8 ));
    InMux I__6102 (
            .O(N__29363),
            .I(N__29360));
    LocalMux I__6101 (
            .O(N__29360),
            .I(\b2v_inst6.curr_state_1_0 ));
    CascadeMux I__6100 (
            .O(N__29357),
            .I(\b2v_inst6.curr_state_7_0_cascade_ ));
    InMux I__6099 (
            .O(N__29354),
            .I(N__29351));
    LocalMux I__6098 (
            .O(N__29351),
            .I(\b2v_inst6.N_42 ));
    CascadeMux I__6097 (
            .O(N__29348),
            .I(\b2v_inst6.countZ0Z_6_cascade_ ));
    CascadeMux I__6096 (
            .O(N__29345),
            .I(\b2v_inst6.count_1_i_a3_0_0_cascade_ ));
    InMux I__6095 (
            .O(N__29342),
            .I(N__29338));
    InMux I__6094 (
            .O(N__29341),
            .I(N__29335));
    LocalMux I__6093 (
            .O(N__29338),
            .I(N__29330));
    LocalMux I__6092 (
            .O(N__29335),
            .I(N__29327));
    CascadeMux I__6091 (
            .O(N__29334),
            .I(N__29322));
    CascadeMux I__6090 (
            .O(N__29333),
            .I(N__29319));
    Sp12to4 I__6089 (
            .O(N__29330),
            .I(N__29315));
    Span4Mux_s2_h I__6088 (
            .O(N__29327),
            .I(N__29312));
    InMux I__6087 (
            .O(N__29326),
            .I(N__29301));
    InMux I__6086 (
            .O(N__29325),
            .I(N__29301));
    InMux I__6085 (
            .O(N__29322),
            .I(N__29301));
    InMux I__6084 (
            .O(N__29319),
            .I(N__29301));
    InMux I__6083 (
            .O(N__29318),
            .I(N__29301));
    Odrv12 I__6082 (
            .O(N__29315),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    Odrv4 I__6081 (
            .O(N__29312),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    LocalMux I__6080 (
            .O(N__29301),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    InMux I__6079 (
            .O(N__29294),
            .I(N__29289));
    CascadeMux I__6078 (
            .O(N__29293),
            .I(N__29286));
    InMux I__6077 (
            .O(N__29292),
            .I(N__29279));
    LocalMux I__6076 (
            .O(N__29289),
            .I(N__29276));
    InMux I__6075 (
            .O(N__29286),
            .I(N__29273));
    InMux I__6074 (
            .O(N__29285),
            .I(N__29264));
    InMux I__6073 (
            .O(N__29284),
            .I(N__29264));
    InMux I__6072 (
            .O(N__29283),
            .I(N__29264));
    InMux I__6071 (
            .O(N__29282),
            .I(N__29264));
    LocalMux I__6070 (
            .O(N__29279),
            .I(N__29261));
    Span4Mux_v I__6069 (
            .O(N__29276),
            .I(N__29252));
    LocalMux I__6068 (
            .O(N__29273),
            .I(N__29252));
    LocalMux I__6067 (
            .O(N__29264),
            .I(N__29252));
    Span4Mux_v I__6066 (
            .O(N__29261),
            .I(N__29252));
    Odrv4 I__6065 (
            .O(N__29252),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    InMux I__6064 (
            .O(N__29249),
            .I(N__29239));
    InMux I__6063 (
            .O(N__29248),
            .I(N__29228));
    InMux I__6062 (
            .O(N__29247),
            .I(N__29228));
    InMux I__6061 (
            .O(N__29246),
            .I(N__29228));
    InMux I__6060 (
            .O(N__29245),
            .I(N__29228));
    InMux I__6059 (
            .O(N__29244),
            .I(N__29228));
    CascadeMux I__6058 (
            .O(N__29243),
            .I(N__29225));
    InMux I__6057 (
            .O(N__29242),
            .I(N__29222));
    LocalMux I__6056 (
            .O(N__29239),
            .I(N__29217));
    LocalMux I__6055 (
            .O(N__29228),
            .I(N__29217));
    InMux I__6054 (
            .O(N__29225),
            .I(N__29214));
    LocalMux I__6053 (
            .O(N__29222),
            .I(N__29211));
    Span4Mux_h I__6052 (
            .O(N__29217),
            .I(N__29206));
    LocalMux I__6051 (
            .O(N__29214),
            .I(N__29206));
    Span4Mux_h I__6050 (
            .O(N__29211),
            .I(N__29203));
    Sp12to4 I__6049 (
            .O(N__29206),
            .I(N__29198));
    Sp12to4 I__6048 (
            .O(N__29203),
            .I(N__29198));
    Span12Mux_v I__6047 (
            .O(N__29198),
            .I(N__29195));
    Odrv12 I__6046 (
            .O(N__29195),
            .I(v33dsw_ok));
    CascadeMux I__6045 (
            .O(N__29192),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_ ));
    InMux I__6044 (
            .O(N__29189),
            .I(N__29185));
    InMux I__6043 (
            .O(N__29188),
            .I(N__29182));
    LocalMux I__6042 (
            .O(N__29185),
            .I(N__29179));
    LocalMux I__6041 (
            .O(N__29182),
            .I(N__29176));
    Span4Mux_h I__6040 (
            .O(N__29179),
            .I(N__29173));
    Odrv12 I__6039 (
            .O(N__29176),
            .I(\b2v_inst36.countZ0Z_9 ));
    Odrv4 I__6038 (
            .O(N__29173),
            .I(\b2v_inst36.countZ0Z_9 ));
    InMux I__6037 (
            .O(N__29168),
            .I(N__29162));
    InMux I__6036 (
            .O(N__29167),
            .I(N__29162));
    LocalMux I__6035 (
            .O(N__29162),
            .I(N__29159));
    Odrv4 I__6034 (
            .O(N__29159),
            .I(\b2v_inst36.count_rst_5 ));
    InMux I__6033 (
            .O(N__29156),
            .I(N__29153));
    LocalMux I__6032 (
            .O(N__29153),
            .I(\b2v_inst36.count_2_9 ));
    CascadeMux I__6031 (
            .O(N__29150),
            .I(N__29142));
    InMux I__6030 (
            .O(N__29149),
            .I(N__29136));
    CEMux I__6029 (
            .O(N__29148),
            .I(N__29136));
    InMux I__6028 (
            .O(N__29147),
            .I(N__29127));
    CEMux I__6027 (
            .O(N__29146),
            .I(N__29127));
    CEMux I__6026 (
            .O(N__29145),
            .I(N__29123));
    InMux I__6025 (
            .O(N__29142),
            .I(N__29111));
    CEMux I__6024 (
            .O(N__29141),
            .I(N__29111));
    LocalMux I__6023 (
            .O(N__29136),
            .I(N__29103));
    InMux I__6022 (
            .O(N__29135),
            .I(N__29098));
    InMux I__6021 (
            .O(N__29134),
            .I(N__29098));
    InMux I__6020 (
            .O(N__29133),
            .I(N__29088));
    CEMux I__6019 (
            .O(N__29132),
            .I(N__29088));
    LocalMux I__6018 (
            .O(N__29127),
            .I(N__29085));
    CEMux I__6017 (
            .O(N__29126),
            .I(N__29082));
    LocalMux I__6016 (
            .O(N__29123),
            .I(N__29079));
    InMux I__6015 (
            .O(N__29122),
            .I(N__29070));
    InMux I__6014 (
            .O(N__29121),
            .I(N__29070));
    InMux I__6013 (
            .O(N__29120),
            .I(N__29070));
    InMux I__6012 (
            .O(N__29119),
            .I(N__29070));
    InMux I__6011 (
            .O(N__29118),
            .I(N__29063));
    InMux I__6010 (
            .O(N__29117),
            .I(N__29063));
    InMux I__6009 (
            .O(N__29116),
            .I(N__29063));
    LocalMux I__6008 (
            .O(N__29111),
            .I(N__29060));
    InMux I__6007 (
            .O(N__29110),
            .I(N__29053));
    InMux I__6006 (
            .O(N__29109),
            .I(N__29053));
    InMux I__6005 (
            .O(N__29108),
            .I(N__29053));
    InMux I__6004 (
            .O(N__29107),
            .I(N__29048));
    InMux I__6003 (
            .O(N__29106),
            .I(N__29048));
    Span4Mux_h I__6002 (
            .O(N__29103),
            .I(N__29043));
    LocalMux I__6001 (
            .O(N__29098),
            .I(N__29043));
    InMux I__6000 (
            .O(N__29097),
            .I(N__29032));
    CEMux I__5999 (
            .O(N__29096),
            .I(N__29032));
    InMux I__5998 (
            .O(N__29095),
            .I(N__29032));
    InMux I__5997 (
            .O(N__29094),
            .I(N__29032));
    InMux I__5996 (
            .O(N__29093),
            .I(N__29032));
    LocalMux I__5995 (
            .O(N__29088),
            .I(N__29029));
    Span4Mux_h I__5994 (
            .O(N__29085),
            .I(N__29024));
    LocalMux I__5993 (
            .O(N__29082),
            .I(N__29024));
    Span4Mux_s3_v I__5992 (
            .O(N__29079),
            .I(N__29021));
    LocalMux I__5991 (
            .O(N__29070),
            .I(N__29016));
    LocalMux I__5990 (
            .O(N__29063),
            .I(N__29016));
    Span4Mux_s1_v I__5989 (
            .O(N__29060),
            .I(N__29005));
    LocalMux I__5988 (
            .O(N__29053),
            .I(N__29005));
    LocalMux I__5987 (
            .O(N__29048),
            .I(N__29005));
    Span4Mux_s1_v I__5986 (
            .O(N__29043),
            .I(N__29005));
    LocalMux I__5985 (
            .O(N__29032),
            .I(N__29005));
    Span4Mux_h I__5984 (
            .O(N__29029),
            .I(N__29002));
    Sp12to4 I__5983 (
            .O(N__29024),
            .I(N__28999));
    Span4Mux_v I__5982 (
            .O(N__29021),
            .I(N__28994));
    Span4Mux_s3_v I__5981 (
            .O(N__29016),
            .I(N__28994));
    Span4Mux_h I__5980 (
            .O(N__29005),
            .I(N__28991));
    Odrv4 I__5979 (
            .O(N__29002),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    Odrv12 I__5978 (
            .O(N__28999),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    Odrv4 I__5977 (
            .O(N__28994),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    Odrv4 I__5976 (
            .O(N__28991),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    SRMux I__5975 (
            .O(N__28982),
            .I(N__28977));
    SRMux I__5974 (
            .O(N__28981),
            .I(N__28969));
    SRMux I__5973 (
            .O(N__28980),
            .I(N__28966));
    LocalMux I__5972 (
            .O(N__28977),
            .I(N__28956));
    InMux I__5971 (
            .O(N__28976),
            .I(N__28951));
    InMux I__5970 (
            .O(N__28975),
            .I(N__28951));
    InMux I__5969 (
            .O(N__28974),
            .I(N__28946));
    InMux I__5968 (
            .O(N__28973),
            .I(N__28946));
    SRMux I__5967 (
            .O(N__28972),
            .I(N__28942));
    LocalMux I__5966 (
            .O(N__28969),
            .I(N__28931));
    LocalMux I__5965 (
            .O(N__28966),
            .I(N__28928));
    InMux I__5964 (
            .O(N__28965),
            .I(N__28921));
    InMux I__5963 (
            .O(N__28964),
            .I(N__28921));
    InMux I__5962 (
            .O(N__28963),
            .I(N__28921));
    SRMux I__5961 (
            .O(N__28962),
            .I(N__28911));
    InMux I__5960 (
            .O(N__28961),
            .I(N__28904));
    InMux I__5959 (
            .O(N__28960),
            .I(N__28904));
    SRMux I__5958 (
            .O(N__28959),
            .I(N__28904));
    Span4Mux_s2_v I__5957 (
            .O(N__28956),
            .I(N__28899));
    LocalMux I__5956 (
            .O(N__28951),
            .I(N__28899));
    LocalMux I__5955 (
            .O(N__28946),
            .I(N__28896));
    InMux I__5954 (
            .O(N__28945),
            .I(N__28893));
    LocalMux I__5953 (
            .O(N__28942),
            .I(N__28890));
    InMux I__5952 (
            .O(N__28941),
            .I(N__28883));
    InMux I__5951 (
            .O(N__28940),
            .I(N__28883));
    InMux I__5950 (
            .O(N__28939),
            .I(N__28883));
    SRMux I__5949 (
            .O(N__28938),
            .I(N__28878));
    InMux I__5948 (
            .O(N__28937),
            .I(N__28878));
    InMux I__5947 (
            .O(N__28936),
            .I(N__28871));
    InMux I__5946 (
            .O(N__28935),
            .I(N__28871));
    InMux I__5945 (
            .O(N__28934),
            .I(N__28871));
    Span4Mux_h I__5944 (
            .O(N__28931),
            .I(N__28866));
    Span4Mux_h I__5943 (
            .O(N__28928),
            .I(N__28866));
    LocalMux I__5942 (
            .O(N__28921),
            .I(N__28863));
    InMux I__5941 (
            .O(N__28920),
            .I(N__28856));
    InMux I__5940 (
            .O(N__28919),
            .I(N__28856));
    InMux I__5939 (
            .O(N__28918),
            .I(N__28856));
    InMux I__5938 (
            .O(N__28917),
            .I(N__28853));
    InMux I__5937 (
            .O(N__28916),
            .I(N__28850));
    InMux I__5936 (
            .O(N__28915),
            .I(N__28845));
    InMux I__5935 (
            .O(N__28914),
            .I(N__28845));
    LocalMux I__5934 (
            .O(N__28911),
            .I(N__28834));
    LocalMux I__5933 (
            .O(N__28904),
            .I(N__28834));
    Span4Mux_v I__5932 (
            .O(N__28899),
            .I(N__28834));
    Span4Mux_h I__5931 (
            .O(N__28896),
            .I(N__28834));
    LocalMux I__5930 (
            .O(N__28893),
            .I(N__28834));
    Span4Mux_v I__5929 (
            .O(N__28890),
            .I(N__28827));
    LocalMux I__5928 (
            .O(N__28883),
            .I(N__28827));
    LocalMux I__5927 (
            .O(N__28878),
            .I(N__28827));
    LocalMux I__5926 (
            .O(N__28871),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__5925 (
            .O(N__28866),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__5924 (
            .O(N__28863),
            .I(\b2v_inst36.count_0_sqmuxa ));
    LocalMux I__5923 (
            .O(N__28856),
            .I(\b2v_inst36.count_0_sqmuxa ));
    LocalMux I__5922 (
            .O(N__28853),
            .I(\b2v_inst36.count_0_sqmuxa ));
    LocalMux I__5921 (
            .O(N__28850),
            .I(\b2v_inst36.count_0_sqmuxa ));
    LocalMux I__5920 (
            .O(N__28845),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__5919 (
            .O(N__28834),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__5918 (
            .O(N__28827),
            .I(\b2v_inst36.count_0_sqmuxa ));
    InMux I__5917 (
            .O(N__28808),
            .I(N__28802));
    InMux I__5916 (
            .O(N__28807),
            .I(N__28802));
    LocalMux I__5915 (
            .O(N__28802),
            .I(N__28799));
    Odrv4 I__5914 (
            .O(N__28799),
            .I(\b2v_inst6.count_0_10 ));
    InMux I__5913 (
            .O(N__28796),
            .I(N__28791));
    InMux I__5912 (
            .O(N__28795),
            .I(N__28788));
    InMux I__5911 (
            .O(N__28794),
            .I(N__28785));
    LocalMux I__5910 (
            .O(N__28791),
            .I(N__28780));
    LocalMux I__5909 (
            .O(N__28788),
            .I(N__28780));
    LocalMux I__5908 (
            .O(N__28785),
            .I(\b2v_inst6.count_rst_4 ));
    Odrv4 I__5907 (
            .O(N__28780),
            .I(\b2v_inst6.count_rst_4 ));
    InMux I__5906 (
            .O(N__28775),
            .I(N__28772));
    LocalMux I__5905 (
            .O(N__28772),
            .I(N__28769));
    Odrv4 I__5904 (
            .O(N__28769),
            .I(\b2v_inst6.un2_count_1_axb_10 ));
    InMux I__5903 (
            .O(N__28766),
            .I(N__28763));
    LocalMux I__5902 (
            .O(N__28763),
            .I(N__28760));
    Sp12to4 I__5901 (
            .O(N__28760),
            .I(N__28757));
    Span12Mux_v I__5900 (
            .O(N__28757),
            .I(N__28754));
    Odrv12 I__5899 (
            .O(N__28754),
            .I(v33a_ok));
    InMux I__5898 (
            .O(N__28751),
            .I(N__28748));
    LocalMux I__5897 (
            .O(N__28748),
            .I(N__28745));
    Span4Mux_v I__5896 (
            .O(N__28745),
            .I(N__28742));
    Odrv4 I__5895 (
            .O(N__28742),
            .I(vccst_cpu_ok));
    CascadeMux I__5894 (
            .O(N__28739),
            .I(N__28736));
    InMux I__5893 (
            .O(N__28736),
            .I(N__28733));
    LocalMux I__5892 (
            .O(N__28733),
            .I(N__28730));
    Span4Mux_v I__5891 (
            .O(N__28730),
            .I(N__28727));
    Span4Mux_v I__5890 (
            .O(N__28727),
            .I(N__28724));
    Sp12to4 I__5889 (
            .O(N__28724),
            .I(N__28721));
    Odrv12 I__5888 (
            .O(N__28721),
            .I(v1p8a_ok));
    InMux I__5887 (
            .O(N__28718),
            .I(N__28715));
    LocalMux I__5886 (
            .O(N__28715),
            .I(N__28712));
    Odrv12 I__5885 (
            .O(N__28712),
            .I(v5a_ok));
    CascadeMux I__5884 (
            .O(N__28709),
            .I(\b2v_inst6.count_rst_5_cascade_ ));
    InMux I__5883 (
            .O(N__28706),
            .I(N__28703));
    LocalMux I__5882 (
            .O(N__28703),
            .I(\b2v_inst6.count_0_15 ));
    InMux I__5881 (
            .O(N__28700),
            .I(N__28694));
    InMux I__5880 (
            .O(N__28699),
            .I(N__28694));
    LocalMux I__5879 (
            .O(N__28694),
            .I(\b2v_inst6.count_rst ));
    InMux I__5878 (
            .O(N__28691),
            .I(N__28688));
    LocalMux I__5877 (
            .O(N__28688),
            .I(\b2v_inst6.countZ0Z_15 ));
    CascadeMux I__5876 (
            .O(N__28685),
            .I(\b2v_inst6.countZ0Z_15_cascade_ ));
    InMux I__5875 (
            .O(N__28682),
            .I(N__28678));
    InMux I__5874 (
            .O(N__28681),
            .I(N__28675));
    LocalMux I__5873 (
            .O(N__28678),
            .I(N__28672));
    LocalMux I__5872 (
            .O(N__28675),
            .I(\b2v_inst6.un2_count_1_axb_7 ));
    Odrv4 I__5871 (
            .O(N__28672),
            .I(\b2v_inst6.un2_count_1_axb_7 ));
    CascadeMux I__5870 (
            .O(N__28667),
            .I(N__28664));
    InMux I__5869 (
            .O(N__28664),
            .I(N__28658));
    InMux I__5868 (
            .O(N__28663),
            .I(N__28658));
    LocalMux I__5867 (
            .O(N__28658),
            .I(N__28655));
    Odrv12 I__5866 (
            .O(N__28655),
            .I(\b2v_inst6.un2_count_1_cry_6_THRU_CO ));
    CascadeMux I__5865 (
            .O(N__28652),
            .I(\b2v_inst6.un2_count_1_axb_7_cascade_ ));
    InMux I__5864 (
            .O(N__28649),
            .I(N__28646));
    LocalMux I__5863 (
            .O(N__28646),
            .I(\b2v_inst6.count_rst_7 ));
    InMux I__5862 (
            .O(N__28643),
            .I(N__28637));
    InMux I__5861 (
            .O(N__28642),
            .I(N__28637));
    LocalMux I__5860 (
            .O(N__28637),
            .I(\b2v_inst6.count_0_7 ));
    CascadeMux I__5859 (
            .O(N__28634),
            .I(\b2v_inst6.count_rst_7_cascade_ ));
    CascadeMux I__5858 (
            .O(N__28631),
            .I(\b2v_inst6.count_en_cascade_ ));
    InMux I__5857 (
            .O(N__28628),
            .I(N__28625));
    LocalMux I__5856 (
            .O(N__28625),
            .I(N__28622));
    Odrv4 I__5855 (
            .O(N__28622),
            .I(\b2v_inst6.countZ0Z_6 ));
    InMux I__5854 (
            .O(N__28619),
            .I(bfn_11_2_0_));
    InMux I__5853 (
            .O(N__28616),
            .I(\b2v_inst6.un2_count_1_cry_9 ));
    InMux I__5852 (
            .O(N__28613),
            .I(\b2v_inst6.un2_count_1_cry_10 ));
    InMux I__5851 (
            .O(N__28610),
            .I(\b2v_inst6.un2_count_1_cry_11 ));
    InMux I__5850 (
            .O(N__28607),
            .I(\b2v_inst6.un2_count_1_cry_12 ));
    InMux I__5849 (
            .O(N__28604),
            .I(\b2v_inst6.un2_count_1_cry_13 ));
    InMux I__5848 (
            .O(N__28601),
            .I(\b2v_inst6.un2_count_1_cry_14 ));
    InMux I__5847 (
            .O(N__28598),
            .I(N__28592));
    InMux I__5846 (
            .O(N__28597),
            .I(N__28592));
    LocalMux I__5845 (
            .O(N__28592),
            .I(\b2v_inst11.count_clk_1_13 ));
    InMux I__5844 (
            .O(N__28589),
            .I(N__28586));
    LocalMux I__5843 (
            .O(N__28586),
            .I(\b2v_inst11.count_clk_0_13 ));
    CEMux I__5842 (
            .O(N__28583),
            .I(N__28579));
    CascadeMux I__5841 (
            .O(N__28582),
            .I(N__28576));
    LocalMux I__5840 (
            .O(N__28579),
            .I(N__28573));
    InMux I__5839 (
            .O(N__28576),
            .I(N__28565));
    Span4Mux_s3_v I__5838 (
            .O(N__28573),
            .I(N__28562));
    CEMux I__5837 (
            .O(N__28572),
            .I(N__28559));
    InMux I__5836 (
            .O(N__28571),
            .I(N__28551));
    CEMux I__5835 (
            .O(N__28570),
            .I(N__28548));
    InMux I__5834 (
            .O(N__28569),
            .I(N__28543));
    CEMux I__5833 (
            .O(N__28568),
            .I(N__28543));
    LocalMux I__5832 (
            .O(N__28565),
            .I(N__28531));
    Span4Mux_h I__5831 (
            .O(N__28562),
            .I(N__28531));
    LocalMux I__5830 (
            .O(N__28559),
            .I(N__28531));
    InMux I__5829 (
            .O(N__28558),
            .I(N__28522));
    InMux I__5828 (
            .O(N__28557),
            .I(N__28522));
    InMux I__5827 (
            .O(N__28556),
            .I(N__28522));
    CEMux I__5826 (
            .O(N__28555),
            .I(N__28522));
    InMux I__5825 (
            .O(N__28554),
            .I(N__28519));
    LocalMux I__5824 (
            .O(N__28551),
            .I(N__28516));
    LocalMux I__5823 (
            .O(N__28548),
            .I(N__28513));
    LocalMux I__5822 (
            .O(N__28543),
            .I(N__28510));
    InMux I__5821 (
            .O(N__28542),
            .I(N__28501));
    CEMux I__5820 (
            .O(N__28541),
            .I(N__28501));
    InMux I__5819 (
            .O(N__28540),
            .I(N__28501));
    InMux I__5818 (
            .O(N__28539),
            .I(N__28501));
    CEMux I__5817 (
            .O(N__28538),
            .I(N__28498));
    IoSpan4Mux I__5816 (
            .O(N__28531),
            .I(N__28493));
    LocalMux I__5815 (
            .O(N__28522),
            .I(N__28493));
    LocalMux I__5814 (
            .O(N__28519),
            .I(N__28490));
    Span4Mux_s2_v I__5813 (
            .O(N__28516),
            .I(N__28480));
    Span4Mux_h I__5812 (
            .O(N__28513),
            .I(N__28480));
    Span4Mux_s1_v I__5811 (
            .O(N__28510),
            .I(N__28475));
    LocalMux I__5810 (
            .O(N__28501),
            .I(N__28475));
    LocalMux I__5809 (
            .O(N__28498),
            .I(N__28468));
    Span4Mux_s1_v I__5808 (
            .O(N__28493),
            .I(N__28468));
    Span4Mux_s1_v I__5807 (
            .O(N__28490),
            .I(N__28468));
    InMux I__5806 (
            .O(N__28489),
            .I(N__28465));
    InMux I__5805 (
            .O(N__28488),
            .I(N__28456));
    InMux I__5804 (
            .O(N__28487),
            .I(N__28456));
    InMux I__5803 (
            .O(N__28486),
            .I(N__28456));
    InMux I__5802 (
            .O(N__28485),
            .I(N__28456));
    Odrv4 I__5801 (
            .O(N__28480),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__5800 (
            .O(N__28475),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__5799 (
            .O(N__28468),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__5798 (
            .O(N__28465),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__5797 (
            .O(N__28456),
            .I(\b2v_inst11.count_clk_en ));
    InMux I__5796 (
            .O(N__28445),
            .I(\b2v_inst6.un2_count_1_cry_1 ));
    InMux I__5795 (
            .O(N__28442),
            .I(\b2v_inst6.un2_count_1_cry_2 ));
    InMux I__5794 (
            .O(N__28439),
            .I(\b2v_inst6.un2_count_1_cry_3 ));
    InMux I__5793 (
            .O(N__28436),
            .I(\b2v_inst6.un2_count_1_cry_4 ));
    InMux I__5792 (
            .O(N__28433),
            .I(\b2v_inst6.un2_count_1_cry_5 ));
    InMux I__5791 (
            .O(N__28430),
            .I(\b2v_inst6.un2_count_1_cry_6 ));
    InMux I__5790 (
            .O(N__28427),
            .I(\b2v_inst6.un2_count_1_cry_7 ));
    InMux I__5789 (
            .O(N__28424),
            .I(N__28419));
    InMux I__5788 (
            .O(N__28423),
            .I(N__28414));
    InMux I__5787 (
            .O(N__28422),
            .I(N__28414));
    LocalMux I__5786 (
            .O(N__28419),
            .I(N__28408));
    LocalMux I__5785 (
            .O(N__28414),
            .I(N__28408));
    InMux I__5784 (
            .O(N__28413),
            .I(N__28405));
    Span4Mux_h I__5783 (
            .O(N__28408),
            .I(N__28402));
    LocalMux I__5782 (
            .O(N__28405),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    Odrv4 I__5781 (
            .O(N__28402),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    CascadeMux I__5780 (
            .O(N__28397),
            .I(N__28394));
    InMux I__5779 (
            .O(N__28394),
            .I(N__28388));
    InMux I__5778 (
            .O(N__28393),
            .I(N__28388));
    LocalMux I__5777 (
            .O(N__28388),
            .I(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ));
    InMux I__5776 (
            .O(N__28385),
            .I(N__28382));
    LocalMux I__5775 (
            .O(N__28382),
            .I(\b2v_inst11.count_clk_0_7 ));
    InMux I__5774 (
            .O(N__28379),
            .I(N__28376));
    LocalMux I__5773 (
            .O(N__28376),
            .I(\b2v_inst11.count_clk_0_10 ));
    CascadeMux I__5772 (
            .O(N__28373),
            .I(N__28370));
    InMux I__5771 (
            .O(N__28370),
            .I(N__28366));
    InMux I__5770 (
            .O(N__28369),
            .I(N__28363));
    LocalMux I__5769 (
            .O(N__28366),
            .I(\b2v_inst11.count_clk_1_10 ));
    LocalMux I__5768 (
            .O(N__28363),
            .I(\b2v_inst11.count_clk_1_10 ));
    InMux I__5767 (
            .O(N__28358),
            .I(N__28355));
    LocalMux I__5766 (
            .O(N__28355),
            .I(\b2v_inst11.count_clkZ0Z_13 ));
    InMux I__5765 (
            .O(N__28352),
            .I(N__28348));
    InMux I__5764 (
            .O(N__28351),
            .I(N__28345));
    LocalMux I__5763 (
            .O(N__28348),
            .I(\b2v_inst11.count_clkZ0Z_11 ));
    LocalMux I__5762 (
            .O(N__28345),
            .I(\b2v_inst11.count_clkZ0Z_11 ));
    CascadeMux I__5761 (
            .O(N__28340),
            .I(\b2v_inst11.count_clkZ0Z_13_cascade_ ));
    InMux I__5760 (
            .O(N__28337),
            .I(N__28333));
    InMux I__5759 (
            .O(N__28336),
            .I(N__28330));
    LocalMux I__5758 (
            .O(N__28333),
            .I(\b2v_inst11.count_clkZ0Z_10 ));
    LocalMux I__5757 (
            .O(N__28330),
            .I(\b2v_inst11.count_clkZ0Z_10 ));
    InMux I__5756 (
            .O(N__28325),
            .I(N__28322));
    LocalMux I__5755 (
            .O(N__28322),
            .I(N__28319));
    Odrv4 I__5754 (
            .O(N__28319),
            .I(\b2v_inst11.un2_count_clk_17_0_o2_4 ));
    InMux I__5753 (
            .O(N__28316),
            .I(N__28312));
    InMux I__5752 (
            .O(N__28315),
            .I(N__28309));
    LocalMux I__5751 (
            .O(N__28312),
            .I(\b2v_inst11.count_clk_1_12 ));
    LocalMux I__5750 (
            .O(N__28309),
            .I(\b2v_inst11.count_clk_1_12 ));
    InMux I__5749 (
            .O(N__28304),
            .I(N__28301));
    LocalMux I__5748 (
            .O(N__28301),
            .I(\b2v_inst11.count_clk_0_12 ));
    InMux I__5747 (
            .O(N__28298),
            .I(N__28294));
    InMux I__5746 (
            .O(N__28297),
            .I(N__28291));
    LocalMux I__5745 (
            .O(N__28294),
            .I(\b2v_inst11.count_clkZ0Z_12 ));
    LocalMux I__5744 (
            .O(N__28291),
            .I(\b2v_inst11.count_clkZ0Z_12 ));
    InMux I__5743 (
            .O(N__28286),
            .I(N__28279));
    InMux I__5742 (
            .O(N__28285),
            .I(N__28279));
    InMux I__5741 (
            .O(N__28284),
            .I(N__28276));
    LocalMux I__5740 (
            .O(N__28279),
            .I(N__28273));
    LocalMux I__5739 (
            .O(N__28276),
            .I(\b2v_inst11.func_state_enZ0 ));
    Odrv4 I__5738 (
            .O(N__28273),
            .I(\b2v_inst11.func_state_enZ0 ));
    InMux I__5737 (
            .O(N__28268),
            .I(N__28265));
    LocalMux I__5736 (
            .O(N__28265),
            .I(\b2v_inst11.func_state_1_m2_1 ));
    CascadeMux I__5735 (
            .O(N__28262),
            .I(N__28259));
    InMux I__5734 (
            .O(N__28259),
            .I(N__28255));
    InMux I__5733 (
            .O(N__28258),
            .I(N__28252));
    LocalMux I__5732 (
            .O(N__28255),
            .I(\b2v_inst11.func_stateZ0Z_1 ));
    LocalMux I__5731 (
            .O(N__28252),
            .I(\b2v_inst11.func_stateZ0Z_1 ));
    InMux I__5730 (
            .O(N__28247),
            .I(N__28243));
    InMux I__5729 (
            .O(N__28246),
            .I(N__28240));
    LocalMux I__5728 (
            .O(N__28243),
            .I(N__28237));
    LocalMux I__5727 (
            .O(N__28240),
            .I(N__28234));
    Odrv4 I__5726 (
            .O(N__28237),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_5 ));
    Odrv4 I__5725 (
            .O(N__28234),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_5 ));
    InMux I__5724 (
            .O(N__28229),
            .I(N__28226));
    LocalMux I__5723 (
            .O(N__28226),
            .I(\b2v_inst11.func_state_1_m2s2_i_0 ));
    InMux I__5722 (
            .O(N__28223),
            .I(N__28220));
    LocalMux I__5721 (
            .O(N__28220),
            .I(N__28216));
    CascadeMux I__5720 (
            .O(N__28219),
            .I(N__28211));
    Span4Mux_v I__5719 (
            .O(N__28216),
            .I(N__28208));
    InMux I__5718 (
            .O(N__28215),
            .I(N__28205));
    InMux I__5717 (
            .O(N__28214),
            .I(N__28202));
    InMux I__5716 (
            .O(N__28211),
            .I(N__28199));
    Odrv4 I__5715 (
            .O(N__28208),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    LocalMux I__5714 (
            .O(N__28205),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    LocalMux I__5713 (
            .O(N__28202),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    LocalMux I__5712 (
            .O(N__28199),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    InMux I__5711 (
            .O(N__28190),
            .I(N__28187));
    LocalMux I__5710 (
            .O(N__28187),
            .I(N__28184));
    Span4Mux_s2_v I__5709 (
            .O(N__28184),
            .I(N__28181));
    Odrv4 I__5708 (
            .O(N__28181),
            .I(\b2v_inst11.count_clk_RNIZ0Z_0 ));
    InMux I__5707 (
            .O(N__28178),
            .I(N__28174));
    InMux I__5706 (
            .O(N__28177),
            .I(N__28170));
    LocalMux I__5705 (
            .O(N__28174),
            .I(N__28166));
    InMux I__5704 (
            .O(N__28173),
            .I(N__28163));
    LocalMux I__5703 (
            .O(N__28170),
            .I(N__28160));
    InMux I__5702 (
            .O(N__28169),
            .I(N__28157));
    Span12Mux_s7_h I__5701 (
            .O(N__28166),
            .I(N__28152));
    LocalMux I__5700 (
            .O(N__28163),
            .I(N__28149));
    Span4Mux_h I__5699 (
            .O(N__28160),
            .I(N__28144));
    LocalMux I__5698 (
            .O(N__28157),
            .I(N__28144));
    InMux I__5697 (
            .O(N__28156),
            .I(N__28139));
    InMux I__5696 (
            .O(N__28155),
            .I(N__28139));
    Odrv12 I__5695 (
            .O(N__28152),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    Odrv4 I__5694 (
            .O(N__28149),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    Odrv4 I__5693 (
            .O(N__28144),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    LocalMux I__5692 (
            .O(N__28139),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    InMux I__5691 (
            .O(N__28130),
            .I(N__28123));
    InMux I__5690 (
            .O(N__28129),
            .I(N__28114));
    InMux I__5689 (
            .O(N__28128),
            .I(N__28114));
    InMux I__5688 (
            .O(N__28127),
            .I(N__28114));
    InMux I__5687 (
            .O(N__28126),
            .I(N__28114));
    LocalMux I__5686 (
            .O(N__28123),
            .I(N__28111));
    LocalMux I__5685 (
            .O(N__28114),
            .I(N__28100));
    Span4Mux_v I__5684 (
            .O(N__28111),
            .I(N__28094));
    InMux I__5683 (
            .O(N__28110),
            .I(N__28091));
    InMux I__5682 (
            .O(N__28109),
            .I(N__28080));
    InMux I__5681 (
            .O(N__28108),
            .I(N__28080));
    InMux I__5680 (
            .O(N__28107),
            .I(N__28080));
    InMux I__5679 (
            .O(N__28106),
            .I(N__28080));
    InMux I__5678 (
            .O(N__28105),
            .I(N__28073));
    InMux I__5677 (
            .O(N__28104),
            .I(N__28073));
    InMux I__5676 (
            .O(N__28103),
            .I(N__28073));
    Span4Mux_s2_v I__5675 (
            .O(N__28100),
            .I(N__28070));
    InMux I__5674 (
            .O(N__28099),
            .I(N__28063));
    InMux I__5673 (
            .O(N__28098),
            .I(N__28063));
    InMux I__5672 (
            .O(N__28097),
            .I(N__28063));
    Span4Mux_v I__5671 (
            .O(N__28094),
            .I(N__28060));
    LocalMux I__5670 (
            .O(N__28091),
            .I(N__28057));
    InMux I__5669 (
            .O(N__28090),
            .I(N__28052));
    InMux I__5668 (
            .O(N__28089),
            .I(N__28052));
    LocalMux I__5667 (
            .O(N__28080),
            .I(N__28043));
    LocalMux I__5666 (
            .O(N__28073),
            .I(N__28043));
    Span4Mux_s3_h I__5665 (
            .O(N__28070),
            .I(N__28043));
    LocalMux I__5664 (
            .O(N__28063),
            .I(N__28043));
    Span4Mux_h I__5663 (
            .O(N__28060),
            .I(N__28040));
    Span4Mux_v I__5662 (
            .O(N__28057),
            .I(N__28037));
    LocalMux I__5661 (
            .O(N__28052),
            .I(N__28032));
    Span4Mux_s2_v I__5660 (
            .O(N__28043),
            .I(N__28032));
    Odrv4 I__5659 (
            .O(N__28040),
            .I(\b2v_inst11.func_state_RNINIV94_0_0 ));
    Odrv4 I__5658 (
            .O(N__28037),
            .I(\b2v_inst11.func_state_RNINIV94_0_0 ));
    Odrv4 I__5657 (
            .O(N__28032),
            .I(\b2v_inst11.func_state_RNINIV94_0_0 ));
    InMux I__5656 (
            .O(N__28025),
            .I(N__28022));
    LocalMux I__5655 (
            .O(N__28022),
            .I(\b2v_inst11.count_clk_0_0 ));
    CascadeMux I__5654 (
            .O(N__28019),
            .I(\b2v_inst11.func_state_1_m2_ns_1_0_cascade_ ));
    InMux I__5653 (
            .O(N__28016),
            .I(N__28010));
    InMux I__5652 (
            .O(N__28015),
            .I(N__28010));
    LocalMux I__5651 (
            .O(N__28010),
            .I(\b2v_inst11.func_state_1_m2_0 ));
    InMux I__5650 (
            .O(N__28007),
            .I(N__28004));
    LocalMux I__5649 (
            .O(N__28004),
            .I(\b2v_inst11.N_327 ));
    InMux I__5648 (
            .O(N__28001),
            .I(N__27998));
    LocalMux I__5647 (
            .O(N__27998),
            .I(N__27995));
    Odrv4 I__5646 (
            .O(N__27995),
            .I(\b2v_inst11.func_state_1_m2_ns_1_1_1 ));
    CascadeMux I__5645 (
            .O(N__27992),
            .I(\b2v_inst11.N_382_cascade_ ));
    InMux I__5644 (
            .O(N__27989),
            .I(N__27986));
    LocalMux I__5643 (
            .O(N__27986),
            .I(\b2v_inst11.un1_func_state25_6_0_2 ));
    CascadeMux I__5642 (
            .O(N__27983),
            .I(N__27979));
    CascadeMux I__5641 (
            .O(N__27982),
            .I(N__27976));
    InMux I__5640 (
            .O(N__27979),
            .I(N__27971));
    InMux I__5639 (
            .O(N__27976),
            .I(N__27968));
    CascadeMux I__5638 (
            .O(N__27975),
            .I(N__27965));
    CascadeMux I__5637 (
            .O(N__27974),
            .I(N__27962));
    LocalMux I__5636 (
            .O(N__27971),
            .I(N__27959));
    LocalMux I__5635 (
            .O(N__27968),
            .I(N__27956));
    InMux I__5634 (
            .O(N__27965),
            .I(N__27951));
    InMux I__5633 (
            .O(N__27962),
            .I(N__27951));
    Odrv4 I__5632 (
            .O(N__27959),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_0 ));
    Odrv4 I__5631 (
            .O(N__27956),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_0 ));
    LocalMux I__5630 (
            .O(N__27951),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_0 ));
    InMux I__5629 (
            .O(N__27944),
            .I(N__27941));
    LocalMux I__5628 (
            .O(N__27941),
            .I(N__27938));
    Span4Mux_v I__5627 (
            .O(N__27938),
            .I(N__27935));
    Odrv4 I__5626 (
            .O(N__27935),
            .I(\b2v_inst11.un1_func_state25_6_0_a3_1 ));
    InMux I__5625 (
            .O(N__27932),
            .I(N__27929));
    LocalMux I__5624 (
            .O(N__27929),
            .I(N__27924));
    InMux I__5623 (
            .O(N__27928),
            .I(N__27919));
    InMux I__5622 (
            .O(N__27927),
            .I(N__27919));
    Odrv4 I__5621 (
            .O(N__27924),
            .I(\b2v_inst11.N_406 ));
    LocalMux I__5620 (
            .O(N__27919),
            .I(\b2v_inst11.N_406 ));
    CascadeMux I__5619 (
            .O(N__27914),
            .I(N__27911));
    InMux I__5618 (
            .O(N__27911),
            .I(N__27908));
    LocalMux I__5617 (
            .O(N__27908),
            .I(\b2v_inst11.func_state_1_m2_ns_1_1 ));
    CascadeMux I__5616 (
            .O(N__27905),
            .I(\b2v_inst11.func_state_1_m2_1_cascade_ ));
    CascadeMux I__5615 (
            .O(N__27902),
            .I(\b2v_inst11.func_stateZ0Z_0_cascade_ ));
    InMux I__5614 (
            .O(N__27899),
            .I(N__27896));
    LocalMux I__5613 (
            .O(N__27896),
            .I(N__27893));
    Span4Mux_v I__5612 (
            .O(N__27893),
            .I(N__27890));
    Odrv4 I__5611 (
            .O(N__27890),
            .I(\b2v_inst11.N_337 ));
    CascadeMux I__5610 (
            .O(N__27887),
            .I(\b2v_inst11.N_338_cascade_ ));
    InMux I__5609 (
            .O(N__27884),
            .I(N__27880));
    InMux I__5608 (
            .O(N__27883),
            .I(N__27877));
    LocalMux I__5607 (
            .O(N__27880),
            .I(\b2v_inst11.N_76 ));
    LocalMux I__5606 (
            .O(N__27877),
            .I(\b2v_inst11.N_76 ));
    CascadeMux I__5605 (
            .O(N__27872),
            .I(\b2v_inst11.N_406_cascade_ ));
    InMux I__5604 (
            .O(N__27869),
            .I(N__27863));
    InMux I__5603 (
            .O(N__27868),
            .I(N__27863));
    LocalMux I__5602 (
            .O(N__27863),
            .I(\b2v_inst11.func_stateZ1Z_0 ));
    CascadeMux I__5601 (
            .O(N__27860),
            .I(\b2v_inst11.func_state_enZ0_cascade_ ));
    CascadeMux I__5600 (
            .O(N__27857),
            .I(\b2v_inst11.func_state_cascade_ ));
    CascadeMux I__5599 (
            .O(N__27854),
            .I(N__27851));
    InMux I__5598 (
            .O(N__27851),
            .I(N__27848));
    LocalMux I__5597 (
            .O(N__27848),
            .I(N__27845));
    Span4Mux_h I__5596 (
            .O(N__27845),
            .I(N__27841));
    InMux I__5595 (
            .O(N__27844),
            .I(N__27838));
    Odrv4 I__5594 (
            .O(N__27841),
            .I(\b2v_inst11.N_428 ));
    LocalMux I__5593 (
            .O(N__27838),
            .I(\b2v_inst11.N_428 ));
    CascadeMux I__5592 (
            .O(N__27833),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0_cascade_ ));
    InMux I__5591 (
            .O(N__27830),
            .I(N__27827));
    LocalMux I__5590 (
            .O(N__27827),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0 ));
    InMux I__5589 (
            .O(N__27824),
            .I(N__27818));
    InMux I__5588 (
            .O(N__27823),
            .I(N__27818));
    LocalMux I__5587 (
            .O(N__27818),
            .I(N__27815));
    Span4Mux_v I__5586 (
            .O(N__27815),
            .I(N__27812));
    Odrv4 I__5585 (
            .O(N__27812),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ));
    CascadeMux I__5584 (
            .O(N__27809),
            .I(N__27804));
    InMux I__5583 (
            .O(N__27808),
            .I(N__27798));
    InMux I__5582 (
            .O(N__27807),
            .I(N__27798));
    InMux I__5581 (
            .O(N__27804),
            .I(N__27793));
    InMux I__5580 (
            .O(N__27803),
            .I(N__27793));
    LocalMux I__5579 (
            .O(N__27798),
            .I(\b2v_inst11.N_369 ));
    LocalMux I__5578 (
            .O(N__27793),
            .I(\b2v_inst11.N_369 ));
    CascadeMux I__5577 (
            .O(N__27788),
            .I(\b2v_inst11.func_state_1_m2_ns_1_1_0_cascade_ ));
    CascadeMux I__5576 (
            .O(N__27785),
            .I(N__27782));
    InMux I__5575 (
            .O(N__27782),
            .I(N__27779));
    LocalMux I__5574 (
            .O(N__27779),
            .I(N__27776));
    Span4Mux_v I__5573 (
            .O(N__27776),
            .I(N__27773));
    Odrv4 I__5572 (
            .O(N__27773),
            .I(\b2v_inst11.g0_i_a7_1_2 ));
    InMux I__5571 (
            .O(N__27770),
            .I(N__27766));
    InMux I__5570 (
            .O(N__27769),
            .I(N__27763));
    LocalMux I__5569 (
            .O(N__27766),
            .I(N__27760));
    LocalMux I__5568 (
            .O(N__27763),
            .I(N__27756));
    Span4Mux_h I__5567 (
            .O(N__27760),
            .I(N__27753));
    InMux I__5566 (
            .O(N__27759),
            .I(N__27750));
    Span12Mux_s7_h I__5565 (
            .O(N__27756),
            .I(N__27747));
    Odrv4 I__5564 (
            .O(N__27753),
            .I(\b2v_inst16.curr_state_RNIUCAD1Z0Z_0 ));
    LocalMux I__5563 (
            .O(N__27750),
            .I(\b2v_inst16.curr_state_RNIUCAD1Z0Z_0 ));
    Odrv12 I__5562 (
            .O(N__27747),
            .I(\b2v_inst16.curr_state_RNIUCAD1Z0Z_0 ));
    InMux I__5561 (
            .O(N__27740),
            .I(N__27737));
    LocalMux I__5560 (
            .O(N__27737),
            .I(N__27731));
    InMux I__5559 (
            .O(N__27736),
            .I(N__27726));
    InMux I__5558 (
            .O(N__27735),
            .I(N__27726));
    CascadeMux I__5557 (
            .O(N__27734),
            .I(N__27723));
    Span4Mux_v I__5556 (
            .O(N__27731),
            .I(N__27717));
    LocalMux I__5555 (
            .O(N__27726),
            .I(N__27714));
    InMux I__5554 (
            .O(N__27723),
            .I(N__27709));
    InMux I__5553 (
            .O(N__27722),
            .I(N__27709));
    InMux I__5552 (
            .O(N__27721),
            .I(N__27704));
    InMux I__5551 (
            .O(N__27720),
            .I(N__27704));
    Span4Mux_h I__5550 (
            .O(N__27717),
            .I(N__27699));
    Span4Mux_v I__5549 (
            .O(N__27714),
            .I(N__27699));
    LocalMux I__5548 (
            .O(N__27709),
            .I(N__27694));
    LocalMux I__5547 (
            .O(N__27704),
            .I(N__27694));
    Odrv4 I__5546 (
            .O(N__27699),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    Odrv12 I__5545 (
            .O(N__27694),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    InMux I__5544 (
            .O(N__27689),
            .I(N__27683));
    InMux I__5543 (
            .O(N__27688),
            .I(N__27683));
    LocalMux I__5542 (
            .O(N__27683),
            .I(N__27680));
    Span4Mux_v I__5541 (
            .O(N__27680),
            .I(N__27677));
    Span4Mux_v I__5540 (
            .O(N__27677),
            .I(N__27674));
    Span4Mux_h I__5539 (
            .O(N__27674),
            .I(N__27671));
    Odrv4 I__5538 (
            .O(N__27671),
            .I(\b2v_inst16.N_268 ));
    InMux I__5537 (
            .O(N__27668),
            .I(N__27665));
    LocalMux I__5536 (
            .O(N__27665),
            .I(\b2v_inst11.N_395 ));
    InMux I__5535 (
            .O(N__27662),
            .I(N__27656));
    InMux I__5534 (
            .O(N__27661),
            .I(N__27656));
    LocalMux I__5533 (
            .O(N__27656),
            .I(\b2v_inst11.N_159 ));
    CascadeMux I__5532 (
            .O(N__27653),
            .I(\b2v_inst11.N_159_cascade_ ));
    InMux I__5531 (
            .O(N__27650),
            .I(N__27647));
    LocalMux I__5530 (
            .O(N__27647),
            .I(N__27640));
    InMux I__5529 (
            .O(N__27646),
            .I(N__27637));
    InMux I__5528 (
            .O(N__27645),
            .I(N__27633));
    InMux I__5527 (
            .O(N__27644),
            .I(N__27628));
    InMux I__5526 (
            .O(N__27643),
            .I(N__27628));
    Span4Mux_v I__5525 (
            .O(N__27640),
            .I(N__27623));
    LocalMux I__5524 (
            .O(N__27637),
            .I(N__27623));
    InMux I__5523 (
            .O(N__27636),
            .I(N__27618));
    LocalMux I__5522 (
            .O(N__27633),
            .I(N__27615));
    LocalMux I__5521 (
            .O(N__27628),
            .I(N__27612));
    Span4Mux_h I__5520 (
            .O(N__27623),
            .I(N__27609));
    InMux I__5519 (
            .O(N__27622),
            .I(N__27606));
    InMux I__5518 (
            .O(N__27621),
            .I(N__27603));
    LocalMux I__5517 (
            .O(N__27618),
            .I(\b2v_inst11.N_425 ));
    Odrv4 I__5516 (
            .O(N__27615),
            .I(\b2v_inst11.N_425 ));
    Odrv4 I__5515 (
            .O(N__27612),
            .I(\b2v_inst11.N_425 ));
    Odrv4 I__5514 (
            .O(N__27609),
            .I(\b2v_inst11.N_425 ));
    LocalMux I__5513 (
            .O(N__27606),
            .I(\b2v_inst11.N_425 ));
    LocalMux I__5512 (
            .O(N__27603),
            .I(\b2v_inst11.N_425 ));
    InMux I__5511 (
            .O(N__27590),
            .I(N__27587));
    LocalMux I__5510 (
            .O(N__27587),
            .I(\b2v_inst11.g2 ));
    InMux I__5509 (
            .O(N__27584),
            .I(N__27581));
    LocalMux I__5508 (
            .O(N__27581),
            .I(N__27576));
    InMux I__5507 (
            .O(N__27580),
            .I(N__27570));
    InMux I__5506 (
            .O(N__27579),
            .I(N__27567));
    Span4Mux_s3_h I__5505 (
            .O(N__27576),
            .I(N__27564));
    InMux I__5504 (
            .O(N__27575),
            .I(N__27561));
    InMux I__5503 (
            .O(N__27574),
            .I(N__27558));
    InMux I__5502 (
            .O(N__27573),
            .I(N__27555));
    LocalMux I__5501 (
            .O(N__27570),
            .I(N__27552));
    LocalMux I__5500 (
            .O(N__27567),
            .I(\b2v_inst11.N_366 ));
    Odrv4 I__5499 (
            .O(N__27564),
            .I(\b2v_inst11.N_366 ));
    LocalMux I__5498 (
            .O(N__27561),
            .I(\b2v_inst11.N_366 ));
    LocalMux I__5497 (
            .O(N__27558),
            .I(\b2v_inst11.N_366 ));
    LocalMux I__5496 (
            .O(N__27555),
            .I(\b2v_inst11.N_366 ));
    Odrv4 I__5495 (
            .O(N__27552),
            .I(\b2v_inst11.N_366 ));
    CascadeMux I__5494 (
            .O(N__27539),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_0_cascade_ ));
    CascadeMux I__5493 (
            .O(N__27536),
            .I(\b2v_inst11.N_168_cascade_ ));
    InMux I__5492 (
            .O(N__27533),
            .I(N__27529));
    InMux I__5491 (
            .O(N__27532),
            .I(N__27524));
    LocalMux I__5490 (
            .O(N__27529),
            .I(N__27521));
    InMux I__5489 (
            .O(N__27528),
            .I(N__27518));
    CascadeMux I__5488 (
            .O(N__27527),
            .I(N__27515));
    LocalMux I__5487 (
            .O(N__27524),
            .I(N__27509));
    Span4Mux_v I__5486 (
            .O(N__27521),
            .I(N__27506));
    LocalMux I__5485 (
            .O(N__27518),
            .I(N__27503));
    InMux I__5484 (
            .O(N__27515),
            .I(N__27500));
    CascadeMux I__5483 (
            .O(N__27514),
            .I(N__27496));
    InMux I__5482 (
            .O(N__27513),
            .I(N__27490));
    InMux I__5481 (
            .O(N__27512),
            .I(N__27490));
    Span4Mux_h I__5480 (
            .O(N__27509),
            .I(N__27487));
    Span4Mux_h I__5479 (
            .O(N__27506),
            .I(N__27480));
    Span4Mux_v I__5478 (
            .O(N__27503),
            .I(N__27480));
    LocalMux I__5477 (
            .O(N__27500),
            .I(N__27480));
    InMux I__5476 (
            .O(N__27499),
            .I(N__27473));
    InMux I__5475 (
            .O(N__27496),
            .I(N__27473));
    InMux I__5474 (
            .O(N__27495),
            .I(N__27473));
    LocalMux I__5473 (
            .O(N__27490),
            .I(curr_state_RNID8DP1_0_0));
    Odrv4 I__5472 (
            .O(N__27487),
            .I(curr_state_RNID8DP1_0_0));
    Odrv4 I__5471 (
            .O(N__27480),
            .I(curr_state_RNID8DP1_0_0));
    LocalMux I__5470 (
            .O(N__27473),
            .I(curr_state_RNID8DP1_0_0));
    InMux I__5469 (
            .O(N__27464),
            .I(N__27460));
    InMux I__5468 (
            .O(N__27463),
            .I(N__27455));
    LocalMux I__5467 (
            .O(N__27460),
            .I(N__27452));
    InMux I__5466 (
            .O(N__27459),
            .I(N__27449));
    InMux I__5465 (
            .O(N__27458),
            .I(N__27446));
    LocalMux I__5464 (
            .O(N__27455),
            .I(N__27442));
    Span4Mux_h I__5463 (
            .O(N__27452),
            .I(N__27437));
    LocalMux I__5462 (
            .O(N__27449),
            .I(N__27437));
    LocalMux I__5461 (
            .O(N__27446),
            .I(N__27434));
    CascadeMux I__5460 (
            .O(N__27445),
            .I(N__27429));
    Span4Mux_v I__5459 (
            .O(N__27442),
            .I(N__27424));
    Span4Mux_v I__5458 (
            .O(N__27437),
            .I(N__27424));
    Span12Mux_s3_h I__5457 (
            .O(N__27434),
            .I(N__27421));
    InMux I__5456 (
            .O(N__27433),
            .I(N__27414));
    InMux I__5455 (
            .O(N__27432),
            .I(N__27414));
    InMux I__5454 (
            .O(N__27429),
            .I(N__27414));
    Odrv4 I__5453 (
            .O(N__27424),
            .I(RSMRSTn_0));
    Odrv12 I__5452 (
            .O(N__27421),
            .I(RSMRSTn_0));
    LocalMux I__5451 (
            .O(N__27414),
            .I(RSMRSTn_0));
    CascadeMux I__5450 (
            .O(N__27407),
            .I(\b2v_inst11.count_clk_RNIDQ4A1Z0Z_6_cascade_ ));
    InMux I__5449 (
            .O(N__27404),
            .I(N__27401));
    LocalMux I__5448 (
            .O(N__27401),
            .I(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0 ));
    CascadeMux I__5447 (
            .O(N__27398),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_ ));
    CascadeMux I__5446 (
            .O(N__27395),
            .I(\b2v_inst11.N_186_i_cascade_ ));
    CascadeMux I__5445 (
            .O(N__27392),
            .I(\b2v_inst11.N_115_f0_cascade_ ));
    InMux I__5444 (
            .O(N__27389),
            .I(N__27386));
    LocalMux I__5443 (
            .O(N__27386),
            .I(\b2v_inst11.N_381 ));
    InMux I__5442 (
            .O(N__27383),
            .I(N__27374));
    InMux I__5441 (
            .O(N__27382),
            .I(N__27374));
    InMux I__5440 (
            .O(N__27381),
            .I(N__27374));
    LocalMux I__5439 (
            .O(N__27374),
            .I(N__27370));
    InMux I__5438 (
            .O(N__27373),
            .I(N__27367));
    Odrv4 I__5437 (
            .O(N__27370),
            .I(\b2v_inst5.curr_state_RNIZ0Z_1 ));
    LocalMux I__5436 (
            .O(N__27367),
            .I(\b2v_inst5.curr_state_RNIZ0Z_1 ));
    CascadeMux I__5435 (
            .O(N__27362),
            .I(N__27359));
    InMux I__5434 (
            .O(N__27359),
            .I(N__27352));
    InMux I__5433 (
            .O(N__27358),
            .I(N__27352));
    InMux I__5432 (
            .O(N__27357),
            .I(N__27349));
    LocalMux I__5431 (
            .O(N__27352),
            .I(\b2v_inst5.N_2898_i ));
    LocalMux I__5430 (
            .O(N__27349),
            .I(\b2v_inst5.N_2898_i ));
    InMux I__5429 (
            .O(N__27344),
            .I(N__27336));
    SRMux I__5428 (
            .O(N__27343),
            .I(N__27336));
    CascadeMux I__5427 (
            .O(N__27342),
            .I(N__27332));
    SRMux I__5426 (
            .O(N__27341),
            .I(N__27326));
    LocalMux I__5425 (
            .O(N__27336),
            .I(N__27320));
    InMux I__5424 (
            .O(N__27335),
            .I(N__27315));
    InMux I__5423 (
            .O(N__27332),
            .I(N__27315));
    SRMux I__5422 (
            .O(N__27331),
            .I(N__27310));
    InMux I__5421 (
            .O(N__27330),
            .I(N__27297));
    SRMux I__5420 (
            .O(N__27329),
            .I(N__27297));
    LocalMux I__5419 (
            .O(N__27326),
            .I(N__27294));
    CascadeMux I__5418 (
            .O(N__27325),
            .I(N__27290));
    InMux I__5417 (
            .O(N__27324),
            .I(N__27284));
    SRMux I__5416 (
            .O(N__27323),
            .I(N__27284));
    Span4Mux_h I__5415 (
            .O(N__27320),
            .I(N__27279));
    LocalMux I__5414 (
            .O(N__27315),
            .I(N__27279));
    InMux I__5413 (
            .O(N__27314),
            .I(N__27274));
    InMux I__5412 (
            .O(N__27313),
            .I(N__27274));
    LocalMux I__5411 (
            .O(N__27310),
            .I(N__27271));
    InMux I__5410 (
            .O(N__27309),
            .I(N__27262));
    InMux I__5409 (
            .O(N__27308),
            .I(N__27262));
    InMux I__5408 (
            .O(N__27307),
            .I(N__27262));
    InMux I__5407 (
            .O(N__27306),
            .I(N__27262));
    InMux I__5406 (
            .O(N__27305),
            .I(N__27257));
    InMux I__5405 (
            .O(N__27304),
            .I(N__27257));
    SRMux I__5404 (
            .O(N__27303),
            .I(N__27254));
    SRMux I__5403 (
            .O(N__27302),
            .I(N__27251));
    LocalMux I__5402 (
            .O(N__27297),
            .I(N__27248));
    Span4Mux_h I__5401 (
            .O(N__27294),
            .I(N__27245));
    InMux I__5400 (
            .O(N__27293),
            .I(N__27240));
    InMux I__5399 (
            .O(N__27290),
            .I(N__27240));
    CascadeMux I__5398 (
            .O(N__27289),
            .I(N__27237));
    LocalMux I__5397 (
            .O(N__27284),
            .I(N__27232));
    Span4Mux_s2_v I__5396 (
            .O(N__27279),
            .I(N__27232));
    LocalMux I__5395 (
            .O(N__27274),
            .I(N__27229));
    Span4Mux_v I__5394 (
            .O(N__27271),
            .I(N__27226));
    LocalMux I__5393 (
            .O(N__27262),
            .I(N__27221));
    LocalMux I__5392 (
            .O(N__27257),
            .I(N__27221));
    LocalMux I__5391 (
            .O(N__27254),
            .I(N__27210));
    LocalMux I__5390 (
            .O(N__27251),
            .I(N__27207));
    Span4Mux_v I__5389 (
            .O(N__27248),
            .I(N__27204));
    Span4Mux_v I__5388 (
            .O(N__27245),
            .I(N__27199));
    LocalMux I__5387 (
            .O(N__27240),
            .I(N__27199));
    InMux I__5386 (
            .O(N__27237),
            .I(N__27196));
    Span4Mux_v I__5385 (
            .O(N__27232),
            .I(N__27193));
    Span4Mux_h I__5384 (
            .O(N__27229),
            .I(N__27190));
    Span4Mux_v I__5383 (
            .O(N__27226),
            .I(N__27185));
    Span4Mux_h I__5382 (
            .O(N__27221),
            .I(N__27185));
    InMux I__5381 (
            .O(N__27220),
            .I(N__27174));
    InMux I__5380 (
            .O(N__27219),
            .I(N__27174));
    InMux I__5379 (
            .O(N__27218),
            .I(N__27174));
    InMux I__5378 (
            .O(N__27217),
            .I(N__27174));
    InMux I__5377 (
            .O(N__27216),
            .I(N__27174));
    InMux I__5376 (
            .O(N__27215),
            .I(N__27169));
    InMux I__5375 (
            .O(N__27214),
            .I(N__27169));
    InMux I__5374 (
            .O(N__27213),
            .I(N__27166));
    Odrv12 I__5373 (
            .O(N__27210),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv12 I__5372 (
            .O(N__27207),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__5371 (
            .O(N__27204),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__5370 (
            .O(N__27199),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__5369 (
            .O(N__27196),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__5368 (
            .O(N__27193),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__5367 (
            .O(N__27190),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__5366 (
            .O(N__27185),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__5365 (
            .O(N__27174),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__5364 (
            .O(N__27169),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__5363 (
            .O(N__27166),
            .I(\b2v_inst5.count_0_sqmuxa ));
    CascadeMux I__5362 (
            .O(N__27143),
            .I(N__27136));
    CascadeMux I__5361 (
            .O(N__27142),
            .I(N__27132));
    CascadeMux I__5360 (
            .O(N__27141),
            .I(N__27127));
    CascadeMux I__5359 (
            .O(N__27140),
            .I(N__27123));
    InMux I__5358 (
            .O(N__27139),
            .I(N__27111));
    InMux I__5357 (
            .O(N__27136),
            .I(N__27111));
    InMux I__5356 (
            .O(N__27135),
            .I(N__27111));
    InMux I__5355 (
            .O(N__27132),
            .I(N__27102));
    InMux I__5354 (
            .O(N__27131),
            .I(N__27102));
    InMux I__5353 (
            .O(N__27130),
            .I(N__27102));
    InMux I__5352 (
            .O(N__27127),
            .I(N__27102));
    InMux I__5351 (
            .O(N__27126),
            .I(N__27093));
    InMux I__5350 (
            .O(N__27123),
            .I(N__27093));
    InMux I__5349 (
            .O(N__27122),
            .I(N__27093));
    InMux I__5348 (
            .O(N__27121),
            .I(N__27093));
    InMux I__5347 (
            .O(N__27120),
            .I(N__27086));
    InMux I__5346 (
            .O(N__27119),
            .I(N__27086));
    InMux I__5345 (
            .O(N__27118),
            .I(N__27086));
    LocalMux I__5344 (
            .O(N__27111),
            .I(N__27081));
    LocalMux I__5343 (
            .O(N__27102),
            .I(N__27081));
    LocalMux I__5342 (
            .O(N__27093),
            .I(N__27074));
    LocalMux I__5341 (
            .O(N__27086),
            .I(N__27074));
    Span4Mux_v I__5340 (
            .O(N__27081),
            .I(N__27074));
    Odrv4 I__5339 (
            .O(N__27074),
            .I(\b2v_inst11.N_172_i ));
    CascadeMux I__5338 (
            .O(N__27071),
            .I(N__27068));
    InMux I__5337 (
            .O(N__27068),
            .I(N__27065));
    LocalMux I__5336 (
            .O(N__27065),
            .I(N__27062));
    Span4Mux_h I__5335 (
            .O(N__27062),
            .I(N__27059));
    Odrv4 I__5334 (
            .O(N__27059),
            .I(\b2v_inst11.un1_clk_100khz_2_i_o3_out ));
    CascadeMux I__5333 (
            .O(N__27056),
            .I(\b2v_inst11.N_19_cascade_ ));
    CascadeMux I__5332 (
            .O(N__27053),
            .I(rsmrstn_cascade_));
    CascadeMux I__5331 (
            .O(N__27050),
            .I(N__27047));
    InMux I__5330 (
            .O(N__27047),
            .I(N__27039));
    InMux I__5329 (
            .O(N__27046),
            .I(N__27039));
    InMux I__5328 (
            .O(N__27045),
            .I(N__27036));
    InMux I__5327 (
            .O(N__27044),
            .I(N__27033));
    LocalMux I__5326 (
            .O(N__27039),
            .I(N__27030));
    LocalMux I__5325 (
            .O(N__27036),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    LocalMux I__5324 (
            .O(N__27033),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    Odrv4 I__5323 (
            .O(N__27030),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    InMux I__5322 (
            .O(N__27023),
            .I(N__27020));
    LocalMux I__5321 (
            .O(N__27020),
            .I(N__27016));
    InMux I__5320 (
            .O(N__27019),
            .I(N__27012));
    Span4Mux_v I__5319 (
            .O(N__27016),
            .I(N__27009));
    InMux I__5318 (
            .O(N__27015),
            .I(N__27006));
    LocalMux I__5317 (
            .O(N__27012),
            .I(\b2v_inst5.countZ0Z_9 ));
    Odrv4 I__5316 (
            .O(N__27009),
            .I(\b2v_inst5.countZ0Z_9 ));
    LocalMux I__5315 (
            .O(N__27006),
            .I(\b2v_inst5.countZ0Z_9 ));
    InMux I__5314 (
            .O(N__26999),
            .I(N__26995));
    InMux I__5313 (
            .O(N__26998),
            .I(N__26992));
    LocalMux I__5312 (
            .O(N__26995),
            .I(N__26989));
    LocalMux I__5311 (
            .O(N__26992),
            .I(N__26984));
    Span4Mux_v I__5310 (
            .O(N__26989),
            .I(N__26984));
    Odrv4 I__5309 (
            .O(N__26984),
            .I(\b2v_inst5.un2_count_1_cry_8_THRU_CO ));
    CascadeMux I__5308 (
            .O(N__26981),
            .I(N__26976));
    CascadeMux I__5307 (
            .O(N__26980),
            .I(N__26970));
    InMux I__5306 (
            .O(N__26979),
            .I(N__26965));
    InMux I__5305 (
            .O(N__26976),
            .I(N__26965));
    InMux I__5304 (
            .O(N__26975),
            .I(N__26955));
    InMux I__5303 (
            .O(N__26974),
            .I(N__26955));
    InMux I__5302 (
            .O(N__26973),
            .I(N__26955));
    InMux I__5301 (
            .O(N__26970),
            .I(N__26952));
    LocalMux I__5300 (
            .O(N__26965),
            .I(N__26949));
    InMux I__5299 (
            .O(N__26964),
            .I(N__26942));
    InMux I__5298 (
            .O(N__26963),
            .I(N__26942));
    InMux I__5297 (
            .O(N__26962),
            .I(N__26942));
    LocalMux I__5296 (
            .O(N__26955),
            .I(N__26935));
    LocalMux I__5295 (
            .O(N__26952),
            .I(N__26928));
    Span4Mux_h I__5294 (
            .O(N__26949),
            .I(N__26928));
    LocalMux I__5293 (
            .O(N__26942),
            .I(N__26928));
    InMux I__5292 (
            .O(N__26941),
            .I(N__26921));
    InMux I__5291 (
            .O(N__26940),
            .I(N__26921));
    InMux I__5290 (
            .O(N__26939),
            .I(N__26921));
    InMux I__5289 (
            .O(N__26938),
            .I(N__26918));
    Odrv4 I__5288 (
            .O(N__26935),
            .I(\b2v_inst5.N_1_i ));
    Odrv4 I__5287 (
            .O(N__26928),
            .I(\b2v_inst5.N_1_i ));
    LocalMux I__5286 (
            .O(N__26921),
            .I(\b2v_inst5.N_1_i ));
    LocalMux I__5285 (
            .O(N__26918),
            .I(\b2v_inst5.N_1_i ));
    InMux I__5284 (
            .O(N__26909),
            .I(N__26906));
    LocalMux I__5283 (
            .O(N__26906),
            .I(\b2v_inst5.count_rst_5 ));
    InMux I__5282 (
            .O(N__26903),
            .I(N__26899));
    InMux I__5281 (
            .O(N__26902),
            .I(N__26896));
    LocalMux I__5280 (
            .O(N__26899),
            .I(N__26893));
    LocalMux I__5279 (
            .O(N__26896),
            .I(N__26890));
    Span4Mux_v I__5278 (
            .O(N__26893),
            .I(N__26885));
    Span4Mux_v I__5277 (
            .O(N__26890),
            .I(N__26885));
    Odrv4 I__5276 (
            .O(N__26885),
            .I(\b2v_inst5.count_rst_9 ));
    InMux I__5275 (
            .O(N__26882),
            .I(N__26879));
    LocalMux I__5274 (
            .O(N__26879),
            .I(N__26876));
    Odrv4 I__5273 (
            .O(N__26876),
            .I(\b2v_inst5.count_1_5 ));
    InMux I__5272 (
            .O(N__26873),
            .I(N__26869));
    CEMux I__5271 (
            .O(N__26872),
            .I(N__26866));
    LocalMux I__5270 (
            .O(N__26869),
            .I(N__26858));
    LocalMux I__5269 (
            .O(N__26866),
            .I(N__26858));
    CEMux I__5268 (
            .O(N__26865),
            .I(N__26852));
    InMux I__5267 (
            .O(N__26864),
            .I(N__26849));
    CEMux I__5266 (
            .O(N__26863),
            .I(N__26845));
    Span4Mux_h I__5265 (
            .O(N__26858),
            .I(N__26842));
    InMux I__5264 (
            .O(N__26857),
            .I(N__26835));
    InMux I__5263 (
            .O(N__26856),
            .I(N__26835));
    InMux I__5262 (
            .O(N__26855),
            .I(N__26835));
    LocalMux I__5261 (
            .O(N__26852),
            .I(N__26832));
    LocalMux I__5260 (
            .O(N__26849),
            .I(N__26829));
    CascadeMux I__5259 (
            .O(N__26848),
            .I(N__26822));
    LocalMux I__5258 (
            .O(N__26845),
            .I(N__26816));
    Span4Mux_s2_h I__5257 (
            .O(N__26842),
            .I(N__26808));
    LocalMux I__5256 (
            .O(N__26835),
            .I(N__26808));
    Span4Mux_v I__5255 (
            .O(N__26832),
            .I(N__26803));
    Span4Mux_v I__5254 (
            .O(N__26829),
            .I(N__26803));
    InMux I__5253 (
            .O(N__26828),
            .I(N__26787));
    InMux I__5252 (
            .O(N__26827),
            .I(N__26787));
    InMux I__5251 (
            .O(N__26826),
            .I(N__26787));
    InMux I__5250 (
            .O(N__26825),
            .I(N__26787));
    InMux I__5249 (
            .O(N__26822),
            .I(N__26782));
    CEMux I__5248 (
            .O(N__26821),
            .I(N__26782));
    CEMux I__5247 (
            .O(N__26820),
            .I(N__26779));
    CEMux I__5246 (
            .O(N__26819),
            .I(N__26776));
    Sp12to4 I__5245 (
            .O(N__26816),
            .I(N__26773));
    InMux I__5244 (
            .O(N__26815),
            .I(N__26766));
    InMux I__5243 (
            .O(N__26814),
            .I(N__26766));
    InMux I__5242 (
            .O(N__26813),
            .I(N__26766));
    Span4Mux_h I__5241 (
            .O(N__26808),
            .I(N__26763));
    Span4Mux_h I__5240 (
            .O(N__26803),
            .I(N__26760));
    InMux I__5239 (
            .O(N__26802),
            .I(N__26755));
    InMux I__5238 (
            .O(N__26801),
            .I(N__26755));
    CEMux I__5237 (
            .O(N__26800),
            .I(N__26744));
    InMux I__5236 (
            .O(N__26799),
            .I(N__26744));
    InMux I__5235 (
            .O(N__26798),
            .I(N__26744));
    InMux I__5234 (
            .O(N__26797),
            .I(N__26744));
    InMux I__5233 (
            .O(N__26796),
            .I(N__26744));
    LocalMux I__5232 (
            .O(N__26787),
            .I(N__26741));
    LocalMux I__5231 (
            .O(N__26782),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__5230 (
            .O(N__26779),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__5229 (
            .O(N__26776),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    Odrv12 I__5228 (
            .O(N__26773),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__5227 (
            .O(N__26766),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    Odrv4 I__5226 (
            .O(N__26763),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    Odrv4 I__5225 (
            .O(N__26760),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__5224 (
            .O(N__26755),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__5223 (
            .O(N__26744),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    Odrv4 I__5222 (
            .O(N__26741),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    CascadeMux I__5221 (
            .O(N__26720),
            .I(\b2v_inst5.curr_stateZ0Z_0_cascade_ ));
    InMux I__5220 (
            .O(N__26717),
            .I(N__26714));
    LocalMux I__5219 (
            .O(N__26714),
            .I(\b2v_inst5.m4_0 ));
    CascadeMux I__5218 (
            .O(N__26711),
            .I(\b2v_inst5.N_2898_i_cascade_ ));
    InMux I__5217 (
            .O(N__26708),
            .I(N__26699));
    InMux I__5216 (
            .O(N__26707),
            .I(N__26699));
    InMux I__5215 (
            .O(N__26706),
            .I(N__26699));
    LocalMux I__5214 (
            .O(N__26699),
            .I(N_413));
    InMux I__5213 (
            .O(N__26696),
            .I(N__26693));
    LocalMux I__5212 (
            .O(N__26693),
            .I(\b2v_inst5.curr_state_0_0 ));
    InMux I__5211 (
            .O(N__26690),
            .I(N__26681));
    InMux I__5210 (
            .O(N__26689),
            .I(N__26681));
    InMux I__5209 (
            .O(N__26688),
            .I(N__26681));
    LocalMux I__5208 (
            .O(N__26681),
            .I(\b2v_inst5.curr_stateZ0Z_0 ));
    CascadeMux I__5207 (
            .O(N__26678),
            .I(\b2v_inst5.countZ0Z_9_cascade_ ));
    CascadeMux I__5206 (
            .O(N__26675),
            .I(N__26672));
    InMux I__5205 (
            .O(N__26672),
            .I(N__26669));
    LocalMux I__5204 (
            .O(N__26669),
            .I(\b2v_inst5.count_1_9 ));
    InMux I__5203 (
            .O(N__26666),
            .I(N__26660));
    InMux I__5202 (
            .O(N__26665),
            .I(N__26660));
    LocalMux I__5201 (
            .O(N__26660),
            .I(N__26657));
    Span4Mux_h I__5200 (
            .O(N__26657),
            .I(N__26654));
    Odrv4 I__5199 (
            .O(N__26654),
            .I(\b2v_inst5.un2_count_1_cry_9_THRU_CO ));
    InMux I__5198 (
            .O(N__26651),
            .I(N__26648));
    LocalMux I__5197 (
            .O(N__26648),
            .I(N__26644));
    InMux I__5196 (
            .O(N__26647),
            .I(N__26641));
    Span4Mux_h I__5195 (
            .O(N__26644),
            .I(N__26638));
    LocalMux I__5194 (
            .O(N__26641),
            .I(\b2v_inst5.un2_count_1_axb_10 ));
    Odrv4 I__5193 (
            .O(N__26638),
            .I(\b2v_inst5.un2_count_1_axb_10 ));
    InMux I__5192 (
            .O(N__26633),
            .I(N__26627));
    InMux I__5191 (
            .O(N__26632),
            .I(N__26627));
    LocalMux I__5190 (
            .O(N__26627),
            .I(\b2v_inst5.count_rst_4 ));
    CascadeMux I__5189 (
            .O(N__26624),
            .I(\b2v_inst5.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__5188 (
            .O(N__26621),
            .I(\b2v_inst5.curr_state_RNIZ0Z_1_cascade_ ));
    CascadeMux I__5187 (
            .O(N__26618),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_ ));
    InMux I__5186 (
            .O(N__26615),
            .I(N__26611));
    InMux I__5185 (
            .O(N__26614),
            .I(N__26608));
    LocalMux I__5184 (
            .O(N__26611),
            .I(N__26605));
    LocalMux I__5183 (
            .O(N__26608),
            .I(\b2v_inst5.countZ0Z_15 ));
    Odrv12 I__5182 (
            .O(N__26605),
            .I(\b2v_inst5.countZ0Z_15 ));
    InMux I__5181 (
            .O(N__26600),
            .I(N__26594));
    InMux I__5180 (
            .O(N__26599),
            .I(N__26594));
    LocalMux I__5179 (
            .O(N__26594),
            .I(N__26591));
    Odrv4 I__5178 (
            .O(N__26591),
            .I(\b2v_inst5.count_rst ));
    InMux I__5177 (
            .O(N__26588),
            .I(N__26585));
    LocalMux I__5176 (
            .O(N__26585),
            .I(\b2v_inst5.count_1_15 ));
    InMux I__5175 (
            .O(N__26582),
            .I(N__26579));
    LocalMux I__5174 (
            .O(N__26579),
            .I(\b2v_inst5.curr_stateZ0Z_1 ));
    InMux I__5173 (
            .O(N__26576),
            .I(N__26570));
    InMux I__5172 (
            .O(N__26575),
            .I(N__26570));
    LocalMux I__5171 (
            .O(N__26570),
            .I(N__26567));
    Span4Mux_h I__5170 (
            .O(N__26567),
            .I(N__26564));
    Odrv4 I__5169 (
            .O(N__26564),
            .I(\b2v_inst5.count_rst_11 ));
    InMux I__5168 (
            .O(N__26561),
            .I(N__26558));
    LocalMux I__5167 (
            .O(N__26558),
            .I(\b2v_inst5.count_1_3 ));
    CascadeMux I__5166 (
            .O(N__26555),
            .I(N__26552));
    InMux I__5165 (
            .O(N__26552),
            .I(N__26549));
    LocalMux I__5164 (
            .O(N__26549),
            .I(N__26546));
    Span4Mux_v I__5163 (
            .O(N__26546),
            .I(N__26543));
    Odrv4 I__5162 (
            .O(N__26543),
            .I(\b2v_inst5.countZ0Z_3 ));
    InMux I__5161 (
            .O(N__26540),
            .I(N__26537));
    LocalMux I__5160 (
            .O(N__26537),
            .I(N__26532));
    InMux I__5159 (
            .O(N__26536),
            .I(N__26529));
    InMux I__5158 (
            .O(N__26535),
            .I(N__26526));
    Odrv4 I__5157 (
            .O(N__26532),
            .I(\b2v_inst5.countZ0Z_13 ));
    LocalMux I__5156 (
            .O(N__26529),
            .I(\b2v_inst5.countZ0Z_13 ));
    LocalMux I__5155 (
            .O(N__26526),
            .I(\b2v_inst5.countZ0Z_13 ));
    InMux I__5154 (
            .O(N__26519),
            .I(N__26516));
    LocalMux I__5153 (
            .O(N__26516),
            .I(N__26512));
    InMux I__5152 (
            .O(N__26515),
            .I(N__26509));
    Span4Mux_h I__5151 (
            .O(N__26512),
            .I(N__26506));
    LocalMux I__5150 (
            .O(N__26509),
            .I(\b2v_inst5.countZ0Z_1 ));
    Odrv4 I__5149 (
            .O(N__26506),
            .I(\b2v_inst5.countZ0Z_1 ));
    CascadeMux I__5148 (
            .O(N__26501),
            .I(\b2v_inst5.countZ0Z_3_cascade_ ));
    InMux I__5147 (
            .O(N__26498),
            .I(N__26495));
    LocalMux I__5146 (
            .O(N__26495),
            .I(N__26491));
    InMux I__5145 (
            .O(N__26494),
            .I(N__26488));
    Span4Mux_h I__5144 (
            .O(N__26491),
            .I(N__26485));
    LocalMux I__5143 (
            .O(N__26488),
            .I(\b2v_inst5.countZ0Z_2 ));
    Odrv4 I__5142 (
            .O(N__26485),
            .I(\b2v_inst5.countZ0Z_2 ));
    InMux I__5141 (
            .O(N__26480),
            .I(N__26477));
    LocalMux I__5140 (
            .O(N__26477),
            .I(N__26474));
    Odrv4 I__5139 (
            .O(N__26474),
            .I(\b2v_inst5.un12_clk_100khz_11 ));
    InMux I__5138 (
            .O(N__26471),
            .I(N__26468));
    LocalMux I__5137 (
            .O(N__26468),
            .I(N__26465));
    Odrv4 I__5136 (
            .O(N__26465),
            .I(\b2v_inst5.un12_clk_100khz_4 ));
    CascadeMux I__5135 (
            .O(N__26462),
            .I(\b2v_inst5.un12_clk_100khz_5_cascade_ ));
    CascadeMux I__5134 (
            .O(N__26459),
            .I(\b2v_inst5.un2_count_1_axb_10_cascade_ ));
    CascadeMux I__5133 (
            .O(N__26456),
            .I(N__26452));
    CascadeMux I__5132 (
            .O(N__26455),
            .I(N__26449));
    InMux I__5131 (
            .O(N__26452),
            .I(N__26444));
    InMux I__5130 (
            .O(N__26449),
            .I(N__26444));
    LocalMux I__5129 (
            .O(N__26444),
            .I(\b2v_inst5.count_1_10 ));
    InMux I__5128 (
            .O(N__26441),
            .I(N__26438));
    LocalMux I__5127 (
            .O(N__26438),
            .I(N__26435));
    Span4Mux_v I__5126 (
            .O(N__26435),
            .I(N__26432));
    Odrv4 I__5125 (
            .O(N__26432),
            .I(\b2v_inst5.un12_clk_100khz_1 ));
    InMux I__5124 (
            .O(N__26429),
            .I(N__26426));
    LocalMux I__5123 (
            .O(N__26426),
            .I(N__26422));
    InMux I__5122 (
            .O(N__26425),
            .I(N__26419));
    Span4Mux_h I__5121 (
            .O(N__26422),
            .I(N__26416));
    LocalMux I__5120 (
            .O(N__26419),
            .I(\b2v_inst5.countZ0Z_5 ));
    Odrv4 I__5119 (
            .O(N__26416),
            .I(\b2v_inst5.countZ0Z_5 ));
    CascadeMux I__5118 (
            .O(N__26411),
            .I(N__26408));
    InMux I__5117 (
            .O(N__26408),
            .I(N__26405));
    LocalMux I__5116 (
            .O(N__26405),
            .I(\b2v_inst5.un12_clk_100khz_9 ));
    InMux I__5115 (
            .O(N__26402),
            .I(N__26399));
    LocalMux I__5114 (
            .O(N__26399),
            .I(N__26395));
    InMux I__5113 (
            .O(N__26398),
            .I(N__26392));
    Span4Mux_v I__5112 (
            .O(N__26395),
            .I(N__26389));
    LocalMux I__5111 (
            .O(N__26392),
            .I(N__26386));
    Span4Mux_v I__5110 (
            .O(N__26389),
            .I(N__26383));
    Span4Mux_v I__5109 (
            .O(N__26386),
            .I(N__26380));
    Odrv4 I__5108 (
            .O(N__26383),
            .I(\b2v_inst5.countZ0Z_6 ));
    Odrv4 I__5107 (
            .O(N__26380),
            .I(\b2v_inst5.countZ0Z_6 ));
    InMux I__5106 (
            .O(N__26375),
            .I(N__26372));
    LocalMux I__5105 (
            .O(N__26372),
            .I(\b2v_inst5.un12_clk_100khz_12 ));
    InMux I__5104 (
            .O(N__26369),
            .I(N__26364));
    InMux I__5103 (
            .O(N__26368),
            .I(N__26359));
    InMux I__5102 (
            .O(N__26367),
            .I(N__26359));
    LocalMux I__5101 (
            .O(N__26364),
            .I(\b2v_inst36.count_rst_8 ));
    LocalMux I__5100 (
            .O(N__26359),
            .I(\b2v_inst36.count_rst_8 ));
    CascadeMux I__5099 (
            .O(N__26354),
            .I(\b2v_inst36.countZ0Z_4_cascade_ ));
    InMux I__5098 (
            .O(N__26351),
            .I(N__26345));
    InMux I__5097 (
            .O(N__26350),
            .I(N__26345));
    LocalMux I__5096 (
            .O(N__26345),
            .I(\b2v_inst36.count_2_6 ));
    InMux I__5095 (
            .O(N__26342),
            .I(N__26339));
    LocalMux I__5094 (
            .O(N__26339),
            .I(\b2v_inst36.un12_clk_100khz_0 ));
    InMux I__5093 (
            .O(N__26336),
            .I(N__26333));
    LocalMux I__5092 (
            .O(N__26333),
            .I(\b2v_inst36.un2_count_1_axb_12 ));
    InMux I__5091 (
            .O(N__26330),
            .I(N__26324));
    InMux I__5090 (
            .O(N__26329),
            .I(N__26324));
    LocalMux I__5089 (
            .O(N__26324),
            .I(\b2v_inst36.count_2_12 ));
    CascadeMux I__5088 (
            .O(N__26321),
            .I(N__26318));
    InMux I__5087 (
            .O(N__26318),
            .I(N__26313));
    InMux I__5086 (
            .O(N__26317),
            .I(N__26308));
    InMux I__5085 (
            .O(N__26316),
            .I(N__26308));
    LocalMux I__5084 (
            .O(N__26313),
            .I(\b2v_inst36.count_rst_2 ));
    LocalMux I__5083 (
            .O(N__26308),
            .I(\b2v_inst36.count_rst_2 ));
    InMux I__5082 (
            .O(N__26303),
            .I(N__26300));
    LocalMux I__5081 (
            .O(N__26300),
            .I(\b2v_inst36.un12_clk_100khz_1 ));
    InMux I__5080 (
            .O(N__26297),
            .I(N__26291));
    InMux I__5079 (
            .O(N__26296),
            .I(N__26291));
    LocalMux I__5078 (
            .O(N__26291),
            .I(N__26288));
    Span4Mux_v I__5077 (
            .O(N__26288),
            .I(N__26285));
    Odrv4 I__5076 (
            .O(N__26285),
            .I(\b2v_inst5.count_rst_13 ));
    InMux I__5075 (
            .O(N__26282),
            .I(N__26279));
    LocalMux I__5074 (
            .O(N__26279),
            .I(\b2v_inst5.count_1_1 ));
    InMux I__5073 (
            .O(N__26276),
            .I(N__26270));
    InMux I__5072 (
            .O(N__26275),
            .I(N__26270));
    LocalMux I__5071 (
            .O(N__26270),
            .I(N__26267));
    Span4Mux_h I__5070 (
            .O(N__26267),
            .I(N__26264));
    Odrv4 I__5069 (
            .O(N__26264),
            .I(\b2v_inst5.count_rst_12 ));
    InMux I__5068 (
            .O(N__26261),
            .I(N__26258));
    LocalMux I__5067 (
            .O(N__26258),
            .I(\b2v_inst5.count_1_2 ));
    InMux I__5066 (
            .O(N__26255),
            .I(N__26252));
    LocalMux I__5065 (
            .O(N__26252),
            .I(\b2v_inst36.un12_clk_100khz_5 ));
    InMux I__5064 (
            .O(N__26249),
            .I(N__26246));
    LocalMux I__5063 (
            .O(N__26246),
            .I(\b2v_inst36.un12_clk_100khz_4 ));
    CascadeMux I__5062 (
            .O(N__26243),
            .I(\b2v_inst36.un12_clk_100khz_6_cascade_ ));
    InMux I__5061 (
            .O(N__26240),
            .I(N__26237));
    LocalMux I__5060 (
            .O(N__26237),
            .I(N__26234));
    Span4Mux_v I__5059 (
            .O(N__26234),
            .I(N__26231));
    Odrv4 I__5058 (
            .O(N__26231),
            .I(\b2v_inst36.un12_clk_100khz_7 ));
    InMux I__5057 (
            .O(N__26228),
            .I(N__26225));
    LocalMux I__5056 (
            .O(N__26225),
            .I(N__26222));
    Odrv12 I__5055 (
            .O(N__26222),
            .I(\b2v_inst36.un12_clk_100khz_9 ));
    CascadeMux I__5054 (
            .O(N__26219),
            .I(\b2v_inst36.un12_clk_100khz_13_cascade_ ));
    CascadeMux I__5053 (
            .O(N__26216),
            .I(\b2v_inst36.N_1_i_cascade_ ));
    InMux I__5052 (
            .O(N__26213),
            .I(N__26210));
    LocalMux I__5051 (
            .O(N__26210),
            .I(\b2v_inst36.count_rst_4 ));
    CascadeMux I__5050 (
            .O(N__26207),
            .I(\b2v_inst36.count_rst_4_cascade_ ));
    InMux I__5049 (
            .O(N__26204),
            .I(N__26201));
    LocalMux I__5048 (
            .O(N__26201),
            .I(N__26197));
    InMux I__5047 (
            .O(N__26200),
            .I(N__26194));
    Odrv4 I__5046 (
            .O(N__26197),
            .I(\b2v_inst36.un2_count_1_axb_10 ));
    LocalMux I__5045 (
            .O(N__26194),
            .I(\b2v_inst36.un2_count_1_axb_10 ));
    InMux I__5044 (
            .O(N__26189),
            .I(N__26183));
    InMux I__5043 (
            .O(N__26188),
            .I(N__26183));
    LocalMux I__5042 (
            .O(N__26183),
            .I(N__26180));
    Odrv4 I__5041 (
            .O(N__26180),
            .I(\b2v_inst36.un2_count_1_cry_9_THRU_CO ));
    CascadeMux I__5040 (
            .O(N__26177),
            .I(\b2v_inst36.un2_count_1_axb_10_cascade_ ));
    CascadeMux I__5039 (
            .O(N__26174),
            .I(N__26166));
    InMux I__5038 (
            .O(N__26173),
            .I(N__26163));
    InMux I__5037 (
            .O(N__26172),
            .I(N__26156));
    InMux I__5036 (
            .O(N__26171),
            .I(N__26156));
    InMux I__5035 (
            .O(N__26170),
            .I(N__26156));
    CascadeMux I__5034 (
            .O(N__26169),
            .I(N__26149));
    InMux I__5033 (
            .O(N__26166),
            .I(N__26139));
    LocalMux I__5032 (
            .O(N__26163),
            .I(N__26134));
    LocalMux I__5031 (
            .O(N__26156),
            .I(N__26134));
    InMux I__5030 (
            .O(N__26155),
            .I(N__26127));
    InMux I__5029 (
            .O(N__26154),
            .I(N__26127));
    InMux I__5028 (
            .O(N__26153),
            .I(N__26124));
    InMux I__5027 (
            .O(N__26152),
            .I(N__26119));
    InMux I__5026 (
            .O(N__26149),
            .I(N__26119));
    InMux I__5025 (
            .O(N__26148),
            .I(N__26112));
    InMux I__5024 (
            .O(N__26147),
            .I(N__26112));
    InMux I__5023 (
            .O(N__26146),
            .I(N__26112));
    InMux I__5022 (
            .O(N__26145),
            .I(N__26103));
    InMux I__5021 (
            .O(N__26144),
            .I(N__26103));
    InMux I__5020 (
            .O(N__26143),
            .I(N__26103));
    InMux I__5019 (
            .O(N__26142),
            .I(N__26103));
    LocalMux I__5018 (
            .O(N__26139),
            .I(N__26100));
    Span4Mux_s1_v I__5017 (
            .O(N__26134),
            .I(N__26097));
    InMux I__5016 (
            .O(N__26133),
            .I(N__26092));
    InMux I__5015 (
            .O(N__26132),
            .I(N__26092));
    LocalMux I__5014 (
            .O(N__26127),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__5013 (
            .O(N__26124),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__5012 (
            .O(N__26119),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__5011 (
            .O(N__26112),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__5010 (
            .O(N__26103),
            .I(\b2v_inst36.N_1_i ));
    Odrv4 I__5009 (
            .O(N__26100),
            .I(\b2v_inst36.N_1_i ));
    Odrv4 I__5008 (
            .O(N__26097),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__5007 (
            .O(N__26092),
            .I(\b2v_inst36.N_1_i ));
    InMux I__5006 (
            .O(N__26075),
            .I(N__26069));
    InMux I__5005 (
            .O(N__26074),
            .I(N__26069));
    LocalMux I__5004 (
            .O(N__26069),
            .I(\b2v_inst36.count_2_10 ));
    InMux I__5003 (
            .O(N__26066),
            .I(N__26063));
    LocalMux I__5002 (
            .O(N__26063),
            .I(\b2v_inst36.un2_count_1_axb_6 ));
    InMux I__5001 (
            .O(N__26060),
            .I(N__26054));
    InMux I__5000 (
            .O(N__26059),
            .I(N__26054));
    LocalMux I__4999 (
            .O(N__26054),
            .I(\b2v_inst36.count_rst_10 ));
    InMux I__4998 (
            .O(N__26051),
            .I(N__26048));
    LocalMux I__4997 (
            .O(N__26048),
            .I(\b2v_inst36.count_2_4 ));
    InMux I__4996 (
            .O(N__26045),
            .I(N__26042));
    LocalMux I__4995 (
            .O(N__26042),
            .I(\b2v_inst36.countZ0Z_4 ));
    CascadeMux I__4994 (
            .O(N__26039),
            .I(\b2v_inst36.curr_stateZ0Z_0_cascade_ ));
    InMux I__4993 (
            .O(N__26036),
            .I(N__26033));
    LocalMux I__4992 (
            .O(N__26033),
            .I(\b2v_inst36.curr_state_0_0 ));
    InMux I__4991 (
            .O(N__26030),
            .I(N__26027));
    LocalMux I__4990 (
            .O(N__26027),
            .I(\b2v_inst36.curr_state_0_1 ));
    InMux I__4989 (
            .O(N__26024),
            .I(N__26021));
    LocalMux I__4988 (
            .O(N__26021),
            .I(\b2v_inst36.curr_state_7_1 ));
    CascadeMux I__4987 (
            .O(N__26018),
            .I(\b2v_inst36.curr_stateZ0Z_1_cascade_ ));
    InMux I__4986 (
            .O(N__26015),
            .I(N__26012));
    LocalMux I__4985 (
            .O(N__26012),
            .I(N__26009));
    Span4Mux_v I__4984 (
            .O(N__26009),
            .I(N__26006));
    Odrv4 I__4983 (
            .O(N__26006),
            .I(\b2v_inst36.DSW_PWROK_0 ));
    CascadeMux I__4982 (
            .O(N__26003),
            .I(N__26000));
    InMux I__4981 (
            .O(N__26000),
            .I(N__25996));
    InMux I__4980 (
            .O(N__25999),
            .I(N__25993));
    LocalMux I__4979 (
            .O(N__25996),
            .I(N__25990));
    LocalMux I__4978 (
            .O(N__25993),
            .I(N__25987));
    Odrv4 I__4977 (
            .O(N__25990),
            .I(\b2v_inst36.un2_count_1_cry_7_THRU_CO ));
    Odrv4 I__4976 (
            .O(N__25987),
            .I(\b2v_inst36.un2_count_1_cry_7_THRU_CO ));
    InMux I__4975 (
            .O(N__25982),
            .I(N__25979));
    LocalMux I__4974 (
            .O(N__25979),
            .I(\b2v_inst36.count_2_8 ));
    InMux I__4973 (
            .O(N__25976),
            .I(N__25973));
    LocalMux I__4972 (
            .O(N__25973),
            .I(\b2v_inst36.count_rst_6 ));
    CascadeMux I__4971 (
            .O(N__25970),
            .I(N__25966));
    CascadeMux I__4970 (
            .O(N__25969),
            .I(N__25963));
    InMux I__4969 (
            .O(N__25966),
            .I(N__25959));
    InMux I__4968 (
            .O(N__25963),
            .I(N__25956));
    InMux I__4967 (
            .O(N__25962),
            .I(N__25953));
    LocalMux I__4966 (
            .O(N__25959),
            .I(N__25948));
    LocalMux I__4965 (
            .O(N__25956),
            .I(N__25948));
    LocalMux I__4964 (
            .O(N__25953),
            .I(\b2v_inst36.countZ0Z_8 ));
    Odrv4 I__4963 (
            .O(N__25948),
            .I(\b2v_inst36.countZ0Z_8 ));
    CascadeMux I__4962 (
            .O(N__25943),
            .I(\b2v_inst36.countZ0Z_8_cascade_ ));
    InMux I__4961 (
            .O(N__25940),
            .I(\b2v_inst11.un1_count_clk_2_cry_10 ));
    InMux I__4960 (
            .O(N__25937),
            .I(\b2v_inst11.un1_count_clk_2_cry_11 ));
    InMux I__4959 (
            .O(N__25934),
            .I(\b2v_inst11.un1_count_clk_2_cry_12 ));
    InMux I__4958 (
            .O(N__25931),
            .I(N__25927));
    InMux I__4957 (
            .O(N__25930),
            .I(N__25924));
    LocalMux I__4956 (
            .O(N__25927),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    LocalMux I__4955 (
            .O(N__25924),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    InMux I__4954 (
            .O(N__25919),
            .I(N__25913));
    InMux I__4953 (
            .O(N__25918),
            .I(N__25913));
    LocalMux I__4952 (
            .O(N__25913),
            .I(\b2v_inst11.count_clk_1_14 ));
    InMux I__4951 (
            .O(N__25910),
            .I(\b2v_inst11.un1_count_clk_2_cry_13 ));
    InMux I__4950 (
            .O(N__25907),
            .I(N__25904));
    LocalMux I__4949 (
            .O(N__25904),
            .I(\b2v_inst11.count_clkZ0Z_15 ));
    InMux I__4948 (
            .O(N__25901),
            .I(\b2v_inst11.un1_count_clk_2_cry_14 ));
    InMux I__4947 (
            .O(N__25898),
            .I(N__25892));
    InMux I__4946 (
            .O(N__25897),
            .I(N__25892));
    LocalMux I__4945 (
            .O(N__25892),
            .I(\b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ));
    InMux I__4944 (
            .O(N__25889),
            .I(N__25886));
    LocalMux I__4943 (
            .O(N__25886),
            .I(\b2v_inst11.count_clk_0_11 ));
    InMux I__4942 (
            .O(N__25883),
            .I(N__25879));
    InMux I__4941 (
            .O(N__25882),
            .I(N__25876));
    LocalMux I__4940 (
            .O(N__25879),
            .I(\b2v_inst11.count_clk_1_11 ));
    LocalMux I__4939 (
            .O(N__25876),
            .I(\b2v_inst11.count_clk_1_11 ));
    CascadeMux I__4938 (
            .O(N__25871),
            .I(\b2v_inst36.curr_state_7_0_cascade_ ));
    InMux I__4937 (
            .O(N__25868),
            .I(N__25865));
    LocalMux I__4936 (
            .O(N__25865),
            .I(N__25860));
    InMux I__4935 (
            .O(N__25864),
            .I(N__25857));
    InMux I__4934 (
            .O(N__25863),
            .I(N__25854));
    Odrv12 I__4933 (
            .O(N__25860),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    LocalMux I__4932 (
            .O(N__25857),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    LocalMux I__4931 (
            .O(N__25854),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    InMux I__4930 (
            .O(N__25847),
            .I(N__25841));
    InMux I__4929 (
            .O(N__25846),
            .I(N__25841));
    LocalMux I__4928 (
            .O(N__25841),
            .I(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ));
    InMux I__4927 (
            .O(N__25838),
            .I(\b2v_inst11.un1_count_clk_2_cry_2 ));
    CascadeMux I__4926 (
            .O(N__25835),
            .I(N__25832));
    InMux I__4925 (
            .O(N__25832),
            .I(N__25827));
    InMux I__4924 (
            .O(N__25831),
            .I(N__25822));
    InMux I__4923 (
            .O(N__25830),
            .I(N__25822));
    LocalMux I__4922 (
            .O(N__25827),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    LocalMux I__4921 (
            .O(N__25822),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    CascadeMux I__4920 (
            .O(N__25817),
            .I(N__25814));
    InMux I__4919 (
            .O(N__25814),
            .I(N__25808));
    InMux I__4918 (
            .O(N__25813),
            .I(N__25808));
    LocalMux I__4917 (
            .O(N__25808),
            .I(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ));
    InMux I__4916 (
            .O(N__25805),
            .I(\b2v_inst11.un1_count_clk_2_cry_3 ));
    InMux I__4915 (
            .O(N__25802),
            .I(N__25798));
    InMux I__4914 (
            .O(N__25801),
            .I(N__25795));
    LocalMux I__4913 (
            .O(N__25798),
            .I(N__25792));
    LocalMux I__4912 (
            .O(N__25795),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    Odrv4 I__4911 (
            .O(N__25792),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    CascadeMux I__4910 (
            .O(N__25787),
            .I(N__25784));
    InMux I__4909 (
            .O(N__25784),
            .I(N__25778));
    InMux I__4908 (
            .O(N__25783),
            .I(N__25778));
    LocalMux I__4907 (
            .O(N__25778),
            .I(N__25775));
    Odrv4 I__4906 (
            .O(N__25775),
            .I(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ));
    InMux I__4905 (
            .O(N__25772),
            .I(\b2v_inst11.un1_count_clk_2_cry_4 ));
    CascadeMux I__4904 (
            .O(N__25769),
            .I(N__25766));
    InMux I__4903 (
            .O(N__25766),
            .I(N__25761));
    InMux I__4902 (
            .O(N__25765),
            .I(N__25756));
    InMux I__4901 (
            .O(N__25764),
            .I(N__25756));
    LocalMux I__4900 (
            .O(N__25761),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    LocalMux I__4899 (
            .O(N__25756),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    CascadeMux I__4898 (
            .O(N__25751),
            .I(N__25748));
    InMux I__4897 (
            .O(N__25748),
            .I(N__25742));
    InMux I__4896 (
            .O(N__25747),
            .I(N__25742));
    LocalMux I__4895 (
            .O(N__25742),
            .I(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ));
    InMux I__4894 (
            .O(N__25739),
            .I(\b2v_inst11.un1_count_clk_2_cry_5 ));
    InMux I__4893 (
            .O(N__25736),
            .I(\b2v_inst11.un1_count_clk_2_cry_6 ));
    InMux I__4892 (
            .O(N__25733),
            .I(N__25729));
    InMux I__4891 (
            .O(N__25732),
            .I(N__25726));
    LocalMux I__4890 (
            .O(N__25729),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    LocalMux I__4889 (
            .O(N__25726),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    CascadeMux I__4888 (
            .O(N__25721),
            .I(N__25718));
    InMux I__4887 (
            .O(N__25718),
            .I(N__25712));
    InMux I__4886 (
            .O(N__25717),
            .I(N__25712));
    LocalMux I__4885 (
            .O(N__25712),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ));
    InMux I__4884 (
            .O(N__25709),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ));
    InMux I__4883 (
            .O(N__25706),
            .I(N__25702));
    InMux I__4882 (
            .O(N__25705),
            .I(N__25699));
    LocalMux I__4881 (
            .O(N__25702),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    LocalMux I__4880 (
            .O(N__25699),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    InMux I__4879 (
            .O(N__25694),
            .I(N__25688));
    InMux I__4878 (
            .O(N__25693),
            .I(N__25688));
    LocalMux I__4877 (
            .O(N__25688),
            .I(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ));
    InMux I__4876 (
            .O(N__25685),
            .I(bfn_8_16_0_));
    InMux I__4875 (
            .O(N__25682),
            .I(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ));
    InMux I__4874 (
            .O(N__25679),
            .I(N__25676));
    LocalMux I__4873 (
            .O(N__25676),
            .I(\b2v_inst11.count_clk_0_2 ));
    InMux I__4872 (
            .O(N__25673),
            .I(N__25670));
    LocalMux I__4871 (
            .O(N__25670),
            .I(\b2v_inst11.count_clk_0_3 ));
    InMux I__4870 (
            .O(N__25667),
            .I(N__25664));
    LocalMux I__4869 (
            .O(N__25664),
            .I(\b2v_inst11.count_clk_0_4 ));
    InMux I__4868 (
            .O(N__25661),
            .I(N__25658));
    LocalMux I__4867 (
            .O(N__25658),
            .I(\b2v_inst11.count_clk_0_6 ));
    InMux I__4866 (
            .O(N__25655),
            .I(N__25650));
    InMux I__4865 (
            .O(N__25654),
            .I(N__25647));
    InMux I__4864 (
            .O(N__25653),
            .I(N__25644));
    LocalMux I__4863 (
            .O(N__25650),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    LocalMux I__4862 (
            .O(N__25647),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    LocalMux I__4861 (
            .O(N__25644),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    CascadeMux I__4860 (
            .O(N__25637),
            .I(N__25634));
    InMux I__4859 (
            .O(N__25634),
            .I(N__25628));
    InMux I__4858 (
            .O(N__25633),
            .I(N__25628));
    LocalMux I__4857 (
            .O(N__25628),
            .I(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ));
    InMux I__4856 (
            .O(N__25625),
            .I(\b2v_inst11.un1_count_clk_2_cry_1 ));
    CascadeMux I__4855 (
            .O(N__25622),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ));
    InMux I__4854 (
            .O(N__25619),
            .I(N__25616));
    LocalMux I__4853 (
            .O(N__25616),
            .I(N__25613));
    Odrv4 I__4852 (
            .O(N__25613),
            .I(\b2v_inst11.count_clk_en_0 ));
    CascadeMux I__4851 (
            .O(N__25610),
            .I(\b2v_inst11.N_328_cascade_ ));
    InMux I__4850 (
            .O(N__25607),
            .I(N__25604));
    LocalMux I__4849 (
            .O(N__25604),
            .I(N__25601));
    Span12Mux_v I__4848 (
            .O(N__25601),
            .I(N__25598));
    Odrv12 I__4847 (
            .O(N__25598),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_0 ));
    CascadeMux I__4846 (
            .O(N__25595),
            .I(\b2v_inst11.count_clk_en_cascade_ ));
    InMux I__4845 (
            .O(N__25592),
            .I(N__25589));
    LocalMux I__4844 (
            .O(N__25589),
            .I(N__25586));
    Span4Mux_v I__4843 (
            .O(N__25586),
            .I(N__25583));
    Odrv4 I__4842 (
            .O(N__25583),
            .I(\b2v_inst11.N_218 ));
    CascadeMux I__4841 (
            .O(N__25580),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_329_N_cascade_ ));
    InMux I__4840 (
            .O(N__25577),
            .I(N__25574));
    LocalMux I__4839 (
            .O(N__25574),
            .I(\b2v_inst11.un1_func_state25_6_0_0 ));
    CascadeMux I__4838 (
            .O(N__25571),
            .I(\b2v_inst11.count_clk_RNIDQ4A1Z0Z_7_cascade_ ));
    CascadeMux I__4837 (
            .O(N__25568),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_ ));
    InMux I__4836 (
            .O(N__25565),
            .I(N__25562));
    LocalMux I__4835 (
            .O(N__25562),
            .I(\b2v_inst11.g0_4_2 ));
    InMux I__4834 (
            .O(N__25559),
            .I(N__25556));
    LocalMux I__4833 (
            .O(N__25556),
            .I(\b2v_inst11.g0_0_0 ));
    CascadeMux I__4832 (
            .O(N__25553),
            .I(N__25550));
    InMux I__4831 (
            .O(N__25550),
            .I(N__25544));
    InMux I__4830 (
            .O(N__25549),
            .I(N__25544));
    LocalMux I__4829 (
            .O(N__25544),
            .I(N__25541));
    Odrv4 I__4828 (
            .O(N__25541),
            .I(\b2v_inst11.un1_clk_100khz_36_and_i_o3_0_c_0 ));
    InMux I__4827 (
            .O(N__25538),
            .I(N__25535));
    LocalMux I__4826 (
            .O(N__25535),
            .I(\b2v_inst11.g0_0_0_1 ));
    InMux I__4825 (
            .O(N__25532),
            .I(N__25526));
    InMux I__4824 (
            .O(N__25531),
            .I(N__25526));
    LocalMux I__4823 (
            .O(N__25526),
            .I(N__25523));
    Span4Mux_h I__4822 (
            .O(N__25523),
            .I(N__25518));
    InMux I__4821 (
            .O(N__25522),
            .I(N__25513));
    InMux I__4820 (
            .O(N__25521),
            .I(N__25513));
    Span4Mux_v I__4819 (
            .O(N__25518),
            .I(N__25509));
    LocalMux I__4818 (
            .O(N__25513),
            .I(N__25506));
    InMux I__4817 (
            .O(N__25512),
            .I(N__25503));
    Odrv4 I__4816 (
            .O(N__25509),
            .I(\b2v_inst11.func_state_RNI8H551Z0Z_0 ));
    Odrv4 I__4815 (
            .O(N__25506),
            .I(\b2v_inst11.func_state_RNI8H551Z0Z_0 ));
    LocalMux I__4814 (
            .O(N__25503),
            .I(\b2v_inst11.func_state_RNI8H551Z0Z_0 ));
    CascadeMux I__4813 (
            .O(N__25496),
            .I(N__25493));
    InMux I__4812 (
            .O(N__25493),
            .I(N__25487));
    InMux I__4811 (
            .O(N__25492),
            .I(N__25487));
    LocalMux I__4810 (
            .O(N__25487),
            .I(N__25484));
    Span4Mux_h I__4809 (
            .O(N__25484),
            .I(N__25480));
    InMux I__4808 (
            .O(N__25483),
            .I(N__25476));
    Span4Mux_v I__4807 (
            .O(N__25480),
            .I(N__25473));
    InMux I__4806 (
            .O(N__25479),
            .I(N__25470));
    LocalMux I__4805 (
            .O(N__25476),
            .I(N__25467));
    Odrv4 I__4804 (
            .O(N__25473),
            .I(\b2v_inst11.func_state_RNIDUQ02Z0Z_1 ));
    LocalMux I__4803 (
            .O(N__25470),
            .I(\b2v_inst11.func_state_RNIDUQ02Z0Z_1 ));
    Odrv4 I__4802 (
            .O(N__25467),
            .I(\b2v_inst11.func_state_RNIDUQ02Z0Z_1 ));
    CascadeMux I__4801 (
            .O(N__25460),
            .I(N__25456));
    InMux I__4800 (
            .O(N__25459),
            .I(N__25444));
    InMux I__4799 (
            .O(N__25456),
            .I(N__25444));
    InMux I__4798 (
            .O(N__25455),
            .I(N__25439));
    InMux I__4797 (
            .O(N__25454),
            .I(N__25439));
    InMux I__4796 (
            .O(N__25453),
            .I(N__25430));
    InMux I__4795 (
            .O(N__25452),
            .I(N__25430));
    InMux I__4794 (
            .O(N__25451),
            .I(N__25430));
    InMux I__4793 (
            .O(N__25450),
            .I(N__25430));
    CascadeMux I__4792 (
            .O(N__25449),
            .I(N__25427));
    LocalMux I__4791 (
            .O(N__25444),
            .I(N__25419));
    LocalMux I__4790 (
            .O(N__25439),
            .I(N__25416));
    LocalMux I__4789 (
            .O(N__25430),
            .I(N__25411));
    InMux I__4788 (
            .O(N__25427),
            .I(N__25408));
    InMux I__4787 (
            .O(N__25426),
            .I(N__25403));
    InMux I__4786 (
            .O(N__25425),
            .I(N__25403));
    InMux I__4785 (
            .O(N__25424),
            .I(N__25398));
    InMux I__4784 (
            .O(N__25423),
            .I(N__25398));
    InMux I__4783 (
            .O(N__25422),
            .I(N__25395));
    Span4Mux_v I__4782 (
            .O(N__25419),
            .I(N__25392));
    Span4Mux_h I__4781 (
            .O(N__25416),
            .I(N__25389));
    InMux I__4780 (
            .O(N__25415),
            .I(N__25384));
    InMux I__4779 (
            .O(N__25414),
            .I(N__25384));
    Span4Mux_h I__4778 (
            .O(N__25411),
            .I(N__25381));
    LocalMux I__4777 (
            .O(N__25408),
            .I(N__25368));
    LocalMux I__4776 (
            .O(N__25403),
            .I(N__25368));
    LocalMux I__4775 (
            .O(N__25398),
            .I(N__25368));
    LocalMux I__4774 (
            .O(N__25395),
            .I(N__25368));
    Span4Mux_h I__4773 (
            .O(N__25392),
            .I(N__25368));
    Span4Mux_v I__4772 (
            .O(N__25389),
            .I(N__25368));
    LocalMux I__4771 (
            .O(N__25384),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ));
    Odrv4 I__4770 (
            .O(N__25381),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ));
    Odrv4 I__4769 (
            .O(N__25368),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ));
    CascadeMux I__4768 (
            .O(N__25361),
            .I(\b2v_inst11.dutycycle_eena_5_d_1_1_cascade_ ));
    CascadeMux I__4767 (
            .O(N__25358),
            .I(\b2v_inst11.dutycycle_eena_5_0_1_cascade_ ));
    InMux I__4766 (
            .O(N__25355),
            .I(N__25352));
    LocalMux I__4765 (
            .O(N__25352),
            .I(N__25349));
    Odrv4 I__4764 (
            .O(N__25349),
            .I(\b2v_inst11.un1_clk_100khz_36_and_i_0 ));
    InMux I__4763 (
            .O(N__25346),
            .I(N__25342));
    InMux I__4762 (
            .O(N__25345),
            .I(N__25339));
    LocalMux I__4761 (
            .O(N__25342),
            .I(N__25334));
    LocalMux I__4760 (
            .O(N__25339),
            .I(N__25334));
    Span4Mux_v I__4759 (
            .O(N__25334),
            .I(N__25331));
    Span4Mux_h I__4758 (
            .O(N__25331),
            .I(N__25328));
    Odrv4 I__4757 (
            .O(N__25328),
            .I(\b2v_inst11.dutycycle_RNI2IQ6CZ0Z_7 ));
    CascadeMux I__4756 (
            .O(N__25325),
            .I(\b2v_inst11.func_state_RNIDUQ02Z0Z_1_cascade_ ));
    InMux I__4755 (
            .O(N__25322),
            .I(N__25317));
    InMux I__4754 (
            .O(N__25321),
            .I(N__25313));
    InMux I__4753 (
            .O(N__25320),
            .I(N__25309));
    LocalMux I__4752 (
            .O(N__25317),
            .I(N__25306));
    InMux I__4751 (
            .O(N__25316),
            .I(N__25303));
    LocalMux I__4750 (
            .O(N__25313),
            .I(N__25298));
    InMux I__4749 (
            .O(N__25312),
            .I(N__25295));
    LocalMux I__4748 (
            .O(N__25309),
            .I(N__25290));
    Span4Mux_v I__4747 (
            .O(N__25306),
            .I(N__25290));
    LocalMux I__4746 (
            .O(N__25303),
            .I(N__25287));
    InMux I__4745 (
            .O(N__25302),
            .I(N__25282));
    InMux I__4744 (
            .O(N__25301),
            .I(N__25282));
    Odrv4 I__4743 (
            .O(N__25298),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0 ));
    LocalMux I__4742 (
            .O(N__25295),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0 ));
    Odrv4 I__4741 (
            .O(N__25290),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0 ));
    Odrv4 I__4740 (
            .O(N__25287),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0 ));
    LocalMux I__4739 (
            .O(N__25282),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0 ));
    CascadeMux I__4738 (
            .O(N__25271),
            .I(\b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf0_cascade_ ));
    InMux I__4737 (
            .O(N__25268),
            .I(N__25265));
    LocalMux I__4736 (
            .O(N__25265),
            .I(\b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf1 ));
    CascadeMux I__4735 (
            .O(N__25262),
            .I(\b2v_inst11.N_14_0_cascade_ ));
    CascadeMux I__4734 (
            .O(N__25259),
            .I(N__25256));
    InMux I__4733 (
            .O(N__25256),
            .I(N__25253));
    LocalMux I__4732 (
            .O(N__25253),
            .I(\b2v_inst11.g2_i_2 ));
    CascadeMux I__4731 (
            .O(N__25250),
            .I(N__25247));
    InMux I__4730 (
            .O(N__25247),
            .I(N__25241));
    InMux I__4729 (
            .O(N__25246),
            .I(N__25241));
    LocalMux I__4728 (
            .O(N__25241),
            .I(N__25235));
    InMux I__4727 (
            .O(N__25240),
            .I(N__25228));
    InMux I__4726 (
            .O(N__25239),
            .I(N__25228));
    InMux I__4725 (
            .O(N__25238),
            .I(N__25228));
    Odrv4 I__4724 (
            .O(N__25235),
            .I(\b2v_inst11.func_state_RNI_6Z0Z_0 ));
    LocalMux I__4723 (
            .O(N__25228),
            .I(\b2v_inst11.func_state_RNI_6Z0Z_0 ));
    CascadeMux I__4722 (
            .O(N__25223),
            .I(\b2v_inst11.N_395_cascade_ ));
    InMux I__4721 (
            .O(N__25220),
            .I(N__25212));
    InMux I__4720 (
            .O(N__25219),
            .I(N__25207));
    InMux I__4719 (
            .O(N__25218),
            .I(N__25207));
    InMux I__4718 (
            .O(N__25217),
            .I(N__25204));
    InMux I__4717 (
            .O(N__25216),
            .I(N__25201));
    InMux I__4716 (
            .O(N__25215),
            .I(N__25198));
    LocalMux I__4715 (
            .O(N__25212),
            .I(N__25193));
    LocalMux I__4714 (
            .O(N__25207),
            .I(N__25190));
    LocalMux I__4713 (
            .O(N__25204),
            .I(N__25187));
    LocalMux I__4712 (
            .O(N__25201),
            .I(N__25182));
    LocalMux I__4711 (
            .O(N__25198),
            .I(N__25182));
    InMux I__4710 (
            .O(N__25197),
            .I(N__25179));
    CascadeMux I__4709 (
            .O(N__25196),
            .I(N__25174));
    Span4Mux_h I__4708 (
            .O(N__25193),
            .I(N__25171));
    Span4Mux_h I__4707 (
            .O(N__25190),
            .I(N__25168));
    Span4Mux_h I__4706 (
            .O(N__25187),
            .I(N__25161));
    Span4Mux_v I__4705 (
            .O(N__25182),
            .I(N__25161));
    LocalMux I__4704 (
            .O(N__25179),
            .I(N__25161));
    InMux I__4703 (
            .O(N__25178),
            .I(N__25156));
    InMux I__4702 (
            .O(N__25177),
            .I(N__25156));
    InMux I__4701 (
            .O(N__25174),
            .I(N__25153));
    Odrv4 I__4700 (
            .O(N__25171),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv4 I__4699 (
            .O(N__25168),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv4 I__4698 (
            .O(N__25161),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__4697 (
            .O(N__25156),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__4696 (
            .O(N__25153),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    CascadeMux I__4695 (
            .O(N__25142),
            .I(N__25135));
    CascadeMux I__4694 (
            .O(N__25141),
            .I(N__25131));
    CascadeMux I__4693 (
            .O(N__25140),
            .I(N__25128));
    InMux I__4692 (
            .O(N__25139),
            .I(N__25125));
    InMux I__4691 (
            .O(N__25138),
            .I(N__25116));
    InMux I__4690 (
            .O(N__25135),
            .I(N__25116));
    InMux I__4689 (
            .O(N__25134),
            .I(N__25116));
    InMux I__4688 (
            .O(N__25131),
            .I(N__25116));
    InMux I__4687 (
            .O(N__25128),
            .I(N__25113));
    LocalMux I__4686 (
            .O(N__25125),
            .I(N__25104));
    LocalMux I__4685 (
            .O(N__25116),
            .I(N__25104));
    LocalMux I__4684 (
            .O(N__25113),
            .I(N__25104));
    InMux I__4683 (
            .O(N__25112),
            .I(N__25099));
    InMux I__4682 (
            .O(N__25111),
            .I(N__25099));
    Span4Mux_v I__4681 (
            .O(N__25104),
            .I(N__25096));
    LocalMux I__4680 (
            .O(N__25099),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    Odrv4 I__4679 (
            .O(N__25096),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    CascadeMux I__4678 (
            .O(N__25091),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ));
    CascadeMux I__4677 (
            .O(N__25088),
            .I(N__25082));
    InMux I__4676 (
            .O(N__25087),
            .I(N__25076));
    InMux I__4675 (
            .O(N__25086),
            .I(N__25071));
    InMux I__4674 (
            .O(N__25085),
            .I(N__25071));
    InMux I__4673 (
            .O(N__25082),
            .I(N__25068));
    InMux I__4672 (
            .O(N__25081),
            .I(N__25065));
    InMux I__4671 (
            .O(N__25080),
            .I(N__25062));
    CascadeMux I__4670 (
            .O(N__25079),
            .I(N__25057));
    LocalMux I__4669 (
            .O(N__25076),
            .I(N__25053));
    LocalMux I__4668 (
            .O(N__25071),
            .I(N__25050));
    LocalMux I__4667 (
            .O(N__25068),
            .I(N__25043));
    LocalMux I__4666 (
            .O(N__25065),
            .I(N__25043));
    LocalMux I__4665 (
            .O(N__25062),
            .I(N__25043));
    InMux I__4664 (
            .O(N__25061),
            .I(N__25038));
    InMux I__4663 (
            .O(N__25060),
            .I(N__25038));
    InMux I__4662 (
            .O(N__25057),
            .I(N__25030));
    InMux I__4661 (
            .O(N__25056),
            .I(N__25030));
    Span4Mux_h I__4660 (
            .O(N__25053),
            .I(N__25027));
    Span4Mux_h I__4659 (
            .O(N__25050),
            .I(N__25020));
    Span4Mux_v I__4658 (
            .O(N__25043),
            .I(N__25020));
    LocalMux I__4657 (
            .O(N__25038),
            .I(N__25020));
    InMux I__4656 (
            .O(N__25037),
            .I(N__25017));
    InMux I__4655 (
            .O(N__25036),
            .I(N__25012));
    InMux I__4654 (
            .O(N__25035),
            .I(N__25012));
    LocalMux I__4653 (
            .O(N__25030),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__4652 (
            .O(N__25027),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__4651 (
            .O(N__25020),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__4650 (
            .O(N__25017),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__4649 (
            .O(N__25012),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    CascadeMux I__4648 (
            .O(N__25001),
            .I(\b2v_inst11.N_365_cascade_ ));
    CascadeMux I__4647 (
            .O(N__24998),
            .I(\b2v_inst11.N_366_cascade_ ));
    InMux I__4646 (
            .O(N__24995),
            .I(N__24988));
    InMux I__4645 (
            .O(N__24994),
            .I(N__24988));
    InMux I__4644 (
            .O(N__24993),
            .I(N__24983));
    LocalMux I__4643 (
            .O(N__24988),
            .I(N__24980));
    InMux I__4642 (
            .O(N__24987),
            .I(N__24977));
    InMux I__4641 (
            .O(N__24986),
            .I(N__24974));
    LocalMux I__4640 (
            .O(N__24983),
            .I(N__24969));
    Span4Mux_v I__4639 (
            .O(N__24980),
            .I(N__24969));
    LocalMux I__4638 (
            .O(N__24977),
            .I(N__24964));
    LocalMux I__4637 (
            .O(N__24974),
            .I(N__24964));
    Span4Mux_v I__4636 (
            .O(N__24969),
            .I(N__24961));
    Odrv4 I__4635 (
            .O(N__24964),
            .I(\b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1 ));
    Odrv4 I__4634 (
            .O(N__24961),
            .I(\b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1 ));
    InMux I__4633 (
            .O(N__24956),
            .I(N__24952));
    InMux I__4632 (
            .O(N__24955),
            .I(N__24947));
    LocalMux I__4631 (
            .O(N__24952),
            .I(N__24944));
    InMux I__4630 (
            .O(N__24951),
            .I(N__24940));
    CascadeMux I__4629 (
            .O(N__24950),
            .I(N__24936));
    LocalMux I__4628 (
            .O(N__24947),
            .I(N__24932));
    Span4Mux_v I__4627 (
            .O(N__24944),
            .I(N__24929));
    InMux I__4626 (
            .O(N__24943),
            .I(N__24926));
    LocalMux I__4625 (
            .O(N__24940),
            .I(N__24923));
    InMux I__4624 (
            .O(N__24939),
            .I(N__24918));
    InMux I__4623 (
            .O(N__24936),
            .I(N__24918));
    CascadeMux I__4622 (
            .O(N__24935),
            .I(N__24913));
    Span4Mux_v I__4621 (
            .O(N__24932),
            .I(N__24908));
    Span4Mux_h I__4620 (
            .O(N__24929),
            .I(N__24908));
    LocalMux I__4619 (
            .O(N__24926),
            .I(N__24905));
    Span4Mux_h I__4618 (
            .O(N__24923),
            .I(N__24902));
    LocalMux I__4617 (
            .O(N__24918),
            .I(N__24899));
    InMux I__4616 (
            .O(N__24917),
            .I(N__24896));
    InMux I__4615 (
            .O(N__24916),
            .I(N__24893));
    InMux I__4614 (
            .O(N__24913),
            .I(N__24890));
    Odrv4 I__4613 (
            .O(N__24908),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__4612 (
            .O(N__24905),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__4611 (
            .O(N__24902),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv12 I__4610 (
            .O(N__24899),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__4609 (
            .O(N__24896),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__4608 (
            .O(N__24893),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__4607 (
            .O(N__24890),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    CascadeMux I__4606 (
            .O(N__24875),
            .I(N__24872));
    InMux I__4605 (
            .O(N__24872),
            .I(N__24869));
    LocalMux I__4604 (
            .O(N__24869),
            .I(\b2v_inst11.N_153_N ));
    InMux I__4603 (
            .O(N__24866),
            .I(N__24863));
    LocalMux I__4602 (
            .O(N__24863),
            .I(N__24860));
    Span4Mux_v I__4601 (
            .O(N__24860),
            .I(N__24857));
    Odrv4 I__4600 (
            .O(N__24857),
            .I(\b2v_inst11.g2_i_a6_0 ));
    InMux I__4599 (
            .O(N__24854),
            .I(N__24850));
    InMux I__4598 (
            .O(N__24853),
            .I(N__24847));
    LocalMux I__4597 (
            .O(N__24850),
            .I(N__24844));
    LocalMux I__4596 (
            .O(N__24847),
            .I(N__24841));
    Span4Mux_v I__4595 (
            .O(N__24844),
            .I(N__24838));
    Span4Mux_v I__4594 (
            .O(N__24841),
            .I(N__24835));
    Span4Mux_h I__4593 (
            .O(N__24838),
            .I(N__24830));
    Span4Mux_h I__4592 (
            .O(N__24835),
            .I(N__24830));
    Odrv4 I__4591 (
            .O(N__24830),
            .I(\b2v_inst11.N_363 ));
    InMux I__4590 (
            .O(N__24827),
            .I(N__24824));
    LocalMux I__4589 (
            .O(N__24824),
            .I(N__24821));
    Odrv4 I__4588 (
            .O(N__24821),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ));
    CascadeMux I__4587 (
            .O(N__24818),
            .I(\b2v_inst11.N_396_N_cascade_ ));
    CascadeMux I__4586 (
            .O(N__24815),
            .I(\b2v_inst11.N_234_N_cascade_ ));
    InMux I__4585 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__4584 (
            .O(N__24809),
            .I(N__24806));
    Odrv4 I__4583 (
            .O(N__24806),
            .I(\b2v_inst11.dutycycle_eena_9 ));
    InMux I__4582 (
            .O(N__24803),
            .I(N__24800));
    LocalMux I__4581 (
            .O(N__24800),
            .I(N__24796));
    InMux I__4580 (
            .O(N__24799),
            .I(N__24793));
    Odrv4 I__4579 (
            .O(N__24796),
            .I(\b2v_inst11.dutycycle_rst_8 ));
    LocalMux I__4578 (
            .O(N__24793),
            .I(\b2v_inst11.dutycycle_rst_8 ));
    InMux I__4577 (
            .O(N__24788),
            .I(N__24782));
    InMux I__4576 (
            .O(N__24787),
            .I(N__24782));
    LocalMux I__4575 (
            .O(N__24782),
            .I(\b2v_inst11.dutycycleZ1Z_12 ));
    CascadeMux I__4574 (
            .O(N__24779),
            .I(\b2v_inst11.dutycycle_eena_9_cascade_ ));
    CascadeMux I__4573 (
            .O(N__24776),
            .I(N__24773));
    InMux I__4572 (
            .O(N__24773),
            .I(N__24770));
    LocalMux I__4571 (
            .O(N__24770),
            .I(\b2v_inst11.N_234_N ));
    InMux I__4570 (
            .O(N__24767),
            .I(N__24764));
    LocalMux I__4569 (
            .O(N__24764),
            .I(\b2v_inst11.dutycycle_eena_7 ));
    CascadeMux I__4568 (
            .O(N__24761),
            .I(N__24758));
    InMux I__4567 (
            .O(N__24758),
            .I(N__24755));
    LocalMux I__4566 (
            .O(N__24755),
            .I(N__24751));
    InMux I__4565 (
            .O(N__24754),
            .I(N__24748));
    Odrv4 I__4564 (
            .O(N__24751),
            .I(\b2v_inst11.dutycycleZ1Z_11 ));
    LocalMux I__4563 (
            .O(N__24748),
            .I(\b2v_inst11.dutycycleZ1Z_11 ));
    CascadeMux I__4562 (
            .O(N__24743),
            .I(\b2v_inst11.dutycycle_eena_7_cascade_ ));
    InMux I__4561 (
            .O(N__24740),
            .I(N__24734));
    InMux I__4560 (
            .O(N__24739),
            .I(N__24734));
    LocalMux I__4559 (
            .O(N__24734),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUFZ0Z1 ));
    CascadeMux I__4558 (
            .O(N__24731),
            .I(N__24728));
    InMux I__4557 (
            .O(N__24728),
            .I(N__24722));
    InMux I__4556 (
            .O(N__24727),
            .I(N__24722));
    LocalMux I__4555 (
            .O(N__24722),
            .I(N__24719));
    Span4Mux_h I__4554 (
            .O(N__24719),
            .I(N__24716));
    Odrv4 I__4553 (
            .O(N__24716),
            .I(\b2v_inst11.dutycycle_RNIT35D7Z0Z_13 ));
    CascadeMux I__4552 (
            .O(N__24713),
            .I(N__24708));
    InMux I__4551 (
            .O(N__24712),
            .I(N__24705));
    CascadeMux I__4550 (
            .O(N__24711),
            .I(N__24700));
    InMux I__4549 (
            .O(N__24708),
            .I(N__24696));
    LocalMux I__4548 (
            .O(N__24705),
            .I(N__24693));
    InMux I__4547 (
            .O(N__24704),
            .I(N__24690));
    CascadeMux I__4546 (
            .O(N__24703),
            .I(N__24685));
    InMux I__4545 (
            .O(N__24700),
            .I(N__24680));
    InMux I__4544 (
            .O(N__24699),
            .I(N__24680));
    LocalMux I__4543 (
            .O(N__24696),
            .I(N__24677));
    Span4Mux_h I__4542 (
            .O(N__24693),
            .I(N__24671));
    LocalMux I__4541 (
            .O(N__24690),
            .I(N__24671));
    InMux I__4540 (
            .O(N__24689),
            .I(N__24666));
    InMux I__4539 (
            .O(N__24688),
            .I(N__24666));
    InMux I__4538 (
            .O(N__24685),
            .I(N__24663));
    LocalMux I__4537 (
            .O(N__24680),
            .I(N__24658));
    Span4Mux_v I__4536 (
            .O(N__24677),
            .I(N__24658));
    InMux I__4535 (
            .O(N__24676),
            .I(N__24655));
    Odrv4 I__4534 (
            .O(N__24671),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    LocalMux I__4533 (
            .O(N__24666),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    LocalMux I__4532 (
            .O(N__24663),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    Odrv4 I__4531 (
            .O(N__24658),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    LocalMux I__4530 (
            .O(N__24655),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    InMux I__4529 (
            .O(N__24644),
            .I(N__24641));
    LocalMux I__4528 (
            .O(N__24641),
            .I(N__24638));
    Span4Mux_h I__4527 (
            .O(N__24638),
            .I(N__24635));
    Odrv4 I__4526 (
            .O(N__24635),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_11 ));
    InMux I__4525 (
            .O(N__24632),
            .I(N__24624));
    CascadeMux I__4524 (
            .O(N__24631),
            .I(N__24617));
    InMux I__4523 (
            .O(N__24630),
            .I(N__24614));
    InMux I__4522 (
            .O(N__24629),
            .I(N__24609));
    InMux I__4521 (
            .O(N__24628),
            .I(N__24609));
    CascadeMux I__4520 (
            .O(N__24627),
            .I(N__24605));
    LocalMux I__4519 (
            .O(N__24624),
            .I(N__24602));
    InMux I__4518 (
            .O(N__24623),
            .I(N__24599));
    CascadeMux I__4517 (
            .O(N__24622),
            .I(N__24592));
    CascadeMux I__4516 (
            .O(N__24621),
            .I(N__24589));
    InMux I__4515 (
            .O(N__24620),
            .I(N__24583));
    InMux I__4514 (
            .O(N__24617),
            .I(N__24583));
    LocalMux I__4513 (
            .O(N__24614),
            .I(N__24580));
    LocalMux I__4512 (
            .O(N__24609),
            .I(N__24577));
    InMux I__4511 (
            .O(N__24608),
            .I(N__24572));
    InMux I__4510 (
            .O(N__24605),
            .I(N__24572));
    Span4Mux_v I__4509 (
            .O(N__24602),
            .I(N__24569));
    LocalMux I__4508 (
            .O(N__24599),
            .I(N__24564));
    InMux I__4507 (
            .O(N__24598),
            .I(N__24561));
    InMux I__4506 (
            .O(N__24597),
            .I(N__24558));
    CascadeMux I__4505 (
            .O(N__24596),
            .I(N__24552));
    InMux I__4504 (
            .O(N__24595),
            .I(N__24543));
    InMux I__4503 (
            .O(N__24592),
            .I(N__24543));
    InMux I__4502 (
            .O(N__24589),
            .I(N__24543));
    InMux I__4501 (
            .O(N__24588),
            .I(N__24543));
    LocalMux I__4500 (
            .O(N__24583),
            .I(N__24540));
    Span4Mux_h I__4499 (
            .O(N__24580),
            .I(N__24537));
    Span4Mux_v I__4498 (
            .O(N__24577),
            .I(N__24530));
    LocalMux I__4497 (
            .O(N__24572),
            .I(N__24530));
    Span4Mux_s3_h I__4496 (
            .O(N__24569),
            .I(N__24530));
    InMux I__4495 (
            .O(N__24568),
            .I(N__24525));
    InMux I__4494 (
            .O(N__24567),
            .I(N__24525));
    Span4Mux_v I__4493 (
            .O(N__24564),
            .I(N__24518));
    LocalMux I__4492 (
            .O(N__24561),
            .I(N__24518));
    LocalMux I__4491 (
            .O(N__24558),
            .I(N__24518));
    InMux I__4490 (
            .O(N__24557),
            .I(N__24511));
    InMux I__4489 (
            .O(N__24556),
            .I(N__24511));
    InMux I__4488 (
            .O(N__24555),
            .I(N__24511));
    InMux I__4487 (
            .O(N__24552),
            .I(N__24508));
    LocalMux I__4486 (
            .O(N__24543),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__4485 (
            .O(N__24540),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__4484 (
            .O(N__24537),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__4483 (
            .O(N__24530),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    LocalMux I__4482 (
            .O(N__24525),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__4481 (
            .O(N__24518),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    LocalMux I__4480 (
            .O(N__24511),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    LocalMux I__4479 (
            .O(N__24508),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    CascadeMux I__4478 (
            .O(N__24491),
            .I(N__24488));
    InMux I__4477 (
            .O(N__24488),
            .I(N__24485));
    LocalMux I__4476 (
            .O(N__24485),
            .I(N__24482));
    Odrv4 I__4475 (
            .O(N__24482),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_5 ));
    CascadeMux I__4474 (
            .O(N__24479),
            .I(\b2v_inst5.count_rst_6_cascade_ ));
    CascadeMux I__4473 (
            .O(N__24476),
            .I(N__24473));
    InMux I__4472 (
            .O(N__24473),
            .I(N__24469));
    InMux I__4471 (
            .O(N__24472),
            .I(N__24466));
    LocalMux I__4470 (
            .O(N__24469),
            .I(\b2v_inst5.un2_count_1_axb_8 ));
    LocalMux I__4469 (
            .O(N__24466),
            .I(\b2v_inst5.un2_count_1_axb_8 ));
    InMux I__4468 (
            .O(N__24461),
            .I(N__24455));
    InMux I__4467 (
            .O(N__24460),
            .I(N__24455));
    LocalMux I__4466 (
            .O(N__24455),
            .I(\b2v_inst5.un2_count_1_cry_7_THRU_CO ));
    CascadeMux I__4465 (
            .O(N__24452),
            .I(\b2v_inst5.un2_count_1_axb_8_cascade_ ));
    InMux I__4464 (
            .O(N__24449),
            .I(N__24443));
    InMux I__4463 (
            .O(N__24448),
            .I(N__24443));
    LocalMux I__4462 (
            .O(N__24443),
            .I(\b2v_inst5.count_1_8 ));
    CascadeMux I__4461 (
            .O(N__24440),
            .I(\b2v_inst5.count_rst_10_cascade_ ));
    InMux I__4460 (
            .O(N__24437),
            .I(N__24434));
    LocalMux I__4459 (
            .O(N__24434),
            .I(N__24429));
    InMux I__4458 (
            .O(N__24433),
            .I(N__24424));
    InMux I__4457 (
            .O(N__24432),
            .I(N__24424));
    Span4Mux_h I__4456 (
            .O(N__24429),
            .I(N__24421));
    LocalMux I__4455 (
            .O(N__24424),
            .I(\b2v_inst5.countZ0Z_4 ));
    Odrv4 I__4454 (
            .O(N__24421),
            .I(\b2v_inst5.countZ0Z_4 ));
    CascadeMux I__4453 (
            .O(N__24416),
            .I(N__24412));
    InMux I__4452 (
            .O(N__24415),
            .I(N__24407));
    InMux I__4451 (
            .O(N__24412),
            .I(N__24407));
    LocalMux I__4450 (
            .O(N__24407),
            .I(N__24404));
    Span4Mux_h I__4449 (
            .O(N__24404),
            .I(N__24401));
    Odrv4 I__4448 (
            .O(N__24401),
            .I(\b2v_inst5.un2_count_1_cry_3_THRU_CO ));
    CascadeMux I__4447 (
            .O(N__24398),
            .I(\b2v_inst5.countZ0Z_4_cascade_ ));
    InMux I__4446 (
            .O(N__24395),
            .I(N__24392));
    LocalMux I__4445 (
            .O(N__24392),
            .I(\b2v_inst5.count_1_4 ));
    InMux I__4444 (
            .O(N__24389),
            .I(N__24385));
    InMux I__4443 (
            .O(N__24388),
            .I(N__24382));
    LocalMux I__4442 (
            .O(N__24385),
            .I(\b2v_inst5.un2_count_1_cry_12_THRU_CO ));
    LocalMux I__4441 (
            .O(N__24382),
            .I(\b2v_inst5.un2_count_1_cry_12_THRU_CO ));
    InMux I__4440 (
            .O(N__24377),
            .I(N__24374));
    LocalMux I__4439 (
            .O(N__24374),
            .I(\b2v_inst5.count_rst_1 ));
    CascadeMux I__4438 (
            .O(N__24371),
            .I(\b2v_inst5.countZ0Z_13_cascade_ ));
    InMux I__4437 (
            .O(N__24368),
            .I(N__24365));
    LocalMux I__4436 (
            .O(N__24365),
            .I(\b2v_inst5.count_1_13 ));
    CascadeMux I__4435 (
            .O(N__24362),
            .I(\b2v_inst5.count_i_0_cascade_ ));
    InMux I__4434 (
            .O(N__24359),
            .I(N__24356));
    LocalMux I__4433 (
            .O(N__24356),
            .I(\b2v_inst5.count_rst_14 ));
    InMux I__4432 (
            .O(N__24353),
            .I(N__24347));
    InMux I__4431 (
            .O(N__24352),
            .I(N__24347));
    LocalMux I__4430 (
            .O(N__24347),
            .I(\b2v_inst5.count_1_0 ));
    CascadeMux I__4429 (
            .O(N__24344),
            .I(\b2v_inst5.count_rst_14_cascade_ ));
    CascadeMux I__4428 (
            .O(N__24341),
            .I(N__24338));
    InMux I__4427 (
            .O(N__24338),
            .I(N__24335));
    LocalMux I__4426 (
            .O(N__24335),
            .I(\b2v_inst5.un2_count_1_axb_0 ));
    InMux I__4425 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__4424 (
            .O(N__24329),
            .I(N__24325));
    InMux I__4423 (
            .O(N__24328),
            .I(N__24322));
    Odrv12 I__4422 (
            .O(N__24325),
            .I(\b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2 ));
    LocalMux I__4421 (
            .O(N__24322),
            .I(\b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2 ));
    InMux I__4420 (
            .O(N__24317),
            .I(N__24314));
    LocalMux I__4419 (
            .O(N__24314),
            .I(N__24311));
    Odrv4 I__4418 (
            .O(N__24311),
            .I(\b2v_inst5.count_1_14 ));
    InMux I__4417 (
            .O(N__24308),
            .I(N__24305));
    LocalMux I__4416 (
            .O(N__24305),
            .I(\b2v_inst5.countZ0Z_14 ));
    InMux I__4415 (
            .O(N__24302),
            .I(N__24296));
    InMux I__4414 (
            .O(N__24301),
            .I(N__24296));
    LocalMux I__4413 (
            .O(N__24296),
            .I(\b2v_inst5.count_i_0 ));
    CascadeMux I__4412 (
            .O(N__24293),
            .I(\b2v_inst5.countZ0Z_14_cascade_ ));
    InMux I__4411 (
            .O(N__24290),
            .I(N__24286));
    InMux I__4410 (
            .O(N__24289),
            .I(N__24283));
    LocalMux I__4409 (
            .O(N__24286),
            .I(N__24280));
    LocalMux I__4408 (
            .O(N__24283),
            .I(N__24277));
    Odrv4 I__4407 (
            .O(N__24280),
            .I(\b2v_inst5.countZ0Z_12 ));
    Odrv4 I__4406 (
            .O(N__24277),
            .I(\b2v_inst5.countZ0Z_12 ));
    InMux I__4405 (
            .O(N__24272),
            .I(N__24269));
    LocalMux I__4404 (
            .O(N__24269),
            .I(N__24266));
    Odrv4 I__4403 (
            .O(N__24266),
            .I(\b2v_inst5.count_rst_6 ));
    InMux I__4402 (
            .O(N__24263),
            .I(N__24257));
    InMux I__4401 (
            .O(N__24262),
            .I(N__24257));
    LocalMux I__4400 (
            .O(N__24257),
            .I(N__24254));
    Odrv4 I__4399 (
            .O(N__24254),
            .I(\b2v_inst36.count_rst ));
    InMux I__4398 (
            .O(N__24251),
            .I(N__24248));
    LocalMux I__4397 (
            .O(N__24248),
            .I(N__24245));
    Span4Mux_v I__4396 (
            .O(N__24245),
            .I(N__24242));
    Odrv4 I__4395 (
            .O(N__24242),
            .I(\b2v_inst20.counter_1_cry_1_THRU_CO ));
    InMux I__4394 (
            .O(N__24239),
            .I(N__24235));
    InMux I__4393 (
            .O(N__24238),
            .I(N__24232));
    LocalMux I__4392 (
            .O(N__24235),
            .I(N__24229));
    LocalMux I__4391 (
            .O(N__24232),
            .I(N__24223));
    Span4Mux_h I__4390 (
            .O(N__24229),
            .I(N__24223));
    InMux I__4389 (
            .O(N__24228),
            .I(N__24220));
    Odrv4 I__4388 (
            .O(N__24223),
            .I(\b2v_inst20.counterZ0Z_2 ));
    LocalMux I__4387 (
            .O(N__24220),
            .I(\b2v_inst20.counterZ0Z_2 ));
    CascadeMux I__4386 (
            .O(N__24215),
            .I(\b2v_inst36.curr_state_RNI3E27Z0Z_0_cascade_ ));
    IoInMux I__4385 (
            .O(N__24212),
            .I(N__24209));
    LocalMux I__4384 (
            .O(N__24209),
            .I(N__24206));
    Span4Mux_s3_h I__4383 (
            .O(N__24206),
            .I(N__24203));
    Span4Mux_h I__4382 (
            .O(N__24203),
            .I(N__24200));
    Span4Mux_v I__4381 (
            .O(N__24200),
            .I(N__24197));
    Odrv4 I__4380 (
            .O(N__24197),
            .I(dsw_pwrok));
    CascadeMux I__4379 (
            .O(N__24194),
            .I(N__24187));
    InMux I__4378 (
            .O(N__24193),
            .I(N__24176));
    InMux I__4377 (
            .O(N__24192),
            .I(N__24176));
    InMux I__4376 (
            .O(N__24191),
            .I(N__24176));
    InMux I__4375 (
            .O(N__24190),
            .I(N__24176));
    InMux I__4374 (
            .O(N__24187),
            .I(N__24176));
    LocalMux I__4373 (
            .O(N__24176),
            .I(N__24167));
    InMux I__4372 (
            .O(N__24175),
            .I(N__24164));
    InMux I__4371 (
            .O(N__24174),
            .I(N__24153));
    InMux I__4370 (
            .O(N__24173),
            .I(N__24153));
    InMux I__4369 (
            .O(N__24172),
            .I(N__24153));
    InMux I__4368 (
            .O(N__24171),
            .I(N__24153));
    InMux I__4367 (
            .O(N__24170),
            .I(N__24153));
    Span4Mux_v I__4366 (
            .O(N__24167),
            .I(N__24150));
    LocalMux I__4365 (
            .O(N__24164),
            .I(N__24145));
    LocalMux I__4364 (
            .O(N__24153),
            .I(N__24145));
    Odrv4 I__4363 (
            .O(N__24150),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    Odrv4 I__4362 (
            .O(N__24145),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    InMux I__4361 (
            .O(N__24140),
            .I(N__24137));
    LocalMux I__4360 (
            .O(N__24137),
            .I(N__24134));
    Span4Mux_h I__4359 (
            .O(N__24134),
            .I(N__24131));
    Odrv4 I__4358 (
            .O(N__24131),
            .I(\b2v_inst20.counter_1_cry_2_THRU_CO ));
    InMux I__4357 (
            .O(N__24128),
            .I(N__24125));
    LocalMux I__4356 (
            .O(N__24125),
            .I(N__24121));
    InMux I__4355 (
            .O(N__24124),
            .I(N__24117));
    Span4Mux_h I__4354 (
            .O(N__24121),
            .I(N__24114));
    InMux I__4353 (
            .O(N__24120),
            .I(N__24111));
    LocalMux I__4352 (
            .O(N__24117),
            .I(\b2v_inst20.counterZ0Z_3 ));
    Odrv4 I__4351 (
            .O(N__24114),
            .I(\b2v_inst20.counterZ0Z_3 ));
    LocalMux I__4350 (
            .O(N__24111),
            .I(\b2v_inst20.counterZ0Z_3 ));
    CascadeMux I__4349 (
            .O(N__24104),
            .I(N__24100));
    InMux I__4348 (
            .O(N__24103),
            .I(N__24094));
    InMux I__4347 (
            .O(N__24100),
            .I(N__24094));
    InMux I__4346 (
            .O(N__24099),
            .I(N__24091));
    LocalMux I__4345 (
            .O(N__24094),
            .I(\b2v_inst36.un2_count_1_axb_7 ));
    LocalMux I__4344 (
            .O(N__24091),
            .I(\b2v_inst36.un2_count_1_axb_7 ));
    CascadeMux I__4343 (
            .O(N__24086),
            .I(N__24083));
    InMux I__4342 (
            .O(N__24083),
            .I(N__24079));
    InMux I__4341 (
            .O(N__24082),
            .I(N__24076));
    LocalMux I__4340 (
            .O(N__24079),
            .I(N__24073));
    LocalMux I__4339 (
            .O(N__24076),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    Odrv4 I__4338 (
            .O(N__24073),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    InMux I__4337 (
            .O(N__24068),
            .I(\b2v_inst36.un2_count_1_cry_6 ));
    InMux I__4336 (
            .O(N__24065),
            .I(bfn_8_4_0_));
    InMux I__4335 (
            .O(N__24062),
            .I(\b2v_inst36.un2_count_1_cry_8 ));
    InMux I__4334 (
            .O(N__24059),
            .I(\b2v_inst36.un2_count_1_cry_9 ));
    InMux I__4333 (
            .O(N__24056),
            .I(N__24051));
    InMux I__4332 (
            .O(N__24055),
            .I(N__24046));
    InMux I__4331 (
            .O(N__24054),
            .I(N__24046));
    LocalMux I__4330 (
            .O(N__24051),
            .I(N__24043));
    LocalMux I__4329 (
            .O(N__24046),
            .I(\b2v_inst36.countZ0Z_11 ));
    Odrv4 I__4328 (
            .O(N__24043),
            .I(\b2v_inst36.countZ0Z_11 ));
    CascadeMux I__4327 (
            .O(N__24038),
            .I(N__24034));
    InMux I__4326 (
            .O(N__24037),
            .I(N__24029));
    InMux I__4325 (
            .O(N__24034),
            .I(N__24029));
    LocalMux I__4324 (
            .O(N__24029),
            .I(N__24026));
    Odrv4 I__4323 (
            .O(N__24026),
            .I(\b2v_inst36.un2_count_1_cry_10_THRU_CO ));
    InMux I__4322 (
            .O(N__24023),
            .I(\b2v_inst36.un2_count_1_cry_10 ));
    InMux I__4321 (
            .O(N__24020),
            .I(\b2v_inst36.un2_count_1_cry_11 ));
    InMux I__4320 (
            .O(N__24017),
            .I(N__24013));
    InMux I__4319 (
            .O(N__24016),
            .I(N__24010));
    LocalMux I__4318 (
            .O(N__24013),
            .I(N__24007));
    LocalMux I__4317 (
            .O(N__24010),
            .I(\b2v_inst36.countZ0Z_13 ));
    Odrv4 I__4316 (
            .O(N__24007),
            .I(\b2v_inst36.countZ0Z_13 ));
    InMux I__4315 (
            .O(N__24002),
            .I(N__23996));
    InMux I__4314 (
            .O(N__24001),
            .I(N__23996));
    LocalMux I__4313 (
            .O(N__23996),
            .I(N__23993));
    Odrv4 I__4312 (
            .O(N__23993),
            .I(\b2v_inst36.count_rst_1 ));
    InMux I__4311 (
            .O(N__23990),
            .I(\b2v_inst36.un2_count_1_cry_12 ));
    InMux I__4310 (
            .O(N__23987),
            .I(N__23983));
    InMux I__4309 (
            .O(N__23986),
            .I(N__23980));
    LocalMux I__4308 (
            .O(N__23983),
            .I(N__23977));
    LocalMux I__4307 (
            .O(N__23980),
            .I(\b2v_inst36.countZ0Z_14 ));
    Odrv4 I__4306 (
            .O(N__23977),
            .I(\b2v_inst36.countZ0Z_14 ));
    InMux I__4305 (
            .O(N__23972),
            .I(N__23966));
    InMux I__4304 (
            .O(N__23971),
            .I(N__23966));
    LocalMux I__4303 (
            .O(N__23966),
            .I(N__23963));
    Span4Mux_h I__4302 (
            .O(N__23963),
            .I(N__23960));
    Odrv4 I__4301 (
            .O(N__23960),
            .I(\b2v_inst36.count_rst_0 ));
    InMux I__4300 (
            .O(N__23957),
            .I(\b2v_inst36.un2_count_1_cry_13 ));
    InMux I__4299 (
            .O(N__23954),
            .I(N__23951));
    LocalMux I__4298 (
            .O(N__23951),
            .I(N__23947));
    InMux I__4297 (
            .O(N__23950),
            .I(N__23944));
    Odrv4 I__4296 (
            .O(N__23947),
            .I(\b2v_inst36.countZ0Z_15 ));
    LocalMux I__4295 (
            .O(N__23944),
            .I(\b2v_inst36.countZ0Z_15 ));
    InMux I__4294 (
            .O(N__23939),
            .I(\b2v_inst36.un2_count_1_cry_14 ));
    InMux I__4293 (
            .O(N__23936),
            .I(N__23932));
    InMux I__4292 (
            .O(N__23935),
            .I(N__23929));
    LocalMux I__4291 (
            .O(N__23932),
            .I(\b2v_inst36.count_2_0 ));
    LocalMux I__4290 (
            .O(N__23929),
            .I(\b2v_inst36.count_2_0 ));
    InMux I__4289 (
            .O(N__23924),
            .I(N__23920));
    InMux I__4288 (
            .O(N__23923),
            .I(N__23917));
    LocalMux I__4287 (
            .O(N__23920),
            .I(\b2v_inst36.count_rst_14 ));
    LocalMux I__4286 (
            .O(N__23917),
            .I(\b2v_inst36.count_rst_14 ));
    InMux I__4285 (
            .O(N__23912),
            .I(N__23909));
    LocalMux I__4284 (
            .O(N__23909),
            .I(\b2v_inst36.un2_count_1_axb_0 ));
    InMux I__4283 (
            .O(N__23906),
            .I(N__23903));
    LocalMux I__4282 (
            .O(N__23903),
            .I(N__23900));
    Odrv4 I__4281 (
            .O(N__23900),
            .I(\b2v_inst36.un2_count_1_axb_1 ));
    InMux I__4280 (
            .O(N__23897),
            .I(N__23888));
    InMux I__4279 (
            .O(N__23896),
            .I(N__23888));
    InMux I__4278 (
            .O(N__23895),
            .I(N__23888));
    LocalMux I__4277 (
            .O(N__23888),
            .I(N__23885));
    Odrv4 I__4276 (
            .O(N__23885),
            .I(\b2v_inst36.count_rst_13 ));
    InMux I__4275 (
            .O(N__23882),
            .I(\b2v_inst36.un2_count_1_cry_0 ));
    InMux I__4274 (
            .O(N__23879),
            .I(N__23874));
    InMux I__4273 (
            .O(N__23878),
            .I(N__23869));
    InMux I__4272 (
            .O(N__23877),
            .I(N__23869));
    LocalMux I__4271 (
            .O(N__23874),
            .I(N__23866));
    LocalMux I__4270 (
            .O(N__23869),
            .I(\b2v_inst36.countZ0Z_2 ));
    Odrv4 I__4269 (
            .O(N__23866),
            .I(\b2v_inst36.countZ0Z_2 ));
    InMux I__4268 (
            .O(N__23861),
            .I(N__23855));
    InMux I__4267 (
            .O(N__23860),
            .I(N__23855));
    LocalMux I__4266 (
            .O(N__23855),
            .I(N__23852));
    Odrv4 I__4265 (
            .O(N__23852),
            .I(\b2v_inst36.un2_count_1_cry_1_THRU_CO ));
    InMux I__4264 (
            .O(N__23849),
            .I(\b2v_inst36.un2_count_1_cry_1 ));
    CascadeMux I__4263 (
            .O(N__23846),
            .I(N__23842));
    InMux I__4262 (
            .O(N__23845),
            .I(N__23839));
    InMux I__4261 (
            .O(N__23842),
            .I(N__23836));
    LocalMux I__4260 (
            .O(N__23839),
            .I(N__23833));
    LocalMux I__4259 (
            .O(N__23836),
            .I(\b2v_inst36.un2_count_1_axb_3 ));
    Odrv4 I__4258 (
            .O(N__23833),
            .I(\b2v_inst36.un2_count_1_axb_3 ));
    InMux I__4257 (
            .O(N__23828),
            .I(N__23822));
    InMux I__4256 (
            .O(N__23827),
            .I(N__23822));
    LocalMux I__4255 (
            .O(N__23822),
            .I(N__23819));
    Odrv4 I__4254 (
            .O(N__23819),
            .I(\b2v_inst36.un2_count_1_cry_2_THRU_CO ));
    InMux I__4253 (
            .O(N__23816),
            .I(\b2v_inst36.un2_count_1_cry_2 ));
    InMux I__4252 (
            .O(N__23813),
            .I(\b2v_inst36.un2_count_1_cry_3 ));
    CascadeMux I__4251 (
            .O(N__23810),
            .I(N__23806));
    CascadeMux I__4250 (
            .O(N__23809),
            .I(N__23803));
    InMux I__4249 (
            .O(N__23806),
            .I(N__23799));
    InMux I__4248 (
            .O(N__23803),
            .I(N__23796));
    InMux I__4247 (
            .O(N__23802),
            .I(N__23793));
    LocalMux I__4246 (
            .O(N__23799),
            .I(\b2v_inst36.countZ0Z_5 ));
    LocalMux I__4245 (
            .O(N__23796),
            .I(\b2v_inst36.countZ0Z_5 ));
    LocalMux I__4244 (
            .O(N__23793),
            .I(\b2v_inst36.countZ0Z_5 ));
    InMux I__4243 (
            .O(N__23786),
            .I(N__23783));
    LocalMux I__4242 (
            .O(N__23783),
            .I(N__23779));
    InMux I__4241 (
            .O(N__23782),
            .I(N__23776));
    Odrv4 I__4240 (
            .O(N__23779),
            .I(\b2v_inst36.un2_count_1_cry_4_THRU_CO ));
    LocalMux I__4239 (
            .O(N__23776),
            .I(\b2v_inst36.un2_count_1_cry_4_THRU_CO ));
    InMux I__4238 (
            .O(N__23771),
            .I(\b2v_inst36.un2_count_1_cry_4 ));
    InMux I__4237 (
            .O(N__23768),
            .I(\b2v_inst36.un2_count_1_cry_5 ));
    CascadeMux I__4236 (
            .O(N__23765),
            .I(\b2v_inst36.countZ0Z_2_cascade_ ));
    InMux I__4235 (
            .O(N__23762),
            .I(N__23759));
    LocalMux I__4234 (
            .O(N__23759),
            .I(\b2v_inst36.count_2_2 ));
    CascadeMux I__4233 (
            .O(N__23756),
            .I(\b2v_inst36.count_rst_7_cascade_ ));
    CascadeMux I__4232 (
            .O(N__23753),
            .I(\b2v_inst36.count_rst_9_cascade_ ));
    InMux I__4231 (
            .O(N__23750),
            .I(N__23747));
    LocalMux I__4230 (
            .O(N__23747),
            .I(\b2v_inst36.count_2_5 ));
    InMux I__4229 (
            .O(N__23744),
            .I(N__23738));
    InMux I__4228 (
            .O(N__23743),
            .I(N__23738));
    LocalMux I__4227 (
            .O(N__23738),
            .I(\b2v_inst36.count_2_7 ));
    InMux I__4226 (
            .O(N__23735),
            .I(N__23732));
    LocalMux I__4225 (
            .O(N__23732),
            .I(\b2v_inst36.count_rst_7 ));
    CascadeMux I__4224 (
            .O(N__23729),
            .I(\b2v_inst36.countZ0Z_5_cascade_ ));
    CascadeMux I__4223 (
            .O(N__23726),
            .I(\b2v_inst11.count_clkZ0Z_15_cascade_ ));
    InMux I__4222 (
            .O(N__23723),
            .I(N__23717));
    InMux I__4221 (
            .O(N__23722),
            .I(N__23717));
    LocalMux I__4220 (
            .O(N__23717),
            .I(\b2v_inst11.N_175 ));
    InMux I__4219 (
            .O(N__23714),
            .I(N__23711));
    LocalMux I__4218 (
            .O(N__23711),
            .I(\b2v_inst11.count_clk_0_14 ));
    CascadeMux I__4217 (
            .O(N__23708),
            .I(N__23705));
    InMux I__4216 (
            .O(N__23705),
            .I(N__23702));
    LocalMux I__4215 (
            .O(N__23702),
            .I(\b2v_inst11.count_clk_0_15 ));
    CascadeMux I__4214 (
            .O(N__23699),
            .I(\b2v_inst36.un2_count_1_axb_3_cascade_ ));
    InMux I__4213 (
            .O(N__23696),
            .I(N__23693));
    LocalMux I__4212 (
            .O(N__23693),
            .I(\b2v_inst36.count_rst_11 ));
    CascadeMux I__4211 (
            .O(N__23690),
            .I(\b2v_inst36.count_rst_11_cascade_ ));
    InMux I__4210 (
            .O(N__23687),
            .I(N__23681));
    InMux I__4209 (
            .O(N__23686),
            .I(N__23681));
    LocalMux I__4208 (
            .O(N__23681),
            .I(\b2v_inst36.count_2_3 ));
    CascadeMux I__4207 (
            .O(N__23678),
            .I(\b2v_inst36.count_rst_12_cascade_ ));
    CascadeMux I__4206 (
            .O(N__23675),
            .I(N__23672));
    InMux I__4205 (
            .O(N__23672),
            .I(N__23669));
    LocalMux I__4204 (
            .O(N__23669),
            .I(\b2v_inst11.count_clk_0_9 ));
    CascadeMux I__4203 (
            .O(N__23666),
            .I(\b2v_inst11.count_clkZ0Z_9_cascade_ ));
    InMux I__4202 (
            .O(N__23663),
            .I(N__23657));
    InMux I__4201 (
            .O(N__23662),
            .I(N__23657));
    LocalMux I__4200 (
            .O(N__23657),
            .I(\b2v_inst11.N_190 ));
    InMux I__4199 (
            .O(N__23654),
            .I(N__23651));
    LocalMux I__4198 (
            .O(N__23651),
            .I(\b2v_inst11.count_clk_0_5 ));
    CascadeMux I__4197 (
            .O(N__23648),
            .I(\b2v_inst11.count_clkZ0Z_5_cascade_ ));
    InMux I__4196 (
            .O(N__23645),
            .I(N__23642));
    LocalMux I__4195 (
            .O(N__23642),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2 ));
    CascadeMux I__4194 (
            .O(N__23639),
            .I(\b2v_inst11.count_clkZ0Z_1_cascade_ ));
    InMux I__4193 (
            .O(N__23636),
            .I(N__23633));
    LocalMux I__4192 (
            .O(N__23633),
            .I(\b2v_inst11.count_clk_0_1 ));
    InMux I__4191 (
            .O(N__23630),
            .I(N__23627));
    LocalMux I__4190 (
            .O(N__23627),
            .I(\b2v_inst11.count_clk_0_8 ));
    CascadeMux I__4189 (
            .O(N__23624),
            .I(\b2v_inst11.count_clkZ0Z_8_cascade_ ));
    CascadeMux I__4188 (
            .O(N__23621),
            .I(\b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ));
    CascadeMux I__4187 (
            .O(N__23618),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ));
    InMux I__4186 (
            .O(N__23615),
            .I(N__23612));
    LocalMux I__4185 (
            .O(N__23612),
            .I(\b2v_inst11.N_379 ));
    CascadeMux I__4184 (
            .O(N__23609),
            .I(\b2v_inst11.N_379_cascade_ ));
    CascadeMux I__4183 (
            .O(N__23606),
            .I(N__23602));
    InMux I__4182 (
            .O(N__23605),
            .I(N__23597));
    InMux I__4181 (
            .O(N__23602),
            .I(N__23597));
    LocalMux I__4180 (
            .O(N__23597),
            .I(\b2v_inst11.dutycycle_eena_13_0 ));
    CascadeMux I__4179 (
            .O(N__23594),
            .I(\b2v_inst11.N_200_i_cascade_ ));
    CascadeMux I__4178 (
            .O(N__23591),
            .I(\b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1_cascade_ ));
    InMux I__4177 (
            .O(N__23588),
            .I(N__23582));
    InMux I__4176 (
            .O(N__23587),
            .I(N__23582));
    LocalMux I__4175 (
            .O(N__23582),
            .I(N__23579));
    Span4Mux_v I__4174 (
            .O(N__23579),
            .I(N__23576));
    Odrv4 I__4173 (
            .O(N__23576),
            .I(\b2v_inst11.dutycycle_eena_3 ));
    InMux I__4172 (
            .O(N__23573),
            .I(N__23565));
    InMux I__4171 (
            .O(N__23572),
            .I(N__23558));
    InMux I__4170 (
            .O(N__23571),
            .I(N__23558));
    CascadeMux I__4169 (
            .O(N__23570),
            .I(N__23555));
    InMux I__4168 (
            .O(N__23569),
            .I(N__23550));
    CascadeMux I__4167 (
            .O(N__23568),
            .I(N__23547));
    LocalMux I__4166 (
            .O(N__23565),
            .I(N__23538));
    InMux I__4165 (
            .O(N__23564),
            .I(N__23533));
    InMux I__4164 (
            .O(N__23563),
            .I(N__23533));
    LocalMux I__4163 (
            .O(N__23558),
            .I(N__23528));
    InMux I__4162 (
            .O(N__23555),
            .I(N__23525));
    InMux I__4161 (
            .O(N__23554),
            .I(N__23520));
    InMux I__4160 (
            .O(N__23553),
            .I(N__23520));
    LocalMux I__4159 (
            .O(N__23550),
            .I(N__23517));
    InMux I__4158 (
            .O(N__23547),
            .I(N__23514));
    InMux I__4157 (
            .O(N__23546),
            .I(N__23511));
    InMux I__4156 (
            .O(N__23545),
            .I(N__23506));
    InMux I__4155 (
            .O(N__23544),
            .I(N__23506));
    InMux I__4154 (
            .O(N__23543),
            .I(N__23503));
    InMux I__4153 (
            .O(N__23542),
            .I(N__23498));
    InMux I__4152 (
            .O(N__23541),
            .I(N__23498));
    Span4Mux_v I__4151 (
            .O(N__23538),
            .I(N__23493));
    LocalMux I__4150 (
            .O(N__23533),
            .I(N__23493));
    InMux I__4149 (
            .O(N__23532),
            .I(N__23488));
    InMux I__4148 (
            .O(N__23531),
            .I(N__23488));
    Span4Mux_h I__4147 (
            .O(N__23528),
            .I(N__23485));
    LocalMux I__4146 (
            .O(N__23525),
            .I(N__23480));
    LocalMux I__4145 (
            .O(N__23520),
            .I(N__23480));
    Span4Mux_v I__4144 (
            .O(N__23517),
            .I(N__23475));
    LocalMux I__4143 (
            .O(N__23514),
            .I(N__23475));
    LocalMux I__4142 (
            .O(N__23511),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    LocalMux I__4141 (
            .O(N__23506),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    LocalMux I__4140 (
            .O(N__23503),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    LocalMux I__4139 (
            .O(N__23498),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    Odrv4 I__4138 (
            .O(N__23493),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    LocalMux I__4137 (
            .O(N__23488),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    Odrv4 I__4136 (
            .O(N__23485),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    Odrv4 I__4135 (
            .O(N__23480),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    Odrv4 I__4134 (
            .O(N__23475),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    InMux I__4133 (
            .O(N__23456),
            .I(N__23453));
    LocalMux I__4132 (
            .O(N__23453),
            .I(\b2v_inst11.un1_clk_100khz_32_and_i_0_c ));
    InMux I__4131 (
            .O(N__23450),
            .I(N__23444));
    InMux I__4130 (
            .O(N__23449),
            .I(N__23444));
    LocalMux I__4129 (
            .O(N__23444),
            .I(N__23441));
    Odrv4 I__4128 (
            .O(N__23441),
            .I(\b2v_inst11.un1_clk_100khz_40_and_i_0_c ));
    CascadeMux I__4127 (
            .O(N__23438),
            .I(N__23431));
    InMux I__4126 (
            .O(N__23437),
            .I(N__23426));
    InMux I__4125 (
            .O(N__23436),
            .I(N__23426));
    InMux I__4124 (
            .O(N__23435),
            .I(N__23419));
    InMux I__4123 (
            .O(N__23434),
            .I(N__23414));
    InMux I__4122 (
            .O(N__23431),
            .I(N__23414));
    LocalMux I__4121 (
            .O(N__23426),
            .I(N__23411));
    CascadeMux I__4120 (
            .O(N__23425),
            .I(N__23408));
    InMux I__4119 (
            .O(N__23424),
            .I(N__23405));
    CascadeMux I__4118 (
            .O(N__23423),
            .I(N__23402));
    InMux I__4117 (
            .O(N__23422),
            .I(N__23394));
    LocalMux I__4116 (
            .O(N__23419),
            .I(N__23389));
    LocalMux I__4115 (
            .O(N__23414),
            .I(N__23389));
    Span4Mux_h I__4114 (
            .O(N__23411),
            .I(N__23386));
    InMux I__4113 (
            .O(N__23408),
            .I(N__23383));
    LocalMux I__4112 (
            .O(N__23405),
            .I(N__23380));
    InMux I__4111 (
            .O(N__23402),
            .I(N__23377));
    InMux I__4110 (
            .O(N__23401),
            .I(N__23366));
    InMux I__4109 (
            .O(N__23400),
            .I(N__23366));
    InMux I__4108 (
            .O(N__23399),
            .I(N__23366));
    InMux I__4107 (
            .O(N__23398),
            .I(N__23366));
    InMux I__4106 (
            .O(N__23397),
            .I(N__23366));
    LocalMux I__4105 (
            .O(N__23394),
            .I(N__23363));
    Span4Mux_v I__4104 (
            .O(N__23389),
            .I(N__23360));
    Span4Mux_h I__4103 (
            .O(N__23386),
            .I(N__23355));
    LocalMux I__4102 (
            .O(N__23383),
            .I(N__23355));
    Odrv12 I__4101 (
            .O(N__23380),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__4100 (
            .O(N__23377),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__4099 (
            .O(N__23366),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__4098 (
            .O(N__23363),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__4097 (
            .O(N__23360),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__4096 (
            .O(N__23355),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    InMux I__4095 (
            .O(N__23342),
            .I(N__23339));
    LocalMux I__4094 (
            .O(N__23339),
            .I(\b2v_inst11.mult1_un145_sum ));
    CascadeMux I__4093 (
            .O(N__23336),
            .I(\b2v_inst11.mult1_un145_sum_cascade_ ));
    InMux I__4092 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__4091 (
            .O(N__23330),
            .I(N__23327));
    Span4Mux_s3_v I__4090 (
            .O(N__23327),
            .I(N__23324));
    Odrv4 I__4089 (
            .O(N__23324),
            .I(\b2v_inst11.mult1_un145_sum_i ));
    InMux I__4088 (
            .O(N__23321),
            .I(N__23318));
    LocalMux I__4087 (
            .O(N__23318),
            .I(N__23315));
    Odrv4 I__4086 (
            .O(N__23315),
            .I(\b2v_inst11.N_10 ));
    CascadeMux I__4085 (
            .O(N__23312),
            .I(\b2v_inst11.dutycycleZ0Z_12_cascade_ ));
    CascadeMux I__4084 (
            .O(N__23309),
            .I(N__23306));
    InMux I__4083 (
            .O(N__23306),
            .I(N__23302));
    InMux I__4082 (
            .O(N__23305),
            .I(N__23299));
    LocalMux I__4081 (
            .O(N__23302),
            .I(N__23296));
    LocalMux I__4080 (
            .O(N__23299),
            .I(N__23293));
    Span4Mux_v I__4079 (
            .O(N__23296),
            .I(N__23290));
    Span4Mux_h I__4078 (
            .O(N__23293),
            .I(N__23287));
    Odrv4 I__4077 (
            .O(N__23290),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_13 ));
    Odrv4 I__4076 (
            .O(N__23287),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_13 ));
    InMux I__4075 (
            .O(N__23282),
            .I(N__23279));
    LocalMux I__4074 (
            .O(N__23279),
            .I(N__23276));
    Odrv4 I__4073 (
            .O(N__23276),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_14 ));
    InMux I__4072 (
            .O(N__23273),
            .I(N__23270));
    LocalMux I__4071 (
            .O(N__23270),
            .I(N__23267));
    Odrv12 I__4070 (
            .O(N__23267),
            .I(\b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19 ));
    CascadeMux I__4069 (
            .O(N__23264),
            .I(\b2v_inst11.dutycycle_set_1_cascade_ ));
    CascadeMux I__4068 (
            .O(N__23261),
            .I(N__23258));
    InMux I__4067 (
            .O(N__23258),
            .I(N__23255));
    LocalMux I__4066 (
            .O(N__23255),
            .I(\b2v_inst11.N_300 ));
    CascadeMux I__4065 (
            .O(N__23252),
            .I(\b2v_inst11.N_300_0_cascade_ ));
    InMux I__4064 (
            .O(N__23249),
            .I(N__23246));
    LocalMux I__4063 (
            .O(N__23246),
            .I(N__23243));
    Span4Mux_v I__4062 (
            .O(N__23243),
            .I(N__23240));
    Odrv4 I__4061 (
            .O(N__23240),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29 ));
    InMux I__4060 (
            .O(N__23237),
            .I(N__23234));
    LocalMux I__4059 (
            .O(N__23234),
            .I(\b2v_inst11.dutycycle_set_0_0 ));
    CascadeMux I__4058 (
            .O(N__23231),
            .I(\b2v_inst11.dutycycle_set_0_0_cascade_ ));
    InMux I__4057 (
            .O(N__23228),
            .I(N__23222));
    InMux I__4056 (
            .O(N__23227),
            .I(N__23222));
    LocalMux I__4055 (
            .O(N__23222),
            .I(\b2v_inst11.dutycycle_0_6 ));
    InMux I__4054 (
            .O(N__23219),
            .I(N__23213));
    InMux I__4053 (
            .O(N__23218),
            .I(N__23213));
    LocalMux I__4052 (
            .O(N__23213),
            .I(\b2v_inst11.dutycycle_0_5 ));
    CascadeMux I__4051 (
            .O(N__23210),
            .I(N__23207));
    InMux I__4050 (
            .O(N__23207),
            .I(N__23204));
    LocalMux I__4049 (
            .O(N__23204),
            .I(\b2v_inst11.dutycycle_set_1 ));
    CascadeMux I__4048 (
            .O(N__23201),
            .I(\b2v_inst11.un1_clk_100khz_40_and_i_0_0_0_cascade_ ));
    InMux I__4047 (
            .O(N__23198),
            .I(N__23192));
    InMux I__4046 (
            .O(N__23197),
            .I(N__23192));
    LocalMux I__4045 (
            .O(N__23192),
            .I(N__23189));
    Odrv4 I__4044 (
            .O(N__23189),
            .I(\b2v_inst11.dutycycle_RNIT35D7Z0Z_4 ));
    CascadeMux I__4043 (
            .O(N__23186),
            .I(N__23183));
    InMux I__4042 (
            .O(N__23183),
            .I(N__23180));
    LocalMux I__4041 (
            .O(N__23180),
            .I(N__23177));
    Span4Mux_h I__4040 (
            .O(N__23177),
            .I(N__23174));
    Odrv4 I__4039 (
            .O(N__23174),
            .I(\b2v_inst11.N_155_N ));
    CascadeMux I__4038 (
            .O(N__23171),
            .I(\b2v_inst11.dutycycle_en_11_cascade_ ));
    CascadeMux I__4037 (
            .O(N__23168),
            .I(\b2v_inst11.N_158_N_cascade_ ));
    CascadeMux I__4036 (
            .O(N__23165),
            .I(N__23162));
    InMux I__4035 (
            .O(N__23162),
            .I(N__23159));
    LocalMux I__4034 (
            .O(N__23159),
            .I(\b2v_inst11.dutycycle_RNIT35D7Z0Z_15 ));
    InMux I__4033 (
            .O(N__23156),
            .I(N__23150));
    InMux I__4032 (
            .O(N__23155),
            .I(N__23150));
    LocalMux I__4031 (
            .O(N__23150),
            .I(N__23147));
    Odrv4 I__4030 (
            .O(N__23147),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ));
    CascadeMux I__4029 (
            .O(N__23144),
            .I(\b2v_inst11.dutycycle_RNIT35D7Z0Z_15_cascade_ ));
    InMux I__4028 (
            .O(N__23141),
            .I(N__23135));
    InMux I__4027 (
            .O(N__23140),
            .I(N__23135));
    LocalMux I__4026 (
            .O(N__23135),
            .I(N__23132));
    Odrv4 I__4025 (
            .O(N__23132),
            .I(\b2v_inst11.dutycycleZ0Z_15 ));
    InMux I__4024 (
            .O(N__23129),
            .I(N__23123));
    InMux I__4023 (
            .O(N__23128),
            .I(N__23123));
    LocalMux I__4022 (
            .O(N__23123),
            .I(\b2v_inst11.dutycycleZ0Z_14 ));
    CascadeMux I__4021 (
            .O(N__23120),
            .I(N__23117));
    InMux I__4020 (
            .O(N__23117),
            .I(N__23114));
    LocalMux I__4019 (
            .O(N__23114),
            .I(\b2v_inst11.dutycycle_en_11 ));
    InMux I__4018 (
            .O(N__23111),
            .I(N__23105));
    InMux I__4017 (
            .O(N__23110),
            .I(N__23105));
    LocalMux I__4016 (
            .O(N__23105),
            .I(N__23102));
    Odrv4 I__4015 (
            .O(N__23102),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ));
    CascadeMux I__4014 (
            .O(N__23099),
            .I(N__23096));
    InMux I__4013 (
            .O(N__23096),
            .I(N__23092));
    CascadeMux I__4012 (
            .O(N__23095),
            .I(N__23088));
    LocalMux I__4011 (
            .O(N__23092),
            .I(N__23083));
    InMux I__4010 (
            .O(N__23091),
            .I(N__23080));
    InMux I__4009 (
            .O(N__23088),
            .I(N__23077));
    InMux I__4008 (
            .O(N__23087),
            .I(N__23073));
    CascadeMux I__4007 (
            .O(N__23086),
            .I(N__23070));
    Span4Mux_v I__4006 (
            .O(N__23083),
            .I(N__23065));
    LocalMux I__4005 (
            .O(N__23080),
            .I(N__23065));
    LocalMux I__4004 (
            .O(N__23077),
            .I(N__23062));
    CascadeMux I__4003 (
            .O(N__23076),
            .I(N__23058));
    LocalMux I__4002 (
            .O(N__23073),
            .I(N__23054));
    InMux I__4001 (
            .O(N__23070),
            .I(N__23051));
    Span4Mux_v I__4000 (
            .O(N__23065),
            .I(N__23048));
    Span4Mux_v I__3999 (
            .O(N__23062),
            .I(N__23045));
    InMux I__3998 (
            .O(N__23061),
            .I(N__23040));
    InMux I__3997 (
            .O(N__23058),
            .I(N__23040));
    InMux I__3996 (
            .O(N__23057),
            .I(N__23037));
    Span4Mux_h I__3995 (
            .O(N__23054),
            .I(N__23032));
    LocalMux I__3994 (
            .O(N__23051),
            .I(N__23032));
    Odrv4 I__3993 (
            .O(N__23048),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__3992 (
            .O(N__23045),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    LocalMux I__3991 (
            .O(N__23040),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    LocalMux I__3990 (
            .O(N__23037),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__3989 (
            .O(N__23032),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    InMux I__3988 (
            .O(N__23021),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11_cZ0 ));
    InMux I__3987 (
            .O(N__23018),
            .I(N__23012));
    InMux I__3986 (
            .O(N__23017),
            .I(N__23012));
    LocalMux I__3985 (
            .O(N__23012),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ));
    InMux I__3984 (
            .O(N__23009),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_cZ0 ));
    InMux I__3983 (
            .O(N__23006),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_cZ0 ));
    InMux I__3982 (
            .O(N__23003),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14 ));
    CascadeMux I__3981 (
            .O(N__23000),
            .I(\b2v_inst11.un1_clk_100khz_43_and_i_0_0_0_cascade_ ));
    CascadeMux I__3980 (
            .O(N__22997),
            .I(\b2v_inst11.dutycycleZ0Z_3_cascade_ ));
    CascadeMux I__3979 (
            .O(N__22994),
            .I(N__22991));
    InMux I__3978 (
            .O(N__22991),
            .I(N__22988));
    LocalMux I__3977 (
            .O(N__22988),
            .I(\b2v_inst11.un1_clk_100khz_43_and_i_0_d_0 ));
    InMux I__3976 (
            .O(N__22985),
            .I(N__22982));
    LocalMux I__3975 (
            .O(N__22982),
            .I(N__22979));
    Odrv4 I__3974 (
            .O(N__22979),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ));
    InMux I__3973 (
            .O(N__22976),
            .I(N__22973));
    LocalMux I__3972 (
            .O(N__22973),
            .I(\b2v_inst11.dutycycle_e_1_3 ));
    InMux I__3971 (
            .O(N__22970),
            .I(N__22967));
    LocalMux I__3970 (
            .O(N__22967),
            .I(\b2v_inst11.un1_clk_100khz_43_and_i_0_0_0 ));
    CascadeMux I__3969 (
            .O(N__22964),
            .I(\b2v_inst11.dutycycle_e_1_3_cascade_ ));
    CascadeMux I__3968 (
            .O(N__22961),
            .I(N__22958));
    InMux I__3967 (
            .O(N__22958),
            .I(N__22953));
    InMux I__3966 (
            .O(N__22957),
            .I(N__22948));
    InMux I__3965 (
            .O(N__22956),
            .I(N__22948));
    LocalMux I__3964 (
            .O(N__22953),
            .I(\b2v_inst11.dutycycle_0_3 ));
    LocalMux I__3963 (
            .O(N__22948),
            .I(\b2v_inst11.dutycycle_0_3 ));
    CascadeMux I__3962 (
            .O(N__22943),
            .I(N__22940));
    InMux I__3961 (
            .O(N__22940),
            .I(N__22934));
    InMux I__3960 (
            .O(N__22939),
            .I(N__22934));
    LocalMux I__3959 (
            .O(N__22934),
            .I(N__22931));
    Odrv4 I__3958 (
            .O(N__22931),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ));
    InMux I__3957 (
            .O(N__22928),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3 ));
    InMux I__3956 (
            .O(N__22925),
            .I(\b2v_inst11.un1_dutycycle_94_cry_4 ));
    InMux I__3955 (
            .O(N__22922),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ));
    CascadeMux I__3954 (
            .O(N__22919),
            .I(N__22909));
    InMux I__3953 (
            .O(N__22918),
            .I(N__22905));
    InMux I__3952 (
            .O(N__22917),
            .I(N__22900));
    InMux I__3951 (
            .O(N__22916),
            .I(N__22900));
    InMux I__3950 (
            .O(N__22915),
            .I(N__22895));
    InMux I__3949 (
            .O(N__22914),
            .I(N__22895));
    InMux I__3948 (
            .O(N__22913),
            .I(N__22892));
    InMux I__3947 (
            .O(N__22912),
            .I(N__22889));
    InMux I__3946 (
            .O(N__22909),
            .I(N__22886));
    InMux I__3945 (
            .O(N__22908),
            .I(N__22883));
    LocalMux I__3944 (
            .O(N__22905),
            .I(N__22878));
    LocalMux I__3943 (
            .O(N__22900),
            .I(N__22878));
    LocalMux I__3942 (
            .O(N__22895),
            .I(N__22874));
    LocalMux I__3941 (
            .O(N__22892),
            .I(N__22871));
    LocalMux I__3940 (
            .O(N__22889),
            .I(N__22866));
    LocalMux I__3939 (
            .O(N__22886),
            .I(N__22866));
    LocalMux I__3938 (
            .O(N__22883),
            .I(N__22861));
    Span4Mux_v I__3937 (
            .O(N__22878),
            .I(N__22861));
    InMux I__3936 (
            .O(N__22877),
            .I(N__22858));
    Span4Mux_h I__3935 (
            .O(N__22874),
            .I(N__22853));
    Span4Mux_v I__3934 (
            .O(N__22871),
            .I(N__22853));
    Span4Mux_h I__3933 (
            .O(N__22866),
            .I(N__22850));
    Odrv4 I__3932 (
            .O(N__22861),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    LocalMux I__3931 (
            .O(N__22858),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    Odrv4 I__3930 (
            .O(N__22853),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    Odrv4 I__3929 (
            .O(N__22850),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    CascadeMux I__3928 (
            .O(N__22841),
            .I(N__22837));
    CascadeMux I__3927 (
            .O(N__22840),
            .I(N__22834));
    InMux I__3926 (
            .O(N__22837),
            .I(N__22831));
    InMux I__3925 (
            .O(N__22834),
            .I(N__22828));
    LocalMux I__3924 (
            .O(N__22831),
            .I(N__22823));
    LocalMux I__3923 (
            .O(N__22828),
            .I(N__22823));
    Span4Mux_h I__3922 (
            .O(N__22823),
            .I(N__22820));
    Odrv4 I__3921 (
            .O(N__22820),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ));
    InMux I__3920 (
            .O(N__22817),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ));
    CascadeMux I__3919 (
            .O(N__22814),
            .I(N__22810));
    InMux I__3918 (
            .O(N__22813),
            .I(N__22805));
    InMux I__3917 (
            .O(N__22810),
            .I(N__22805));
    LocalMux I__3916 (
            .O(N__22805),
            .I(N__22802));
    Odrv4 I__3915 (
            .O(N__22802),
            .I(\b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9JZ0Z1 ));
    InMux I__3914 (
            .O(N__22799),
            .I(bfn_7_8_0_));
    CascadeMux I__3913 (
            .O(N__22796),
            .I(N__22792));
    CascadeMux I__3912 (
            .O(N__22795),
            .I(N__22785));
    InMux I__3911 (
            .O(N__22792),
            .I(N__22782));
    CascadeMux I__3910 (
            .O(N__22791),
            .I(N__22765));
    CascadeMux I__3909 (
            .O(N__22790),
            .I(N__22762));
    InMux I__3908 (
            .O(N__22789),
            .I(N__22753));
    InMux I__3907 (
            .O(N__22788),
            .I(N__22753));
    InMux I__3906 (
            .O(N__22785),
            .I(N__22753));
    LocalMux I__3905 (
            .O(N__22782),
            .I(N__22750));
    InMux I__3904 (
            .O(N__22781),
            .I(N__22747));
    InMux I__3903 (
            .O(N__22780),
            .I(N__22742));
    InMux I__3902 (
            .O(N__22779),
            .I(N__22742));
    InMux I__3901 (
            .O(N__22778),
            .I(N__22735));
    InMux I__3900 (
            .O(N__22777),
            .I(N__22735));
    InMux I__3899 (
            .O(N__22776),
            .I(N__22735));
    InMux I__3898 (
            .O(N__22775),
            .I(N__22732));
    InMux I__3897 (
            .O(N__22774),
            .I(N__22723));
    InMux I__3896 (
            .O(N__22773),
            .I(N__22723));
    InMux I__3895 (
            .O(N__22772),
            .I(N__22723));
    InMux I__3894 (
            .O(N__22771),
            .I(N__22723));
    InMux I__3893 (
            .O(N__22770),
            .I(N__22716));
    InMux I__3892 (
            .O(N__22769),
            .I(N__22716));
    InMux I__3891 (
            .O(N__22768),
            .I(N__22716));
    InMux I__3890 (
            .O(N__22765),
            .I(N__22707));
    InMux I__3889 (
            .O(N__22762),
            .I(N__22707));
    InMux I__3888 (
            .O(N__22761),
            .I(N__22707));
    InMux I__3887 (
            .O(N__22760),
            .I(N__22707));
    LocalMux I__3886 (
            .O(N__22753),
            .I(N__22702));
    Span4Mux_h I__3885 (
            .O(N__22750),
            .I(N__22702));
    LocalMux I__3884 (
            .O(N__22747),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3883 (
            .O(N__22742),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3882 (
            .O(N__22735),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3881 (
            .O(N__22732),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3880 (
            .O(N__22723),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3879 (
            .O(N__22716),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3878 (
            .O(N__22707),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__3877 (
            .O(N__22702),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    InMux I__3876 (
            .O(N__22685),
            .I(N__22679));
    InMux I__3875 (
            .O(N__22684),
            .I(N__22679));
    LocalMux I__3874 (
            .O(N__22679),
            .I(N__22676));
    Span4Mux_h I__3873 (
            .O(N__22676),
            .I(N__22673));
    Odrv4 I__3872 (
            .O(N__22673),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJZ0Z1 ));
    InMux I__3871 (
            .O(N__22670),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ));
    CascadeMux I__3870 (
            .O(N__22667),
            .I(N__22662));
    CascadeMux I__3869 (
            .O(N__22666),
            .I(N__22654));
    CascadeMux I__3868 (
            .O(N__22665),
            .I(N__22651));
    InMux I__3867 (
            .O(N__22662),
            .I(N__22647));
    InMux I__3866 (
            .O(N__22661),
            .I(N__22643));
    CascadeMux I__3865 (
            .O(N__22660),
            .I(N__22638));
    CascadeMux I__3864 (
            .O(N__22659),
            .I(N__22632));
    CascadeMux I__3863 (
            .O(N__22658),
            .I(N__22628));
    CascadeMux I__3862 (
            .O(N__22657),
            .I(N__22625));
    InMux I__3861 (
            .O(N__22654),
            .I(N__22620));
    InMux I__3860 (
            .O(N__22651),
            .I(N__22620));
    InMux I__3859 (
            .O(N__22650),
            .I(N__22617));
    LocalMux I__3858 (
            .O(N__22647),
            .I(N__22614));
    InMux I__3857 (
            .O(N__22646),
            .I(N__22611));
    LocalMux I__3856 (
            .O(N__22643),
            .I(N__22608));
    InMux I__3855 (
            .O(N__22642),
            .I(N__22603));
    InMux I__3854 (
            .O(N__22641),
            .I(N__22603));
    InMux I__3853 (
            .O(N__22638),
            .I(N__22596));
    InMux I__3852 (
            .O(N__22637),
            .I(N__22596));
    InMux I__3851 (
            .O(N__22636),
            .I(N__22596));
    InMux I__3850 (
            .O(N__22635),
            .I(N__22591));
    InMux I__3849 (
            .O(N__22632),
            .I(N__22591));
    InMux I__3848 (
            .O(N__22631),
            .I(N__22588));
    InMux I__3847 (
            .O(N__22628),
            .I(N__22583));
    InMux I__3846 (
            .O(N__22625),
            .I(N__22583));
    LocalMux I__3845 (
            .O(N__22620),
            .I(N__22578));
    LocalMux I__3844 (
            .O(N__22617),
            .I(N__22578));
    Span4Mux_v I__3843 (
            .O(N__22614),
            .I(N__22575));
    LocalMux I__3842 (
            .O(N__22611),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__3841 (
            .O(N__22608),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__3840 (
            .O(N__22603),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__3839 (
            .O(N__22596),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__3838 (
            .O(N__22591),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__3837 (
            .O(N__22588),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__3836 (
            .O(N__22583),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__3835 (
            .O(N__22578),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__3834 (
            .O(N__22575),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    InMux I__3833 (
            .O(N__22556),
            .I(N__22550));
    InMux I__3832 (
            .O(N__22555),
            .I(N__22550));
    LocalMux I__3831 (
            .O(N__22550),
            .I(N__22547));
    Span4Mux_v I__3830 (
            .O(N__22547),
            .I(N__22544));
    Odrv4 I__3829 (
            .O(N__22544),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJZ0Z1 ));
    InMux I__3828 (
            .O(N__22541),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9 ));
    InMux I__3827 (
            .O(N__22538),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10 ));
    InMux I__3826 (
            .O(N__22535),
            .I(N__22532));
    LocalMux I__3825 (
            .O(N__22532),
            .I(N__22529));
    Span4Mux_v I__3824 (
            .O(N__22529),
            .I(N__22526));
    Odrv4 I__3823 (
            .O(N__22526),
            .I(\b2v_inst5.un2_count_1_axb_11 ));
    InMux I__3822 (
            .O(N__22523),
            .I(N__22514));
    InMux I__3821 (
            .O(N__22522),
            .I(N__22514));
    InMux I__3820 (
            .O(N__22521),
            .I(N__22514));
    LocalMux I__3819 (
            .O(N__22514),
            .I(N__22511));
    Odrv4 I__3818 (
            .O(N__22511),
            .I(\b2v_inst5.count_rst_3 ));
    InMux I__3817 (
            .O(N__22508),
            .I(\b2v_inst5.un2_count_1_cry_10 ));
    InMux I__3816 (
            .O(N__22505),
            .I(N__22499));
    InMux I__3815 (
            .O(N__22504),
            .I(N__22499));
    LocalMux I__3814 (
            .O(N__22499),
            .I(N__22496));
    Odrv4 I__3813 (
            .O(N__22496),
            .I(\b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2 ));
    InMux I__3812 (
            .O(N__22493),
            .I(\b2v_inst5.un2_count_1_cry_11 ));
    InMux I__3811 (
            .O(N__22490),
            .I(\b2v_inst5.un2_count_1_cry_12 ));
    InMux I__3810 (
            .O(N__22487),
            .I(\b2v_inst5.un2_count_1_cry_13 ));
    InMux I__3809 (
            .O(N__22484),
            .I(\b2v_inst5.un2_count_1_cry_14 ));
    InMux I__3808 (
            .O(N__22481),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ));
    InMux I__3807 (
            .O(N__22478),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ));
    InMux I__3806 (
            .O(N__22475),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2 ));
    InMux I__3805 (
            .O(N__22472),
            .I(\b2v_inst5.un2_count_1_cry_1 ));
    InMux I__3804 (
            .O(N__22469),
            .I(\b2v_inst5.un2_count_1_cry_2 ));
    InMux I__3803 (
            .O(N__22466),
            .I(\b2v_inst5.un2_count_1_cry_3 ));
    InMux I__3802 (
            .O(N__22463),
            .I(\b2v_inst5.un2_count_1_cry_4 ));
    InMux I__3801 (
            .O(N__22460),
            .I(N__22454));
    InMux I__3800 (
            .O(N__22459),
            .I(N__22454));
    LocalMux I__3799 (
            .O(N__22454),
            .I(N__22451));
    Span4Mux_v I__3798 (
            .O(N__22451),
            .I(N__22448));
    Odrv4 I__3797 (
            .O(N__22448),
            .I(\b2v_inst5.count_rst_8 ));
    InMux I__3796 (
            .O(N__22445),
            .I(\b2v_inst5.un2_count_1_cry_5 ));
    InMux I__3795 (
            .O(N__22442),
            .I(N__22439));
    LocalMux I__3794 (
            .O(N__22439),
            .I(N__22436));
    Odrv12 I__3793 (
            .O(N__22436),
            .I(\b2v_inst5.countZ0Z_7 ));
    InMux I__3792 (
            .O(N__22433),
            .I(N__22427));
    InMux I__3791 (
            .O(N__22432),
            .I(N__22427));
    LocalMux I__3790 (
            .O(N__22427),
            .I(N__22424));
    Odrv4 I__3789 (
            .O(N__22424),
            .I(\b2v_inst5.count_rst_7 ));
    InMux I__3788 (
            .O(N__22421),
            .I(\b2v_inst5.un2_count_1_cry_6 ));
    InMux I__3787 (
            .O(N__22418),
            .I(bfn_7_6_0_));
    InMux I__3786 (
            .O(N__22415),
            .I(\b2v_inst5.un2_count_1_cry_8 ));
    InMux I__3785 (
            .O(N__22412),
            .I(\b2v_inst5.un2_count_1_cry_9 ));
    InMux I__3784 (
            .O(N__22409),
            .I(N__22406));
    LocalMux I__3783 (
            .O(N__22406),
            .I(N__22403));
    Odrv4 I__3782 (
            .O(N__22403),
            .I(\b2v_inst20.counter_1_cry_5_THRU_CO ));
    InMux I__3781 (
            .O(N__22400),
            .I(N__22396));
    CascadeMux I__3780 (
            .O(N__22399),
            .I(N__22392));
    LocalMux I__3779 (
            .O(N__22396),
            .I(N__22389));
    InMux I__3778 (
            .O(N__22395),
            .I(N__22384));
    InMux I__3777 (
            .O(N__22392),
            .I(N__22384));
    Odrv4 I__3776 (
            .O(N__22389),
            .I(\b2v_inst20.counterZ0Z_6 ));
    LocalMux I__3775 (
            .O(N__22384),
            .I(\b2v_inst20.counterZ0Z_6 ));
    InMux I__3774 (
            .O(N__22379),
            .I(N__22375));
    CascadeMux I__3773 (
            .O(N__22378),
            .I(N__22372));
    LocalMux I__3772 (
            .O(N__22375),
            .I(N__22368));
    InMux I__3771 (
            .O(N__22372),
            .I(N__22363));
    InMux I__3770 (
            .O(N__22371),
            .I(N__22363));
    Odrv4 I__3769 (
            .O(N__22368),
            .I(\b2v_inst20.counterZ0Z_1 ));
    LocalMux I__3768 (
            .O(N__22363),
            .I(\b2v_inst20.counterZ0Z_1 ));
    CascadeMux I__3767 (
            .O(N__22358),
            .I(N__22355));
    InMux I__3766 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__3765 (
            .O(N__22352),
            .I(N__22346));
    InMux I__3764 (
            .O(N__22351),
            .I(N__22339));
    InMux I__3763 (
            .O(N__22350),
            .I(N__22339));
    InMux I__3762 (
            .O(N__22349),
            .I(N__22339));
    Odrv4 I__3761 (
            .O(N__22346),
            .I(\b2v_inst20.counterZ0Z_0 ));
    LocalMux I__3760 (
            .O(N__22339),
            .I(\b2v_inst20.counterZ0Z_0 ));
    CascadeMux I__3759 (
            .O(N__22334),
            .I(N__22331));
    InMux I__3758 (
            .O(N__22331),
            .I(N__22328));
    LocalMux I__3757 (
            .O(N__22328),
            .I(N__22325));
    Odrv4 I__3756 (
            .O(N__22325),
            .I(\b2v_inst20.un4_counter_0_and ));
    InMux I__3755 (
            .O(N__22322),
            .I(N__22319));
    LocalMux I__3754 (
            .O(N__22319),
            .I(N__22316));
    Span4Mux_h I__3753 (
            .O(N__22316),
            .I(N__22313));
    Odrv4 I__3752 (
            .O(N__22313),
            .I(\b2v_inst20.counter_1_cry_4_THRU_CO ));
    InMux I__3751 (
            .O(N__22310),
            .I(N__22307));
    LocalMux I__3750 (
            .O(N__22307),
            .I(N__22302));
    InMux I__3749 (
            .O(N__22306),
            .I(N__22297));
    InMux I__3748 (
            .O(N__22305),
            .I(N__22297));
    Odrv4 I__3747 (
            .O(N__22302),
            .I(\b2v_inst20.counterZ0Z_5 ));
    LocalMux I__3746 (
            .O(N__22297),
            .I(\b2v_inst20.counterZ0Z_5 ));
    InMux I__3745 (
            .O(N__22292),
            .I(N__22289));
    LocalMux I__3744 (
            .O(N__22289),
            .I(N__22286));
    Odrv4 I__3743 (
            .O(N__22286),
            .I(\b2v_inst20.counter_1_cry_3_THRU_CO ));
    InMux I__3742 (
            .O(N__22283),
            .I(N__22279));
    CascadeMux I__3741 (
            .O(N__22282),
            .I(N__22275));
    LocalMux I__3740 (
            .O(N__22279),
            .I(N__22272));
    InMux I__3739 (
            .O(N__22278),
            .I(N__22267));
    InMux I__3738 (
            .O(N__22275),
            .I(N__22267));
    Odrv4 I__3737 (
            .O(N__22272),
            .I(\b2v_inst20.counterZ0Z_4 ));
    LocalMux I__3736 (
            .O(N__22267),
            .I(\b2v_inst20.counterZ0Z_4 ));
    InMux I__3735 (
            .O(N__22262),
            .I(\b2v_inst5.un2_count_1_cry_0 ));
    InMux I__3734 (
            .O(N__22259),
            .I(N__22256));
    LocalMux I__3733 (
            .O(N__22256),
            .I(\b2v_inst5.count_1_7 ));
    InMux I__3732 (
            .O(N__22253),
            .I(N__22247));
    InMux I__3731 (
            .O(N__22252),
            .I(N__22247));
    LocalMux I__3730 (
            .O(N__22247),
            .I(\b2v_inst5.count_1_11 ));
    CascadeMux I__3729 (
            .O(N__22244),
            .I(\b2v_inst5.countZ0Z_7_cascade_ ));
    InMux I__3728 (
            .O(N__22241),
            .I(N__22238));
    LocalMux I__3727 (
            .O(N__22238),
            .I(\b2v_inst5.count_1_12 ));
    InMux I__3726 (
            .O(N__22235),
            .I(N__22231));
    InMux I__3725 (
            .O(N__22234),
            .I(N__22228));
    LocalMux I__3724 (
            .O(N__22231),
            .I(N__22225));
    LocalMux I__3723 (
            .O(N__22228),
            .I(\b2v_inst20.counterZ0Z_7 ));
    Odrv4 I__3722 (
            .O(N__22225),
            .I(\b2v_inst20.counterZ0Z_7 ));
    CascadeMux I__3721 (
            .O(N__22220),
            .I(N__22217));
    InMux I__3720 (
            .O(N__22217),
            .I(N__22214));
    LocalMux I__3719 (
            .O(N__22214),
            .I(N__22211));
    Odrv12 I__3718 (
            .O(N__22211),
            .I(\b2v_inst20.un4_counter_1_and ));
    InMux I__3717 (
            .O(N__22208),
            .I(N__22205));
    LocalMux I__3716 (
            .O(N__22205),
            .I(\b2v_inst36.count_2_15 ));
    InMux I__3715 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__3714 (
            .O(N__22199),
            .I(\b2v_inst36.count_2_13 ));
    InMux I__3713 (
            .O(N__22196),
            .I(N__22193));
    LocalMux I__3712 (
            .O(N__22193),
            .I(\b2v_inst36.count_2_14 ));
    CascadeMux I__3711 (
            .O(N__22190),
            .I(N__22187));
    InMux I__3710 (
            .O(N__22187),
            .I(N__22182));
    InMux I__3709 (
            .O(N__22186),
            .I(N__22177));
    InMux I__3708 (
            .O(N__22185),
            .I(N__22177));
    LocalMux I__3707 (
            .O(N__22182),
            .I(\b2v_inst36.count_i_0 ));
    LocalMux I__3706 (
            .O(N__22177),
            .I(\b2v_inst36.count_i_0 ));
    InMux I__3705 (
            .O(N__22172),
            .I(N__22169));
    LocalMux I__3704 (
            .O(N__22169),
            .I(\b2v_inst11.mult1_un145_sum_cry_6_s ));
    CascadeMux I__3703 (
            .O(N__22166),
            .I(N__22162));
    CascadeMux I__3702 (
            .O(N__22165),
            .I(N__22158));
    InMux I__3701 (
            .O(N__22162),
            .I(N__22151));
    InMux I__3700 (
            .O(N__22161),
            .I(N__22151));
    InMux I__3699 (
            .O(N__22158),
            .I(N__22151));
    LocalMux I__3698 (
            .O(N__22151),
            .I(\b2v_inst11.mult1_un145_sum_i_0_8 ));
    CascadeMux I__3697 (
            .O(N__22148),
            .I(N__22145));
    InMux I__3696 (
            .O(N__22145),
            .I(N__22142));
    LocalMux I__3695 (
            .O(N__22142),
            .I(\b2v_inst11.mult1_un159_sum_axb_7 ));
    InMux I__3694 (
            .O(N__22139),
            .I(\b2v_inst11.mult1_un152_sum_cry_6 ));
    CascadeMux I__3693 (
            .O(N__22136),
            .I(N__22133));
    InMux I__3692 (
            .O(N__22133),
            .I(N__22130));
    LocalMux I__3691 (
            .O(N__22130),
            .I(\b2v_inst11.mult1_un152_sum_axb_8 ));
    InMux I__3690 (
            .O(N__22127),
            .I(\b2v_inst11.mult1_un152_sum_cry_7 ));
    InMux I__3689 (
            .O(N__22124),
            .I(N__22121));
    LocalMux I__3688 (
            .O(N__22121),
            .I(N__22117));
    CascadeMux I__3687 (
            .O(N__22120),
            .I(N__22113));
    Span4Mux_v I__3686 (
            .O(N__22117),
            .I(N__22109));
    InMux I__3685 (
            .O(N__22116),
            .I(N__22104));
    InMux I__3684 (
            .O(N__22113),
            .I(N__22104));
    InMux I__3683 (
            .O(N__22112),
            .I(N__22101));
    Odrv4 I__3682 (
            .O(N__22109),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    LocalMux I__3681 (
            .O(N__22104),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    LocalMux I__3680 (
            .O(N__22101),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    CascadeMux I__3679 (
            .O(N__22094),
            .I(\b2v_inst11.mult1_un152_sum_s_8_cascade_ ));
    CascadeMux I__3678 (
            .O(N__22091),
            .I(N__22087));
    CascadeMux I__3677 (
            .O(N__22090),
            .I(N__22083));
    InMux I__3676 (
            .O(N__22087),
            .I(N__22076));
    InMux I__3675 (
            .O(N__22086),
            .I(N__22076));
    InMux I__3674 (
            .O(N__22083),
            .I(N__22076));
    LocalMux I__3673 (
            .O(N__22076),
            .I(\b2v_inst11.mult1_un152_sum_i_0_8 ));
    CascadeMux I__3672 (
            .O(N__22073),
            .I(\b2v_inst36.count_rst_3_cascade_ ));
    CascadeMux I__3671 (
            .O(N__22070),
            .I(\b2v_inst36.countZ0Z_11_cascade_ ));
    InMux I__3670 (
            .O(N__22067),
            .I(N__22064));
    LocalMux I__3669 (
            .O(N__22064),
            .I(\b2v_inst36.count_2_11 ));
    InMux I__3668 (
            .O(N__22061),
            .I(N__22055));
    InMux I__3667 (
            .O(N__22060),
            .I(N__22055));
    LocalMux I__3666 (
            .O(N__22055),
            .I(\b2v_inst36.count_2_1 ));
    InMux I__3665 (
            .O(N__22052),
            .I(N__22049));
    LocalMux I__3664 (
            .O(N__22049),
            .I(\b2v_inst11.mult1_un138_sum_cry_6_s ));
    CascadeMux I__3663 (
            .O(N__22046),
            .I(N__22042));
    CascadeMux I__3662 (
            .O(N__22045),
            .I(N__22038));
    InMux I__3661 (
            .O(N__22042),
            .I(N__22031));
    InMux I__3660 (
            .O(N__22041),
            .I(N__22031));
    InMux I__3659 (
            .O(N__22038),
            .I(N__22031));
    LocalMux I__3658 (
            .O(N__22031),
            .I(\b2v_inst11.mult1_un138_sum_i_0_8 ));
    InMux I__3657 (
            .O(N__22028),
            .I(\b2v_inst11.mult1_un145_sum_cry_6 ));
    CascadeMux I__3656 (
            .O(N__22025),
            .I(N__22022));
    InMux I__3655 (
            .O(N__22022),
            .I(N__22019));
    LocalMux I__3654 (
            .O(N__22019),
            .I(\b2v_inst11.mult1_un145_sum_axb_8 ));
    InMux I__3653 (
            .O(N__22016),
            .I(\b2v_inst11.mult1_un145_sum_cry_7 ));
    CascadeMux I__3652 (
            .O(N__22013),
            .I(\b2v_inst11.mult1_un145_sum_s_8_cascade_ ));
    CascadeMux I__3651 (
            .O(N__22010),
            .I(N__22007));
    InMux I__3650 (
            .O(N__22007),
            .I(N__22004));
    LocalMux I__3649 (
            .O(N__22004),
            .I(\b2v_inst11.mult1_un152_sum_cry_3_s ));
    InMux I__3648 (
            .O(N__22001),
            .I(\b2v_inst11.mult1_un152_sum_cry_2 ));
    CascadeMux I__3647 (
            .O(N__21998),
            .I(N__21995));
    InMux I__3646 (
            .O(N__21995),
            .I(N__21992));
    LocalMux I__3645 (
            .O(N__21992),
            .I(\b2v_inst11.mult1_un145_sum_cry_3_s ));
    InMux I__3644 (
            .O(N__21989),
            .I(N__21986));
    LocalMux I__3643 (
            .O(N__21986),
            .I(\b2v_inst11.mult1_un152_sum_cry_4_s ));
    InMux I__3642 (
            .O(N__21983),
            .I(\b2v_inst11.mult1_un152_sum_cry_3 ));
    InMux I__3641 (
            .O(N__21980),
            .I(N__21977));
    LocalMux I__3640 (
            .O(N__21977),
            .I(\b2v_inst11.mult1_un145_sum_cry_4_s ));
    CascadeMux I__3639 (
            .O(N__21974),
            .I(N__21971));
    InMux I__3638 (
            .O(N__21971),
            .I(N__21968));
    LocalMux I__3637 (
            .O(N__21968),
            .I(\b2v_inst11.mult1_un152_sum_cry_5_s ));
    InMux I__3636 (
            .O(N__21965),
            .I(\b2v_inst11.mult1_un152_sum_cry_4 ));
    CascadeMux I__3635 (
            .O(N__21962),
            .I(N__21959));
    InMux I__3634 (
            .O(N__21959),
            .I(N__21955));
    CascadeMux I__3633 (
            .O(N__21958),
            .I(N__21951));
    LocalMux I__3632 (
            .O(N__21955),
            .I(N__21947));
    InMux I__3631 (
            .O(N__21954),
            .I(N__21942));
    InMux I__3630 (
            .O(N__21951),
            .I(N__21942));
    InMux I__3629 (
            .O(N__21950),
            .I(N__21939));
    Odrv4 I__3628 (
            .O(N__21947),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    LocalMux I__3627 (
            .O(N__21942),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    LocalMux I__3626 (
            .O(N__21939),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    CascadeMux I__3625 (
            .O(N__21932),
            .I(N__21929));
    InMux I__3624 (
            .O(N__21929),
            .I(N__21926));
    LocalMux I__3623 (
            .O(N__21926),
            .I(\b2v_inst11.mult1_un145_sum_cry_5_s ));
    InMux I__3622 (
            .O(N__21923),
            .I(N__21920));
    LocalMux I__3621 (
            .O(N__21920),
            .I(\b2v_inst11.mult1_un152_sum_cry_6_s ));
    InMux I__3620 (
            .O(N__21917),
            .I(\b2v_inst11.mult1_un152_sum_cry_5 ));
    InMux I__3619 (
            .O(N__21914),
            .I(\b2v_inst11.mult1_un138_sum_cry_5_c ));
    InMux I__3618 (
            .O(N__21911),
            .I(N__21908));
    LocalMux I__3617 (
            .O(N__21908),
            .I(\b2v_inst11.mult1_un131_sum_cry_6_s ));
    CascadeMux I__3616 (
            .O(N__21905),
            .I(N__21901));
    CascadeMux I__3615 (
            .O(N__21904),
            .I(N__21897));
    InMux I__3614 (
            .O(N__21901),
            .I(N__21890));
    InMux I__3613 (
            .O(N__21900),
            .I(N__21890));
    InMux I__3612 (
            .O(N__21897),
            .I(N__21890));
    LocalMux I__3611 (
            .O(N__21890),
            .I(\b2v_inst11.mult1_un131_sum_i_0_8 ));
    InMux I__3610 (
            .O(N__21887),
            .I(\b2v_inst11.mult1_un138_sum_cry_6_c ));
    CascadeMux I__3609 (
            .O(N__21884),
            .I(N__21881));
    InMux I__3608 (
            .O(N__21881),
            .I(N__21878));
    LocalMux I__3607 (
            .O(N__21878),
            .I(\b2v_inst11.mult1_un138_sum_axb_8 ));
    InMux I__3606 (
            .O(N__21875),
            .I(\b2v_inst11.mult1_un138_sum_cry_7 ));
    CascadeMux I__3605 (
            .O(N__21872),
            .I(\b2v_inst11.mult1_un138_sum_s_8_cascade_ ));
    InMux I__3604 (
            .O(N__21869),
            .I(N__21866));
    LocalMux I__3603 (
            .O(N__21866),
            .I(N__21863));
    Odrv12 I__3602 (
            .O(N__21863),
            .I(\b2v_inst11.mult1_un138_sum_i ));
    InMux I__3601 (
            .O(N__21860),
            .I(\b2v_inst11.mult1_un145_sum_cry_2 ));
    CascadeMux I__3600 (
            .O(N__21857),
            .I(N__21854));
    InMux I__3599 (
            .O(N__21854),
            .I(N__21851));
    LocalMux I__3598 (
            .O(N__21851),
            .I(\b2v_inst11.mult1_un138_sum_cry_3_s ));
    InMux I__3597 (
            .O(N__21848),
            .I(\b2v_inst11.mult1_un145_sum_cry_3 ));
    InMux I__3596 (
            .O(N__21845),
            .I(N__21842));
    LocalMux I__3595 (
            .O(N__21842),
            .I(\b2v_inst11.mult1_un138_sum_cry_4_s ));
    InMux I__3594 (
            .O(N__21839),
            .I(\b2v_inst11.mult1_un145_sum_cry_4 ));
    InMux I__3593 (
            .O(N__21836),
            .I(N__21832));
    CascadeMux I__3592 (
            .O(N__21835),
            .I(N__21828));
    LocalMux I__3591 (
            .O(N__21832),
            .I(N__21824));
    InMux I__3590 (
            .O(N__21831),
            .I(N__21819));
    InMux I__3589 (
            .O(N__21828),
            .I(N__21819));
    InMux I__3588 (
            .O(N__21827),
            .I(N__21816));
    Odrv4 I__3587 (
            .O(N__21824),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    LocalMux I__3586 (
            .O(N__21819),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    LocalMux I__3585 (
            .O(N__21816),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    CascadeMux I__3584 (
            .O(N__21809),
            .I(N__21806));
    InMux I__3583 (
            .O(N__21806),
            .I(N__21803));
    LocalMux I__3582 (
            .O(N__21803),
            .I(\b2v_inst11.mult1_un138_sum_cry_5_s ));
    InMux I__3581 (
            .O(N__21800),
            .I(\b2v_inst11.mult1_un145_sum_cry_5 ));
    InMux I__3580 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__3579 (
            .O(N__21794),
            .I(\b2v_inst5.count_1_6 ));
    InMux I__3578 (
            .O(N__21791),
            .I(N__21788));
    LocalMux I__3577 (
            .O(N__21788),
            .I(N__21785));
    Span4Mux_v I__3576 (
            .O(N__21785),
            .I(N__21782));
    Span4Mux_h I__3575 (
            .O(N__21782),
            .I(N__21779));
    Span4Mux_v I__3574 (
            .O(N__21779),
            .I(N__21776));
    Odrv4 I__3573 (
            .O(N__21776),
            .I(vr_ready_vccinaux));
    InMux I__3572 (
            .O(N__21773),
            .I(N__21770));
    LocalMux I__3571 (
            .O(N__21770),
            .I(N__21767));
    Span12Mux_s7_v I__3570 (
            .O(N__21767),
            .I(N__21764));
    Odrv12 I__3569 (
            .O(N__21764),
            .I(vr_ready_vccin));
    InMux I__3568 (
            .O(N__21761),
            .I(N__21758));
    LocalMux I__3567 (
            .O(N__21758),
            .I(N__21754));
    InMux I__3566 (
            .O(N__21757),
            .I(N__21751));
    Odrv4 I__3565 (
            .O(N__21754),
            .I(\b2v_inst11.mult1_un124_sum_cry_3_s ));
    LocalMux I__3564 (
            .O(N__21751),
            .I(\b2v_inst11.mult1_un124_sum_cry_3_s ));
    CascadeMux I__3563 (
            .O(N__21746),
            .I(N__21741));
    InMux I__3562 (
            .O(N__21745),
            .I(N__21737));
    InMux I__3561 (
            .O(N__21744),
            .I(N__21731));
    InMux I__3560 (
            .O(N__21741),
            .I(N__21731));
    InMux I__3559 (
            .O(N__21740),
            .I(N__21728));
    LocalMux I__3558 (
            .O(N__21737),
            .I(N__21724));
    InMux I__3557 (
            .O(N__21736),
            .I(N__21721));
    LocalMux I__3556 (
            .O(N__21731),
            .I(N__21716));
    LocalMux I__3555 (
            .O(N__21728),
            .I(N__21716));
    InMux I__3554 (
            .O(N__21727),
            .I(N__21713));
    Odrv12 I__3553 (
            .O(N__21724),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__3552 (
            .O(N__21721),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    Odrv4 I__3551 (
            .O(N__21716),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__3550 (
            .O(N__21713),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    CascadeMux I__3549 (
            .O(N__21704),
            .I(N__21701));
    InMux I__3548 (
            .O(N__21701),
            .I(N__21698));
    LocalMux I__3547 (
            .O(N__21698),
            .I(\b2v_inst11.mult1_un131_sum_axb_4_l_fx ));
    InMux I__3546 (
            .O(N__21695),
            .I(N__21691));
    InMux I__3545 (
            .O(N__21694),
            .I(N__21688));
    LocalMux I__3544 (
            .O(N__21691),
            .I(N__21683));
    LocalMux I__3543 (
            .O(N__21688),
            .I(N__21683));
    Odrv12 I__3542 (
            .O(N__21683),
            .I(\b2v_inst11.mult1_un138_sum ));
    InMux I__3541 (
            .O(N__21680),
            .I(N__21677));
    LocalMux I__3540 (
            .O(N__21677),
            .I(N__21674));
    Odrv12 I__3539 (
            .O(N__21674),
            .I(\b2v_inst11.mult1_un131_sum_i ));
    InMux I__3538 (
            .O(N__21671),
            .I(\b2v_inst11.mult1_un138_sum_cry_2_c ));
    CascadeMux I__3537 (
            .O(N__21668),
            .I(N__21665));
    InMux I__3536 (
            .O(N__21665),
            .I(N__21662));
    LocalMux I__3535 (
            .O(N__21662),
            .I(\b2v_inst11.mult1_un131_sum_cry_3_s ));
    InMux I__3534 (
            .O(N__21659),
            .I(\b2v_inst11.mult1_un138_sum_cry_3_c ));
    InMux I__3533 (
            .O(N__21656),
            .I(N__21653));
    LocalMux I__3532 (
            .O(N__21653),
            .I(\b2v_inst11.mult1_un131_sum_cry_4_s ));
    InMux I__3531 (
            .O(N__21650),
            .I(\b2v_inst11.mult1_un138_sum_cry_4_c ));
    CascadeMux I__3530 (
            .O(N__21647),
            .I(N__21642));
    InMux I__3529 (
            .O(N__21646),
            .I(N__21638));
    InMux I__3528 (
            .O(N__21645),
            .I(N__21633));
    InMux I__3527 (
            .O(N__21642),
            .I(N__21633));
    InMux I__3526 (
            .O(N__21641),
            .I(N__21630));
    LocalMux I__3525 (
            .O(N__21638),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__3524 (
            .O(N__21633),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__3523 (
            .O(N__21630),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    CascadeMux I__3522 (
            .O(N__21623),
            .I(N__21620));
    InMux I__3521 (
            .O(N__21620),
            .I(N__21617));
    LocalMux I__3520 (
            .O(N__21617),
            .I(\b2v_inst11.mult1_un131_sum_cry_5_s ));
    CascadeMux I__3519 (
            .O(N__21614),
            .I(N__21611));
    InMux I__3518 (
            .O(N__21611),
            .I(N__21608));
    LocalMux I__3517 (
            .O(N__21608),
            .I(N__21605));
    Odrv4 I__3516 (
            .O(N__21605),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ));
    CascadeMux I__3515 (
            .O(N__21602),
            .I(N__21598));
    CascadeMux I__3514 (
            .O(N__21601),
            .I(N__21595));
    InMux I__3513 (
            .O(N__21598),
            .I(N__21590));
    InMux I__3512 (
            .O(N__21595),
            .I(N__21590));
    LocalMux I__3511 (
            .O(N__21590),
            .I(\b2v_inst11.mult1_un47_sum ));
    InMux I__3510 (
            .O(N__21587),
            .I(\b2v_inst11.un1_dutycycle_53_cry_13 ));
    CascadeMux I__3509 (
            .O(N__21584),
            .I(N__21579));
    InMux I__3508 (
            .O(N__21583),
            .I(N__21569));
    InMux I__3507 (
            .O(N__21582),
            .I(N__21569));
    InMux I__3506 (
            .O(N__21579),
            .I(N__21569));
    InMux I__3505 (
            .O(N__21578),
            .I(N__21569));
    LocalMux I__3504 (
            .O(N__21569),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ));
    InMux I__3503 (
            .O(N__21566),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14 ));
    CascadeMux I__3502 (
            .O(N__21563),
            .I(N__21559));
    InMux I__3501 (
            .O(N__21562),
            .I(N__21551));
    InMux I__3500 (
            .O(N__21559),
            .I(N__21551));
    InMux I__3499 (
            .O(N__21558),
            .I(N__21551));
    LocalMux I__3498 (
            .O(N__21551),
            .I(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ));
    InMux I__3497 (
            .O(N__21548),
            .I(bfn_6_11_0_));
    InMux I__3496 (
            .O(N__21545),
            .I(\b2v_inst11.CO2 ));
    CascadeMux I__3495 (
            .O(N__21542),
            .I(N__21539));
    InMux I__3494 (
            .O(N__21539),
            .I(N__21533));
    InMux I__3493 (
            .O(N__21538),
            .I(N__21533));
    LocalMux I__3492 (
            .O(N__21533),
            .I(\b2v_inst11.CO2_THRU_CO ));
    InMux I__3491 (
            .O(N__21530),
            .I(N__21526));
    InMux I__3490 (
            .O(N__21529),
            .I(N__21523));
    LocalMux I__3489 (
            .O(N__21526),
            .I(N__21518));
    LocalMux I__3488 (
            .O(N__21523),
            .I(N__21518));
    Span4Mux_v I__3487 (
            .O(N__21518),
            .I(N__21515));
    Odrv4 I__3486 (
            .O(N__21515),
            .I(\b2v_inst11.mult1_un131_sum ));
    InMux I__3485 (
            .O(N__21512),
            .I(N__21509));
    LocalMux I__3484 (
            .O(N__21509),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_14 ));
    CascadeMux I__3483 (
            .O(N__21506),
            .I(N__21503));
    InMux I__3482 (
            .O(N__21503),
            .I(N__21500));
    LocalMux I__3481 (
            .O(N__21500),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_5 ));
    InMux I__3480 (
            .O(N__21497),
            .I(N__21493));
    InMux I__3479 (
            .O(N__21496),
            .I(N__21490));
    LocalMux I__3478 (
            .O(N__21493),
            .I(N__21487));
    LocalMux I__3477 (
            .O(N__21490),
            .I(N__21484));
    Span4Mux_h I__3476 (
            .O(N__21487),
            .I(N__21481));
    Span4Mux_v I__3475 (
            .O(N__21484),
            .I(N__21478));
    Odrv4 I__3474 (
            .O(N__21481),
            .I(\b2v_inst11.mult1_un103_sum ));
    Odrv4 I__3473 (
            .O(N__21478),
            .I(\b2v_inst11.mult1_un103_sum ));
    InMux I__3472 (
            .O(N__21473),
            .I(\b2v_inst11.un1_dutycycle_53_cry_5 ));
    CascadeMux I__3471 (
            .O(N__21470),
            .I(N__21467));
    InMux I__3470 (
            .O(N__21467),
            .I(N__21464));
    LocalMux I__3469 (
            .O(N__21464),
            .I(N__21461));
    Span4Mux_v I__3468 (
            .O(N__21461),
            .I(N__21458));
    Odrv4 I__3467 (
            .O(N__21458),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_10 ));
    InMux I__3466 (
            .O(N__21455),
            .I(N__21451));
    InMux I__3465 (
            .O(N__21454),
            .I(N__21448));
    LocalMux I__3464 (
            .O(N__21451),
            .I(N__21445));
    LocalMux I__3463 (
            .O(N__21448),
            .I(N__21440));
    Span4Mux_s1_h I__3462 (
            .O(N__21445),
            .I(N__21440));
    Span4Mux_h I__3461 (
            .O(N__21440),
            .I(N__21437));
    Odrv4 I__3460 (
            .O(N__21437),
            .I(\b2v_inst11.mult1_un96_sum ));
    InMux I__3459 (
            .O(N__21434),
            .I(\b2v_inst11.un1_dutycycle_53_cry_6 ));
    CascadeMux I__3458 (
            .O(N__21431),
            .I(N__21428));
    InMux I__3457 (
            .O(N__21428),
            .I(N__21425));
    LocalMux I__3456 (
            .O(N__21425),
            .I(N__21422));
    Odrv4 I__3455 (
            .O(N__21422),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_11 ));
    InMux I__3454 (
            .O(N__21419),
            .I(N__21415));
    InMux I__3453 (
            .O(N__21418),
            .I(N__21412));
    LocalMux I__3452 (
            .O(N__21415),
            .I(N__21409));
    LocalMux I__3451 (
            .O(N__21412),
            .I(N__21404));
    Span4Mux_s1_h I__3450 (
            .O(N__21409),
            .I(N__21404));
    Span4Mux_h I__3449 (
            .O(N__21404),
            .I(N__21401));
    Odrv4 I__3448 (
            .O(N__21401),
            .I(\b2v_inst11.mult1_un89_sum ));
    InMux I__3447 (
            .O(N__21398),
            .I(bfn_6_10_0_));
    CascadeMux I__3446 (
            .O(N__21395),
            .I(N__21392));
    InMux I__3445 (
            .O(N__21392),
            .I(N__21389));
    LocalMux I__3444 (
            .O(N__21389),
            .I(N__21386));
    Odrv4 I__3443 (
            .O(N__21386),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_12 ));
    InMux I__3442 (
            .O(N__21383),
            .I(N__21380));
    LocalMux I__3441 (
            .O(N__21380),
            .I(N__21376));
    InMux I__3440 (
            .O(N__21379),
            .I(N__21373));
    Span4Mux_h I__3439 (
            .O(N__21376),
            .I(N__21370));
    LocalMux I__3438 (
            .O(N__21373),
            .I(N__21367));
    Odrv4 I__3437 (
            .O(N__21370),
            .I(\b2v_inst11.mult1_un82_sum ));
    Odrv12 I__3436 (
            .O(N__21367),
            .I(\b2v_inst11.mult1_un82_sum ));
    InMux I__3435 (
            .O(N__21362),
            .I(\b2v_inst11.un1_dutycycle_53_cry_8 ));
    InMux I__3434 (
            .O(N__21359),
            .I(N__21356));
    LocalMux I__3433 (
            .O(N__21356),
            .I(N__21353));
    Span4Mux_v I__3432 (
            .O(N__21353),
            .I(N__21350));
    Odrv4 I__3431 (
            .O(N__21350),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_13 ));
    InMux I__3430 (
            .O(N__21347),
            .I(N__21343));
    InMux I__3429 (
            .O(N__21346),
            .I(N__21340));
    LocalMux I__3428 (
            .O(N__21343),
            .I(N__21337));
    LocalMux I__3427 (
            .O(N__21340),
            .I(N__21334));
    Odrv4 I__3426 (
            .O(N__21337),
            .I(\b2v_inst11.mult1_un75_sum ));
    Odrv12 I__3425 (
            .O(N__21334),
            .I(\b2v_inst11.mult1_un75_sum ));
    InMux I__3424 (
            .O(N__21329),
            .I(\b2v_inst11.un1_dutycycle_53_cry_9 ));
    InMux I__3423 (
            .O(N__21326),
            .I(N__21323));
    LocalMux I__3422 (
            .O(N__21323),
            .I(N__21320));
    Span4Mux_h I__3421 (
            .O(N__21320),
            .I(N__21317));
    Odrv4 I__3420 (
            .O(N__21317),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_14 ));
    CascadeMux I__3419 (
            .O(N__21314),
            .I(N__21310));
    InMux I__3418 (
            .O(N__21313),
            .I(N__21307));
    InMux I__3417 (
            .O(N__21310),
            .I(N__21304));
    LocalMux I__3416 (
            .O(N__21307),
            .I(N__21301));
    LocalMux I__3415 (
            .O(N__21304),
            .I(N__21298));
    Span4Mux_v I__3414 (
            .O(N__21301),
            .I(N__21295));
    Span12Mux_s5_h I__3413 (
            .O(N__21298),
            .I(N__21292));
    Odrv4 I__3412 (
            .O(N__21295),
            .I(\b2v_inst11.mult1_un68_sum ));
    Odrv12 I__3411 (
            .O(N__21292),
            .I(\b2v_inst11.mult1_un68_sum ));
    InMux I__3410 (
            .O(N__21287),
            .I(\b2v_inst11.un1_dutycycle_53_cry_10 ));
    CascadeMux I__3409 (
            .O(N__21284),
            .I(N__21281));
    InMux I__3408 (
            .O(N__21281),
            .I(N__21278));
    LocalMux I__3407 (
            .O(N__21278),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_15 ));
    InMux I__3406 (
            .O(N__21275),
            .I(N__21271));
    InMux I__3405 (
            .O(N__21274),
            .I(N__21268));
    LocalMux I__3404 (
            .O(N__21271),
            .I(N__21265));
    LocalMux I__3403 (
            .O(N__21268),
            .I(N__21262));
    Span4Mux_h I__3402 (
            .O(N__21265),
            .I(N__21259));
    Odrv4 I__3401 (
            .O(N__21262),
            .I(\b2v_inst11.mult1_un61_sum ));
    Odrv4 I__3400 (
            .O(N__21259),
            .I(\b2v_inst11.mult1_un61_sum ));
    InMux I__3399 (
            .O(N__21254),
            .I(\b2v_inst11.un1_dutycycle_53_cry_11 ));
    CascadeMux I__3398 (
            .O(N__21251),
            .I(N__21248));
    InMux I__3397 (
            .O(N__21248),
            .I(N__21245));
    LocalMux I__3396 (
            .O(N__21245),
            .I(N__21242));
    Span4Mux_h I__3395 (
            .O(N__21242),
            .I(N__21239));
    Odrv4 I__3394 (
            .O(N__21239),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_13 ));
    CascadeMux I__3393 (
            .O(N__21236),
            .I(N__21233));
    InMux I__3392 (
            .O(N__21233),
            .I(N__21229));
    InMux I__3391 (
            .O(N__21232),
            .I(N__21226));
    LocalMux I__3390 (
            .O(N__21229),
            .I(N__21223));
    LocalMux I__3389 (
            .O(N__21226),
            .I(N__21220));
    Span4Mux_h I__3388 (
            .O(N__21223),
            .I(N__21217));
    Odrv4 I__3387 (
            .O(N__21220),
            .I(\b2v_inst11.mult1_un54_sum ));
    Odrv4 I__3386 (
            .O(N__21217),
            .I(\b2v_inst11.mult1_un54_sum ));
    InMux I__3385 (
            .O(N__21212),
            .I(\b2v_inst11.un1_dutycycle_53_cry_12 ));
    InMux I__3384 (
            .O(N__21209),
            .I(N__21206));
    LocalMux I__3383 (
            .O(N__21206),
            .I(\b2v_inst11.d_i3_mux ));
    InMux I__3382 (
            .O(N__21203),
            .I(N__21200));
    LocalMux I__3381 (
            .O(N__21200),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_0 ));
    InMux I__3380 (
            .O(N__21197),
            .I(\b2v_inst11.un1_dutycycle_53_cry_0 ));
    InMux I__3379 (
            .O(N__21194),
            .I(\b2v_inst11.un1_dutycycle_53_cry_1 ));
    InMux I__3378 (
            .O(N__21191),
            .I(N__21188));
    LocalMux I__3377 (
            .O(N__21188),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_2 ));
    InMux I__3376 (
            .O(N__21185),
            .I(N__21181));
    InMux I__3375 (
            .O(N__21184),
            .I(N__21178));
    LocalMux I__3374 (
            .O(N__21181),
            .I(N__21175));
    LocalMux I__3373 (
            .O(N__21178),
            .I(N__21172));
    Span4Mux_h I__3372 (
            .O(N__21175),
            .I(N__21167));
    Span4Mux_v I__3371 (
            .O(N__21172),
            .I(N__21167));
    Odrv4 I__3370 (
            .O(N__21167),
            .I(\b2v_inst11.mult1_un124_sum ));
    InMux I__3369 (
            .O(N__21164),
            .I(\b2v_inst11.un1_dutycycle_53_cry_2 ));
    InMux I__3368 (
            .O(N__21161),
            .I(N__21157));
    InMux I__3367 (
            .O(N__21160),
            .I(N__21154));
    LocalMux I__3366 (
            .O(N__21157),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_7 ));
    LocalMux I__3365 (
            .O(N__21154),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_7 ));
    CascadeMux I__3364 (
            .O(N__21149),
            .I(N__21146));
    InMux I__3363 (
            .O(N__21146),
            .I(N__21143));
    LocalMux I__3362 (
            .O(N__21143),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ));
    InMux I__3361 (
            .O(N__21140),
            .I(N__21136));
    InMux I__3360 (
            .O(N__21139),
            .I(N__21133));
    LocalMux I__3359 (
            .O(N__21136),
            .I(N__21130));
    LocalMux I__3358 (
            .O(N__21133),
            .I(N__21125));
    Span4Mux_h I__3357 (
            .O(N__21130),
            .I(N__21125));
    Span4Mux_v I__3356 (
            .O(N__21125),
            .I(N__21122));
    Odrv4 I__3355 (
            .O(N__21122),
            .I(\b2v_inst11.mult1_un117_sum ));
    InMux I__3354 (
            .O(N__21119),
            .I(\b2v_inst11.un1_dutycycle_53_cry_3 ));
    InMux I__3353 (
            .O(N__21116),
            .I(N__21113));
    LocalMux I__3352 (
            .O(N__21113),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_7 ));
    InMux I__3351 (
            .O(N__21110),
            .I(N__21106));
    InMux I__3350 (
            .O(N__21109),
            .I(N__21103));
    LocalMux I__3349 (
            .O(N__21106),
            .I(N__21100));
    LocalMux I__3348 (
            .O(N__21103),
            .I(N__21097));
    Span12Mux_s5_h I__3347 (
            .O(N__21100),
            .I(N__21094));
    Odrv4 I__3346 (
            .O(N__21097),
            .I(\b2v_inst11.mult1_un110_sum ));
    Odrv12 I__3345 (
            .O(N__21094),
            .I(\b2v_inst11.mult1_un110_sum ));
    InMux I__3344 (
            .O(N__21089),
            .I(\b2v_inst11.un1_dutycycle_53_cry_4 ));
    CascadeMux I__3343 (
            .O(N__21086),
            .I(\b2v_inst11.dutycycleZ0Z_7_cascade_ ));
    InMux I__3342 (
            .O(N__21083),
            .I(N__21080));
    LocalMux I__3341 (
            .O(N__21080),
            .I(\b2v_inst11.dutycycle_RNI_8Z0Z_7 ));
    CascadeMux I__3340 (
            .O(N__21077),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_4_cascade_ ));
    CascadeMux I__3339 (
            .O(N__21074),
            .I(\b2v_inst11.un1_dutycycle_53_axb_8_cascade_ ));
    InMux I__3338 (
            .O(N__21071),
            .I(N__21068));
    LocalMux I__3337 (
            .O(N__21068),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ));
    CascadeMux I__3336 (
            .O(N__21065),
            .I(\b2v_inst11.un1_dutycycle_53_axb_3_1_0_cascade_ ));
    CascadeMux I__3335 (
            .O(N__21062),
            .I(\b2v_inst11.un1_dutycycle_53_axb_3_cascade_ ));
    CascadeMux I__3334 (
            .O(N__21059),
            .I(\b2v_inst11.un1_i3_mux_cascade_ ));
    InMux I__3333 (
            .O(N__21056),
            .I(N__21050));
    InMux I__3332 (
            .O(N__21055),
            .I(N__21050));
    LocalMux I__3331 (
            .O(N__21050),
            .I(\b2v_inst11.dutycycleZ1Z_8 ));
    InMux I__3330 (
            .O(N__21047),
            .I(N__21044));
    LocalMux I__3329 (
            .O(N__21044),
            .I(\b2v_inst11.un1_dutycycle_53_3_0_tz ));
    CascadeMux I__3328 (
            .O(N__21041),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_3_cascade_ ));
    CascadeMux I__3327 (
            .O(N__21038),
            .I(\b2v_inst11.N_26_i_1_cascade_ ));
    InMux I__3326 (
            .O(N__21035),
            .I(N__21032));
    LocalMux I__3325 (
            .O(N__21032),
            .I(N__21029));
    Odrv4 I__3324 (
            .O(N__21029),
            .I(\b2v_inst11.un1_dutycycle_53_axb_9_1 ));
    InMux I__3323 (
            .O(N__21026),
            .I(N__21020));
    InMux I__3322 (
            .O(N__21025),
            .I(N__21020));
    LocalMux I__3321 (
            .O(N__21020),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    CascadeMux I__3320 (
            .O(N__21017),
            .I(N__21013));
    InMux I__3319 (
            .O(N__21016),
            .I(N__21008));
    InMux I__3318 (
            .O(N__21013),
            .I(N__21008));
    LocalMux I__3317 (
            .O(N__21008),
            .I(\b2v_inst11.dutycycleZ1Z_4 ));
    CascadeMux I__3316 (
            .O(N__21005),
            .I(N__21001));
    InMux I__3315 (
            .O(N__21004),
            .I(N__20998));
    InMux I__3314 (
            .O(N__21001),
            .I(N__20995));
    LocalMux I__3313 (
            .O(N__20998),
            .I(\b2v_inst20.counterZ0Z_27 ));
    LocalMux I__3312 (
            .O(N__20995),
            .I(\b2v_inst20.counterZ0Z_27 ));
    InMux I__3311 (
            .O(N__20990),
            .I(\b2v_inst20.counter_1_cry_26 ));
    InMux I__3310 (
            .O(N__20987),
            .I(\b2v_inst20.counter_1_cry_27 ));
    InMux I__3309 (
            .O(N__20984),
            .I(\b2v_inst20.counter_1_cry_28 ));
    InMux I__3308 (
            .O(N__20981),
            .I(\b2v_inst20.counter_1_cry_29 ));
    InMux I__3307 (
            .O(N__20978),
            .I(\b2v_inst20.counter_1_cry_30 ));
    CascadeMux I__3306 (
            .O(N__20975),
            .I(N__20972));
    InMux I__3305 (
            .O(N__20972),
            .I(N__20966));
    InMux I__3304 (
            .O(N__20971),
            .I(N__20966));
    LocalMux I__3303 (
            .O(N__20966),
            .I(\b2v_inst20.counterZ0Z_28 ));
    CascadeMux I__3302 (
            .O(N__20963),
            .I(N__20960));
    InMux I__3301 (
            .O(N__20960),
            .I(N__20954));
    InMux I__3300 (
            .O(N__20959),
            .I(N__20954));
    LocalMux I__3299 (
            .O(N__20954),
            .I(\b2v_inst20.counterZ0Z_29 ));
    CascadeMux I__3298 (
            .O(N__20951),
            .I(N__20947));
    CascadeMux I__3297 (
            .O(N__20950),
            .I(N__20944));
    InMux I__3296 (
            .O(N__20947),
            .I(N__20939));
    InMux I__3295 (
            .O(N__20944),
            .I(N__20939));
    LocalMux I__3294 (
            .O(N__20939),
            .I(\b2v_inst20.counterZ0Z_30 ));
    InMux I__3293 (
            .O(N__20936),
            .I(N__20930));
    InMux I__3292 (
            .O(N__20935),
            .I(N__20930));
    LocalMux I__3291 (
            .O(N__20930),
            .I(\b2v_inst20.counterZ0Z_31 ));
    InMux I__3290 (
            .O(N__20927),
            .I(N__20924));
    LocalMux I__3289 (
            .O(N__20924),
            .I(\b2v_inst20.un4_counter_7_and ));
    InMux I__3288 (
            .O(N__20921),
            .I(N__20918));
    LocalMux I__3287 (
            .O(N__20918),
            .I(\b2v_inst11.un1_dutycycle_53_9_1_1 ));
    CascadeMux I__3286 (
            .O(N__20915),
            .I(\b2v_inst11.dutycycleZ1Z_5_cascade_ ));
    InMux I__3285 (
            .O(N__20912),
            .I(N__20908));
    InMux I__3284 (
            .O(N__20911),
            .I(N__20905));
    LocalMux I__3283 (
            .O(N__20908),
            .I(\b2v_inst20.counterZ0Z_19 ));
    LocalMux I__3282 (
            .O(N__20905),
            .I(\b2v_inst20.counterZ0Z_19 ));
    InMux I__3281 (
            .O(N__20900),
            .I(\b2v_inst20.counter_1_cry_18 ));
    CascadeMux I__3280 (
            .O(N__20897),
            .I(N__20893));
    InMux I__3279 (
            .O(N__20896),
            .I(N__20890));
    InMux I__3278 (
            .O(N__20893),
            .I(N__20887));
    LocalMux I__3277 (
            .O(N__20890),
            .I(\b2v_inst20.counterZ0Z_20 ));
    LocalMux I__3276 (
            .O(N__20887),
            .I(\b2v_inst20.counterZ0Z_20 ));
    InMux I__3275 (
            .O(N__20882),
            .I(\b2v_inst20.counter_1_cry_19 ));
    InMux I__3274 (
            .O(N__20879),
            .I(N__20875));
    InMux I__3273 (
            .O(N__20878),
            .I(N__20872));
    LocalMux I__3272 (
            .O(N__20875),
            .I(\b2v_inst20.counterZ0Z_21 ));
    LocalMux I__3271 (
            .O(N__20872),
            .I(\b2v_inst20.counterZ0Z_21 ));
    InMux I__3270 (
            .O(N__20867),
            .I(\b2v_inst20.counter_1_cry_20 ));
    InMux I__3269 (
            .O(N__20864),
            .I(N__20860));
    InMux I__3268 (
            .O(N__20863),
            .I(N__20857));
    LocalMux I__3267 (
            .O(N__20860),
            .I(\b2v_inst20.counterZ0Z_22 ));
    LocalMux I__3266 (
            .O(N__20857),
            .I(\b2v_inst20.counterZ0Z_22 ));
    InMux I__3265 (
            .O(N__20852),
            .I(\b2v_inst20.counter_1_cry_21 ));
    InMux I__3264 (
            .O(N__20849),
            .I(N__20845));
    InMux I__3263 (
            .O(N__20848),
            .I(N__20842));
    LocalMux I__3262 (
            .O(N__20845),
            .I(\b2v_inst20.counterZ0Z_23 ));
    LocalMux I__3261 (
            .O(N__20842),
            .I(\b2v_inst20.counterZ0Z_23 ));
    InMux I__3260 (
            .O(N__20837),
            .I(\b2v_inst20.counter_1_cry_22 ));
    InMux I__3259 (
            .O(N__20834),
            .I(N__20830));
    InMux I__3258 (
            .O(N__20833),
            .I(N__20827));
    LocalMux I__3257 (
            .O(N__20830),
            .I(\b2v_inst20.counterZ0Z_24 ));
    LocalMux I__3256 (
            .O(N__20827),
            .I(\b2v_inst20.counterZ0Z_24 ));
    InMux I__3255 (
            .O(N__20822),
            .I(\b2v_inst20.counter_1_cry_23 ));
    InMux I__3254 (
            .O(N__20819),
            .I(N__20815));
    InMux I__3253 (
            .O(N__20818),
            .I(N__20812));
    LocalMux I__3252 (
            .O(N__20815),
            .I(\b2v_inst20.counterZ0Z_25 ));
    LocalMux I__3251 (
            .O(N__20812),
            .I(\b2v_inst20.counterZ0Z_25 ));
    InMux I__3250 (
            .O(N__20807),
            .I(bfn_6_5_0_));
    InMux I__3249 (
            .O(N__20804),
            .I(N__20800));
    InMux I__3248 (
            .O(N__20803),
            .I(N__20797));
    LocalMux I__3247 (
            .O(N__20800),
            .I(\b2v_inst20.counterZ0Z_26 ));
    LocalMux I__3246 (
            .O(N__20797),
            .I(\b2v_inst20.counterZ0Z_26 ));
    InMux I__3245 (
            .O(N__20792),
            .I(\b2v_inst20.counter_1_cry_25 ));
    CascadeMux I__3244 (
            .O(N__20789),
            .I(N__20785));
    InMux I__3243 (
            .O(N__20788),
            .I(N__20782));
    InMux I__3242 (
            .O(N__20785),
            .I(N__20779));
    LocalMux I__3241 (
            .O(N__20782),
            .I(\b2v_inst20.counterZ0Z_10 ));
    LocalMux I__3240 (
            .O(N__20779),
            .I(\b2v_inst20.counterZ0Z_10 ));
    InMux I__3239 (
            .O(N__20774),
            .I(\b2v_inst20.counter_1_cry_9 ));
    InMux I__3238 (
            .O(N__20771),
            .I(N__20767));
    InMux I__3237 (
            .O(N__20770),
            .I(N__20764));
    LocalMux I__3236 (
            .O(N__20767),
            .I(\b2v_inst20.counterZ0Z_11 ));
    LocalMux I__3235 (
            .O(N__20764),
            .I(\b2v_inst20.counterZ0Z_11 ));
    InMux I__3234 (
            .O(N__20759),
            .I(\b2v_inst20.counter_1_cry_10 ));
    InMux I__3233 (
            .O(N__20756),
            .I(N__20752));
    InMux I__3232 (
            .O(N__20755),
            .I(N__20749));
    LocalMux I__3231 (
            .O(N__20752),
            .I(\b2v_inst20.counterZ0Z_12 ));
    LocalMux I__3230 (
            .O(N__20749),
            .I(\b2v_inst20.counterZ0Z_12 ));
    InMux I__3229 (
            .O(N__20744),
            .I(\b2v_inst20.counter_1_cry_11 ));
    InMux I__3228 (
            .O(N__20741),
            .I(N__20737));
    InMux I__3227 (
            .O(N__20740),
            .I(N__20734));
    LocalMux I__3226 (
            .O(N__20737),
            .I(\b2v_inst20.counterZ0Z_13 ));
    LocalMux I__3225 (
            .O(N__20734),
            .I(\b2v_inst20.counterZ0Z_13 ));
    InMux I__3224 (
            .O(N__20729),
            .I(\b2v_inst20.counter_1_cry_12 ));
    CascadeMux I__3223 (
            .O(N__20726),
            .I(N__20722));
    InMux I__3222 (
            .O(N__20725),
            .I(N__20719));
    InMux I__3221 (
            .O(N__20722),
            .I(N__20716));
    LocalMux I__3220 (
            .O(N__20719),
            .I(\b2v_inst20.counterZ0Z_14 ));
    LocalMux I__3219 (
            .O(N__20716),
            .I(\b2v_inst20.counterZ0Z_14 ));
    InMux I__3218 (
            .O(N__20711),
            .I(\b2v_inst20.counter_1_cry_13 ));
    InMux I__3217 (
            .O(N__20708),
            .I(N__20704));
    InMux I__3216 (
            .O(N__20707),
            .I(N__20701));
    LocalMux I__3215 (
            .O(N__20704),
            .I(\b2v_inst20.counterZ0Z_15 ));
    LocalMux I__3214 (
            .O(N__20701),
            .I(\b2v_inst20.counterZ0Z_15 ));
    InMux I__3213 (
            .O(N__20696),
            .I(\b2v_inst20.counter_1_cry_14 ));
    InMux I__3212 (
            .O(N__20693),
            .I(N__20689));
    InMux I__3211 (
            .O(N__20692),
            .I(N__20686));
    LocalMux I__3210 (
            .O(N__20689),
            .I(\b2v_inst20.counterZ0Z_16 ));
    LocalMux I__3209 (
            .O(N__20686),
            .I(\b2v_inst20.counterZ0Z_16 ));
    InMux I__3208 (
            .O(N__20681),
            .I(\b2v_inst20.counter_1_cry_15 ));
    CascadeMux I__3207 (
            .O(N__20678),
            .I(N__20674));
    InMux I__3206 (
            .O(N__20677),
            .I(N__20671));
    InMux I__3205 (
            .O(N__20674),
            .I(N__20668));
    LocalMux I__3204 (
            .O(N__20671),
            .I(\b2v_inst20.counterZ0Z_17 ));
    LocalMux I__3203 (
            .O(N__20668),
            .I(\b2v_inst20.counterZ0Z_17 ));
    InMux I__3202 (
            .O(N__20663),
            .I(bfn_6_4_0_));
    InMux I__3201 (
            .O(N__20660),
            .I(N__20656));
    InMux I__3200 (
            .O(N__20659),
            .I(N__20653));
    LocalMux I__3199 (
            .O(N__20656),
            .I(\b2v_inst20.counterZ0Z_18 ));
    LocalMux I__3198 (
            .O(N__20653),
            .I(\b2v_inst20.counterZ0Z_18 ));
    InMux I__3197 (
            .O(N__20648),
            .I(\b2v_inst20.counter_1_cry_17 ));
    InMux I__3196 (
            .O(N__20645),
            .I(\b2v_inst20.counter_1_cry_1 ));
    InMux I__3195 (
            .O(N__20642),
            .I(\b2v_inst20.counter_1_cry_2 ));
    InMux I__3194 (
            .O(N__20639),
            .I(\b2v_inst20.counter_1_cry_3 ));
    InMux I__3193 (
            .O(N__20636),
            .I(\b2v_inst20.counter_1_cry_4 ));
    InMux I__3192 (
            .O(N__20633),
            .I(\b2v_inst20.counter_1_cry_5 ));
    InMux I__3191 (
            .O(N__20630),
            .I(\b2v_inst20.counter_1_cry_6 ));
    InMux I__3190 (
            .O(N__20627),
            .I(N__20623));
    InMux I__3189 (
            .O(N__20626),
            .I(N__20620));
    LocalMux I__3188 (
            .O(N__20623),
            .I(\b2v_inst20.counterZ0Z_8 ));
    LocalMux I__3187 (
            .O(N__20620),
            .I(\b2v_inst20.counterZ0Z_8 ));
    InMux I__3186 (
            .O(N__20615),
            .I(\b2v_inst20.counter_1_cry_7 ));
    InMux I__3185 (
            .O(N__20612),
            .I(N__20608));
    InMux I__3184 (
            .O(N__20611),
            .I(N__20605));
    LocalMux I__3183 (
            .O(N__20608),
            .I(\b2v_inst20.counterZ0Z_9 ));
    LocalMux I__3182 (
            .O(N__20605),
            .I(\b2v_inst20.counterZ0Z_9 ));
    InMux I__3181 (
            .O(N__20600),
            .I(bfn_6_3_0_));
    CascadeMux I__3180 (
            .O(N__20597),
            .I(N__20594));
    InMux I__3179 (
            .O(N__20594),
            .I(N__20591));
    LocalMux I__3178 (
            .O(N__20591),
            .I(\b2v_inst11.mult1_un159_sum_cry_2_s ));
    InMux I__3177 (
            .O(N__20588),
            .I(\b2v_inst11.mult1_un159_sum_cry_1 ));
    CascadeMux I__3176 (
            .O(N__20585),
            .I(N__20582));
    InMux I__3175 (
            .O(N__20582),
            .I(N__20579));
    LocalMux I__3174 (
            .O(N__20579),
            .I(\b2v_inst11.mult1_un159_sum_cry_3_s ));
    InMux I__3173 (
            .O(N__20576),
            .I(\b2v_inst11.mult1_un159_sum_cry_2 ));
    InMux I__3172 (
            .O(N__20573),
            .I(N__20570));
    LocalMux I__3171 (
            .O(N__20570),
            .I(\b2v_inst11.mult1_un159_sum_cry_4_s ));
    InMux I__3170 (
            .O(N__20567),
            .I(\b2v_inst11.mult1_un159_sum_cry_3 ));
    InMux I__3169 (
            .O(N__20564),
            .I(N__20561));
    LocalMux I__3168 (
            .O(N__20561),
            .I(\b2v_inst11.mult1_un159_sum_cry_5_s ));
    InMux I__3167 (
            .O(N__20558),
            .I(\b2v_inst11.mult1_un159_sum_cry_4 ));
    CascadeMux I__3166 (
            .O(N__20555),
            .I(N__20552));
    InMux I__3165 (
            .O(N__20552),
            .I(N__20549));
    LocalMux I__3164 (
            .O(N__20549),
            .I(\b2v_inst11.mult1_un166_sum_axb_6 ));
    InMux I__3163 (
            .O(N__20546),
            .I(\b2v_inst11.mult1_un159_sum_cry_5 ));
    InMux I__3162 (
            .O(N__20543),
            .I(\b2v_inst11.mult1_un159_sum_cry_6 ));
    InMux I__3161 (
            .O(N__20540),
            .I(N__20536));
    CascadeMux I__3160 (
            .O(N__20539),
            .I(N__20532));
    LocalMux I__3159 (
            .O(N__20536),
            .I(N__20527));
    InMux I__3158 (
            .O(N__20535),
            .I(N__20524));
    InMux I__3157 (
            .O(N__20532),
            .I(N__20517));
    InMux I__3156 (
            .O(N__20531),
            .I(N__20517));
    InMux I__3155 (
            .O(N__20530),
            .I(N__20517));
    Odrv12 I__3154 (
            .O(N__20527),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    LocalMux I__3153 (
            .O(N__20524),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    LocalMux I__3152 (
            .O(N__20517),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    CascadeMux I__3151 (
            .O(N__20510),
            .I(N__20507));
    InMux I__3150 (
            .O(N__20507),
            .I(N__20504));
    LocalMux I__3149 (
            .O(N__20504),
            .I(N__20501));
    Odrv4 I__3148 (
            .O(N__20501),
            .I(\b2v_inst11.mult1_un124_sum_i_0_8 ));
    InMux I__3147 (
            .O(N__20498),
            .I(N__20495));
    LocalMux I__3146 (
            .O(N__20495),
            .I(\b2v_inst11.mult1_un159_sum_i ));
    InMux I__3145 (
            .O(N__20492),
            .I(N__20489));
    LocalMux I__3144 (
            .O(N__20489),
            .I(N__20486));
    Odrv4 I__3143 (
            .O(N__20486),
            .I(\b2v_inst11.mult1_un117_sum_i ));
    InMux I__3142 (
            .O(N__20483),
            .I(\b2v_inst11.mult1_un124_sum_cry_2 ));
    CascadeMux I__3141 (
            .O(N__20480),
            .I(N__20477));
    InMux I__3140 (
            .O(N__20477),
            .I(N__20474));
    LocalMux I__3139 (
            .O(N__20474),
            .I(\b2v_inst11.mult1_un117_sum_cry_3_s ));
    InMux I__3138 (
            .O(N__20471),
            .I(N__20468));
    LocalMux I__3137 (
            .O(N__20468),
            .I(\b2v_inst11.mult1_un124_sum_cry_4_s ));
    InMux I__3136 (
            .O(N__20465),
            .I(\b2v_inst11.mult1_un124_sum_cry_3 ));
    InMux I__3135 (
            .O(N__20462),
            .I(N__20459));
    LocalMux I__3134 (
            .O(N__20459),
            .I(\b2v_inst11.mult1_un117_sum_cry_4_s ));
    CascadeMux I__3133 (
            .O(N__20456),
            .I(N__20453));
    InMux I__3132 (
            .O(N__20453),
            .I(N__20450));
    LocalMux I__3131 (
            .O(N__20450),
            .I(\b2v_inst11.mult1_un124_sum_cry_5_s ));
    InMux I__3130 (
            .O(N__20447),
            .I(\b2v_inst11.mult1_un124_sum_cry_4 ));
    InMux I__3129 (
            .O(N__20444),
            .I(N__20441));
    LocalMux I__3128 (
            .O(N__20441),
            .I(N__20437));
    CascadeMux I__3127 (
            .O(N__20440),
            .I(N__20433));
    Span4Mux_v I__3126 (
            .O(N__20437),
            .I(N__20429));
    InMux I__3125 (
            .O(N__20436),
            .I(N__20424));
    InMux I__3124 (
            .O(N__20433),
            .I(N__20424));
    InMux I__3123 (
            .O(N__20432),
            .I(N__20421));
    Odrv4 I__3122 (
            .O(N__20429),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__3121 (
            .O(N__20424),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__3120 (
            .O(N__20421),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    CascadeMux I__3119 (
            .O(N__20414),
            .I(N__20411));
    InMux I__3118 (
            .O(N__20411),
            .I(N__20408));
    LocalMux I__3117 (
            .O(N__20408),
            .I(\b2v_inst11.mult1_un117_sum_cry_5_s ));
    InMux I__3116 (
            .O(N__20405),
            .I(\b2v_inst11.mult1_un124_sum_cry_5 ));
    InMux I__3115 (
            .O(N__20402),
            .I(N__20399));
    LocalMux I__3114 (
            .O(N__20399),
            .I(\b2v_inst11.mult1_un117_sum_cry_6_s ));
    CascadeMux I__3113 (
            .O(N__20396),
            .I(N__20392));
    CascadeMux I__3112 (
            .O(N__20395),
            .I(N__20388));
    InMux I__3111 (
            .O(N__20392),
            .I(N__20381));
    InMux I__3110 (
            .O(N__20391),
            .I(N__20381));
    InMux I__3109 (
            .O(N__20388),
            .I(N__20381));
    LocalMux I__3108 (
            .O(N__20381),
            .I(\b2v_inst11.mult1_un117_sum_i_0_8 ));
    CascadeMux I__3107 (
            .O(N__20378),
            .I(N__20375));
    InMux I__3106 (
            .O(N__20375),
            .I(N__20372));
    LocalMux I__3105 (
            .O(N__20372),
            .I(\b2v_inst11.mult1_un131_sum_axb_8 ));
    InMux I__3104 (
            .O(N__20369),
            .I(\b2v_inst11.mult1_un124_sum_cry_6 ));
    CascadeMux I__3103 (
            .O(N__20366),
            .I(N__20363));
    InMux I__3102 (
            .O(N__20363),
            .I(N__20360));
    LocalMux I__3101 (
            .O(N__20360),
            .I(\b2v_inst11.mult1_un124_sum_axb_8 ));
    InMux I__3100 (
            .O(N__20357),
            .I(\b2v_inst11.mult1_un124_sum_cry_7 ));
    CascadeMux I__3099 (
            .O(N__20354),
            .I(\b2v_inst11.mult1_un124_sum_s_8_cascade_ ));
    InMux I__3098 (
            .O(N__20351),
            .I(N__20347));
    InMux I__3097 (
            .O(N__20350),
            .I(N__20344));
    LocalMux I__3096 (
            .O(N__20347),
            .I(\b2v_inst11.mult1_un124_sum_cry_6_s ));
    LocalMux I__3095 (
            .O(N__20344),
            .I(\b2v_inst11.mult1_un124_sum_cry_6_s ));
    CascadeMux I__3094 (
            .O(N__20339),
            .I(N__20336));
    InMux I__3093 (
            .O(N__20336),
            .I(N__20333));
    LocalMux I__3092 (
            .O(N__20333),
            .I(\b2v_inst11.mult1_un131_sum_axb_7_l_fx ));
    InMux I__3091 (
            .O(N__20330),
            .I(N__20327));
    LocalMux I__3090 (
            .O(N__20327),
            .I(N__20324));
    Sp12to4 I__3089 (
            .O(N__20324),
            .I(N__20321));
    Odrv12 I__3088 (
            .O(N__20321),
            .I(\b2v_inst11.g3_0 ));
    InMux I__3087 (
            .O(N__20318),
            .I(N__20315));
    LocalMux I__3086 (
            .O(N__20315),
            .I(\b2v_inst11.mult1_un124_sum_i ));
    InMux I__3085 (
            .O(N__20312),
            .I(\b2v_inst11.mult1_un131_sum_cry_2 ));
    InMux I__3084 (
            .O(N__20309),
            .I(\b2v_inst11.mult1_un131_sum_cry_3 ));
    InMux I__3083 (
            .O(N__20306),
            .I(\b2v_inst11.mult1_un131_sum_cry_4 ));
    InMux I__3082 (
            .O(N__20303),
            .I(\b2v_inst11.mult1_un131_sum_cry_5 ));
    InMux I__3081 (
            .O(N__20300),
            .I(\b2v_inst11.mult1_un131_sum_cry_6 ));
    InMux I__3080 (
            .O(N__20297),
            .I(\b2v_inst11.mult1_un131_sum_cry_7 ));
    CascadeMux I__3079 (
            .O(N__20294),
            .I(\b2v_inst11.mult1_un131_sum_s_8_cascade_ ));
    CascadeMux I__3078 (
            .O(N__20291),
            .I(N__20288));
    InMux I__3077 (
            .O(N__20288),
            .I(N__20285));
    LocalMux I__3076 (
            .O(N__20285),
            .I(\b2v_inst11.mult1_un124_sum_i_8 ));
    InMux I__3075 (
            .O(N__20282),
            .I(N__20279));
    LocalMux I__3074 (
            .O(N__20279),
            .I(\b2v_inst11.un85_clk_100khz_2 ));
    CascadeMux I__3073 (
            .O(N__20276),
            .I(N__20273));
    InMux I__3072 (
            .O(N__20273),
            .I(N__20270));
    LocalMux I__3071 (
            .O(N__20270),
            .I(\b2v_inst11.un85_clk_100khz_1 ));
    InMux I__3070 (
            .O(N__20267),
            .I(N__20264));
    LocalMux I__3069 (
            .O(N__20264),
            .I(N__20261));
    Odrv12 I__3068 (
            .O(N__20261),
            .I(\b2v_inst11.mult1_un96_sum_i ));
    InMux I__3067 (
            .O(N__20258),
            .I(N__20255));
    LocalMux I__3066 (
            .O(N__20255),
            .I(\b2v_inst11.mult1_un131_sum_i_8 ));
    InMux I__3065 (
            .O(N__20252),
            .I(N__20249));
    LocalMux I__3064 (
            .O(N__20249),
            .I(\b2v_inst11.un85_clk_100khz_3 ));
    CascadeMux I__3063 (
            .O(N__20246),
            .I(N__20242));
    InMux I__3062 (
            .O(N__20245),
            .I(N__20235));
    InMux I__3061 (
            .O(N__20242),
            .I(N__20235));
    InMux I__3060 (
            .O(N__20241),
            .I(N__20232));
    InMux I__3059 (
            .O(N__20240),
            .I(N__20229));
    LocalMux I__3058 (
            .O(N__20235),
            .I(N__20226));
    LocalMux I__3057 (
            .O(N__20232),
            .I(N__20222));
    LocalMux I__3056 (
            .O(N__20229),
            .I(N__20219));
    Span4Mux_h I__3055 (
            .O(N__20226),
            .I(N__20216));
    InMux I__3054 (
            .O(N__20225),
            .I(N__20213));
    Span4Mux_h I__3053 (
            .O(N__20222),
            .I(N__20210));
    Odrv12 I__3052 (
            .O(N__20219),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    Odrv4 I__3051 (
            .O(N__20216),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    LocalMux I__3050 (
            .O(N__20213),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    Odrv4 I__3049 (
            .O(N__20210),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    InMux I__3048 (
            .O(N__20201),
            .I(N__20198));
    LocalMux I__3047 (
            .O(N__20198),
            .I(\b2v_inst11.mult1_un103_sum_i_8 ));
    CascadeMux I__3046 (
            .O(N__20195),
            .I(N__20192));
    InMux I__3045 (
            .O(N__20192),
            .I(N__20189));
    LocalMux I__3044 (
            .O(N__20189),
            .I(\b2v_inst11.mult1_un40_sum_i_5 ));
    CascadeMux I__3043 (
            .O(N__20186),
            .I(\b2v_inst11.mult1_un40_sum_i_5_cascade_ ));
    InMux I__3042 (
            .O(N__20183),
            .I(N__20179));
    InMux I__3041 (
            .O(N__20182),
            .I(N__20176));
    LocalMux I__3040 (
            .O(N__20179),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ));
    LocalMux I__3039 (
            .O(N__20176),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ));
    InMux I__3038 (
            .O(N__20171),
            .I(N__20166));
    InMux I__3037 (
            .O(N__20170),
            .I(N__20163));
    InMux I__3036 (
            .O(N__20169),
            .I(N__20160));
    LocalMux I__3035 (
            .O(N__20166),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    LocalMux I__3034 (
            .O(N__20163),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    LocalMux I__3033 (
            .O(N__20160),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    CascadeMux I__3032 (
            .O(N__20153),
            .I(N__20150));
    InMux I__3031 (
            .O(N__20150),
            .I(N__20147));
    LocalMux I__3030 (
            .O(N__20147),
            .I(\b2v_inst11.un1_dutycycle_53_i_29 ));
    InMux I__3029 (
            .O(N__20144),
            .I(N__20141));
    LocalMux I__3028 (
            .O(N__20141),
            .I(N__20138));
    Span4Mux_v I__3027 (
            .O(N__20138),
            .I(N__20135));
    Span4Mux_v I__3026 (
            .O(N__20135),
            .I(N__20131));
    InMux I__3025 (
            .O(N__20134),
            .I(N__20128));
    Odrv4 I__3024 (
            .O(N__20131),
            .I(\b2v_inst16.count_rst ));
    LocalMux I__3023 (
            .O(N__20128),
            .I(\b2v_inst16.count_rst ));
    InMux I__3022 (
            .O(N__20123),
            .I(N__20120));
    LocalMux I__3021 (
            .O(N__20120),
            .I(N__20117));
    Span4Mux_h I__3020 (
            .O(N__20117),
            .I(N__20114));
    Span4Mux_v I__3019 (
            .O(N__20114),
            .I(N__20111));
    Odrv4 I__3018 (
            .O(N__20111),
            .I(\b2v_inst16.count_4_10 ));
    CEMux I__3017 (
            .O(N__20108),
            .I(N__20100));
    InMux I__3016 (
            .O(N__20107),
            .I(N__20097));
    CEMux I__3015 (
            .O(N__20106),
            .I(N__20090));
    InMux I__3014 (
            .O(N__20105),
            .I(N__20080));
    CEMux I__3013 (
            .O(N__20104),
            .I(N__20080));
    CEMux I__3012 (
            .O(N__20103),
            .I(N__20072));
    LocalMux I__3011 (
            .O(N__20100),
            .I(N__20069));
    LocalMux I__3010 (
            .O(N__20097),
            .I(N__20066));
    CEMux I__3009 (
            .O(N__20096),
            .I(N__20063));
    InMux I__3008 (
            .O(N__20095),
            .I(N__20056));
    InMux I__3007 (
            .O(N__20094),
            .I(N__20056));
    InMux I__3006 (
            .O(N__20093),
            .I(N__20056));
    LocalMux I__3005 (
            .O(N__20090),
            .I(N__20053));
    InMux I__3004 (
            .O(N__20089),
            .I(N__20050));
    InMux I__3003 (
            .O(N__20088),
            .I(N__20045));
    InMux I__3002 (
            .O(N__20087),
            .I(N__20045));
    InMux I__3001 (
            .O(N__20086),
            .I(N__20040));
    InMux I__3000 (
            .O(N__20085),
            .I(N__20040));
    LocalMux I__2999 (
            .O(N__20080),
            .I(N__20033));
    InMux I__2998 (
            .O(N__20079),
            .I(N__20022));
    CEMux I__2997 (
            .O(N__20078),
            .I(N__20022));
    InMux I__2996 (
            .O(N__20077),
            .I(N__20022));
    InMux I__2995 (
            .O(N__20076),
            .I(N__20022));
    InMux I__2994 (
            .O(N__20075),
            .I(N__20022));
    LocalMux I__2993 (
            .O(N__20072),
            .I(N__20019));
    Span4Mux_s1_v I__2992 (
            .O(N__20069),
            .I(N__20016));
    Span4Mux_v I__2991 (
            .O(N__20066),
            .I(N__20013));
    LocalMux I__2990 (
            .O(N__20063),
            .I(N__20008));
    LocalMux I__2989 (
            .O(N__20056),
            .I(N__20008));
    Span4Mux_s1_v I__2988 (
            .O(N__20053),
            .I(N__20003));
    LocalMux I__2987 (
            .O(N__20050),
            .I(N__20003));
    LocalMux I__2986 (
            .O(N__20045),
            .I(N__20000));
    LocalMux I__2985 (
            .O(N__20040),
            .I(N__19997));
    InMux I__2984 (
            .O(N__20039),
            .I(N__19988));
    CEMux I__2983 (
            .O(N__20038),
            .I(N__19988));
    InMux I__2982 (
            .O(N__20037),
            .I(N__19988));
    InMux I__2981 (
            .O(N__20036),
            .I(N__19988));
    Span4Mux_s3_h I__2980 (
            .O(N__20033),
            .I(N__19985));
    LocalMux I__2979 (
            .O(N__20022),
            .I(N__19982));
    Span4Mux_v I__2978 (
            .O(N__20019),
            .I(N__19965));
    Span4Mux_s1_h I__2977 (
            .O(N__20016),
            .I(N__19965));
    Span4Mux_v I__2976 (
            .O(N__20013),
            .I(N__19965));
    Span4Mux_s1_v I__2975 (
            .O(N__20008),
            .I(N__19965));
    Span4Mux_v I__2974 (
            .O(N__20003),
            .I(N__19965));
    Span4Mux_s1_v I__2973 (
            .O(N__20000),
            .I(N__19965));
    Span4Mux_s1_h I__2972 (
            .O(N__19997),
            .I(N__19965));
    LocalMux I__2971 (
            .O(N__19988),
            .I(N__19965));
    Odrv4 I__2970 (
            .O(N__19985),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__2969 (
            .O(N__19982),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__2968 (
            .O(N__19965),
            .I(\b2v_inst16.count_en ));
    InMux I__2967 (
            .O(N__19958),
            .I(N__19955));
    LocalMux I__2966 (
            .O(N__19955),
            .I(N__19951));
    InMux I__2965 (
            .O(N__19954),
            .I(N__19948));
    Sp12to4 I__2964 (
            .O(N__19951),
            .I(N__19943));
    LocalMux I__2963 (
            .O(N__19948),
            .I(N__19943));
    Span12Mux_s9_v I__2962 (
            .O(N__19943),
            .I(N__19940));
    Odrv12 I__2961 (
            .O(N__19940),
            .I(\b2v_inst16.countZ0Z_10 ));
    InMux I__2960 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__2959 (
            .O(N__19934),
            .I(N__19931));
    Span4Mux_s3_v I__2958 (
            .O(N__19931),
            .I(N__19928));
    Odrv4 I__2957 (
            .O(N__19928),
            .I(\b2v_inst11.mult1_un110_sum_i ));
    CascadeMux I__2956 (
            .O(N__19925),
            .I(N__19922));
    InMux I__2955 (
            .O(N__19922),
            .I(N__19919));
    LocalMux I__2954 (
            .O(N__19919),
            .I(\b2v_inst11.mult1_un117_sum_i_8 ));
    IoInMux I__2953 (
            .O(N__19916),
            .I(N__19913));
    LocalMux I__2952 (
            .O(N__19913),
            .I(N__19910));
    Odrv12 I__2951 (
            .O(N__19910),
            .I(vccst_en));
    InMux I__2950 (
            .O(N__19907),
            .I(N__19904));
    LocalMux I__2949 (
            .O(N__19904),
            .I(\b2v_inst11.un85_clk_100khz_4 ));
    CascadeMux I__2948 (
            .O(N__19901),
            .I(N__19898));
    InMux I__2947 (
            .O(N__19898),
            .I(N__19895));
    LocalMux I__2946 (
            .O(N__19895),
            .I(\b2v_inst11.mult1_un47_sum_cry_4_s ));
    InMux I__2945 (
            .O(N__19892),
            .I(\b2v_inst11.mult1_un47_sum_cry_3 ));
    InMux I__2944 (
            .O(N__19889),
            .I(N__19886));
    LocalMux I__2943 (
            .O(N__19886),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_s ));
    InMux I__2942 (
            .O(N__19883),
            .I(\b2v_inst11.mult1_un47_sum_cry_4 ));
    InMux I__2941 (
            .O(N__19880),
            .I(\b2v_inst11.mult1_un47_sum_cry_5 ));
    CascadeMux I__2940 (
            .O(N__19877),
            .I(N__19874));
    InMux I__2939 (
            .O(N__19874),
            .I(N__19871));
    LocalMux I__2938 (
            .O(N__19871),
            .I(\b2v_inst11.mult1_un47_sum_l_fx_6 ));
    CascadeMux I__2937 (
            .O(N__19868),
            .I(N__19865));
    InMux I__2936 (
            .O(N__19865),
            .I(N__19862));
    LocalMux I__2935 (
            .O(N__19862),
            .I(\b2v_inst11.mult1_un47_sum_i ));
    InMux I__2934 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__2933 (
            .O(N__19856),
            .I(N__19853));
    Odrv4 I__2932 (
            .O(N__19853),
            .I(\b2v_inst11.un1_dutycycle_53_axb_12 ));
    InMux I__2931 (
            .O(N__19850),
            .I(N__19847));
    LocalMux I__2930 (
            .O(N__19847),
            .I(N__19842));
    InMux I__2929 (
            .O(N__19846),
            .I(N__19835));
    InMux I__2928 (
            .O(N__19845),
            .I(N__19835));
    Span4Mux_h I__2927 (
            .O(N__19842),
            .I(N__19832));
    InMux I__2926 (
            .O(N__19841),
            .I(N__19827));
    InMux I__2925 (
            .O(N__19840),
            .I(N__19827));
    LocalMux I__2924 (
            .O(N__19835),
            .I(N__19824));
    Odrv4 I__2923 (
            .O(N__19832),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    LocalMux I__2922 (
            .O(N__19827),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    Odrv4 I__2921 (
            .O(N__19824),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    CascadeMux I__2920 (
            .O(N__19817),
            .I(N__19813));
    CascadeMux I__2919 (
            .O(N__19816),
            .I(N__19808));
    InMux I__2918 (
            .O(N__19813),
            .I(N__19805));
    InMux I__2917 (
            .O(N__19812),
            .I(N__19798));
    InMux I__2916 (
            .O(N__19811),
            .I(N__19798));
    InMux I__2915 (
            .O(N__19808),
            .I(N__19798));
    LocalMux I__2914 (
            .O(N__19805),
            .I(N__19795));
    LocalMux I__2913 (
            .O(N__19798),
            .I(N__19792));
    Odrv4 I__2912 (
            .O(N__19795),
            .I(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv4 I__2911 (
            .O(N__19792),
            .I(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    InMux I__2910 (
            .O(N__19787),
            .I(N__19784));
    LocalMux I__2909 (
            .O(N__19784),
            .I(N__19780));
    CascadeMux I__2908 (
            .O(N__19783),
            .I(N__19775));
    Span4Mux_v I__2907 (
            .O(N__19780),
            .I(N__19772));
    InMux I__2906 (
            .O(N__19779),
            .I(N__19767));
    InMux I__2905 (
            .O(N__19778),
            .I(N__19767));
    InMux I__2904 (
            .O(N__19775),
            .I(N__19764));
    Span4Mux_h I__2903 (
            .O(N__19772),
            .I(N__19759));
    LocalMux I__2902 (
            .O(N__19767),
            .I(N__19759));
    LocalMux I__2901 (
            .O(N__19764),
            .I(\b2v_inst11.count_RNIZ0Z_8 ));
    Odrv4 I__2900 (
            .O(N__19759),
            .I(\b2v_inst11.count_RNIZ0Z_8 ));
    InMux I__2899 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__2898 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_v I__2897 (
            .O(N__19748),
            .I(N__19745));
    Span4Mux_h I__2896 (
            .O(N__19745),
            .I(N__19742));
    Odrv4 I__2895 (
            .O(N__19742),
            .I(\b2v_inst11.curr_state_4_0 ));
    CascadeMux I__2894 (
            .O(N__19739),
            .I(N__19736));
    InMux I__2893 (
            .O(N__19736),
            .I(N__19733));
    LocalMux I__2892 (
            .O(N__19733),
            .I(\b2v_inst11.mult1_un47_sum_s_4_sf ));
    CascadeMux I__2891 (
            .O(N__19730),
            .I(N__19727));
    InMux I__2890 (
            .O(N__19727),
            .I(N__19724));
    LocalMux I__2889 (
            .O(N__19724),
            .I(\b2v_inst11.mult1_un40_sum_i_l_ofx_4 ));
    InMux I__2888 (
            .O(N__19721),
            .I(N__19718));
    LocalMux I__2887 (
            .O(N__19718),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ));
    InMux I__2886 (
            .O(N__19715),
            .I(N__19712));
    LocalMux I__2885 (
            .O(N__19712),
            .I(N__19709));
    Odrv4 I__2884 (
            .O(N__19709),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_7 ));
    CascadeMux I__2883 (
            .O(N__19706),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ));
    InMux I__2882 (
            .O(N__19703),
            .I(N__19700));
    LocalMux I__2881 (
            .O(N__19700),
            .I(\b2v_inst11.dutycycle_RNI_8Z0Z_6 ));
    InMux I__2880 (
            .O(N__19697),
            .I(N__19692));
    InMux I__2879 (
            .O(N__19696),
            .I(N__19687));
    InMux I__2878 (
            .O(N__19695),
            .I(N__19687));
    LocalMux I__2877 (
            .O(N__19692),
            .I(\b2v_inst11.mult1_un47_sum_cry_3_s ));
    LocalMux I__2876 (
            .O(N__19687),
            .I(\b2v_inst11.mult1_un47_sum_cry_3_s ));
    InMux I__2875 (
            .O(N__19682),
            .I(\b2v_inst11.mult1_un47_sum_cry_2 ));
    CascadeMux I__2874 (
            .O(N__19679),
            .I(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_9_cascade_ ));
    InMux I__2873 (
            .O(N__19676),
            .I(N__19672));
    InMux I__2872 (
            .O(N__19675),
            .I(N__19669));
    LocalMux I__2871 (
            .O(N__19672),
            .I(\b2v_inst11.dutycycleZ1Z_9 ));
    LocalMux I__2870 (
            .O(N__19669),
            .I(\b2v_inst11.dutycycleZ1Z_9 ));
    CascadeMux I__2869 (
            .O(N__19664),
            .I(\b2v_inst11.un1_dutycycle_53_30_a1_0_cascade_ ));
    InMux I__2868 (
            .O(N__19661),
            .I(N__19658));
    LocalMux I__2867 (
            .O(N__19658),
            .I(\b2v_inst11.un1_dutycycle_53_44_2 ));
    CascadeMux I__2866 (
            .O(N__19655),
            .I(\b2v_inst11.un1_dutycycle_53_5_1_cascade_ ));
    InMux I__2865 (
            .O(N__19652),
            .I(N__19645));
    InMux I__2864 (
            .O(N__19651),
            .I(N__19645));
    InMux I__2863 (
            .O(N__19650),
            .I(N__19642));
    LocalMux I__2862 (
            .O(N__19645),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_6 ));
    LocalMux I__2861 (
            .O(N__19642),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_6 ));
    InMux I__2860 (
            .O(N__19637),
            .I(N__19633));
    InMux I__2859 (
            .O(N__19636),
            .I(N__19630));
    LocalMux I__2858 (
            .O(N__19633),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_4 ));
    LocalMux I__2857 (
            .O(N__19630),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_4 ));
    InMux I__2856 (
            .O(N__19625),
            .I(N__19622));
    LocalMux I__2855 (
            .O(N__19622),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_8 ));
    CascadeMux I__2854 (
            .O(N__19619),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_8_cascade_ ));
    InMux I__2853 (
            .O(N__19616),
            .I(N__19613));
    LocalMux I__2852 (
            .O(N__19613),
            .I(\b2v_inst11.un1_dutycycle_53_9_1 ));
    InMux I__2851 (
            .O(N__19610),
            .I(N__19607));
    LocalMux I__2850 (
            .O(N__19607),
            .I(\b2v_inst11.un1_dutycycle_53_axb_7 ));
    InMux I__2849 (
            .O(N__19604),
            .I(N__19601));
    LocalMux I__2848 (
            .O(N__19601),
            .I(\b2v_inst20.un4_counter_6_and ));
    InMux I__2847 (
            .O(N__19598),
            .I(N__19595));
    LocalMux I__2846 (
            .O(N__19595),
            .I(\b2v_inst11.un1_dutycycle_53_39_d_0_0 ));
    CascadeMux I__2845 (
            .O(N__19592),
            .I(\b2v_inst11.dutycycle_RNITSFK3Z0Z_10_cascade_ ));
    CascadeMux I__2844 (
            .O(N__19589),
            .I(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_10_cascade_ ));
    InMux I__2843 (
            .O(N__19586),
            .I(N__19583));
    LocalMux I__2842 (
            .O(N__19583),
            .I(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_10 ));
    CascadeMux I__2841 (
            .O(N__19580),
            .I(N__19577));
    InMux I__2840 (
            .O(N__19577),
            .I(N__19571));
    InMux I__2839 (
            .O(N__19576),
            .I(N__19571));
    LocalMux I__2838 (
            .O(N__19571),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    CascadeMux I__2837 (
            .O(N__19568),
            .I(\b2v_inst11.dutycycleZ0Z_1_cascade_ ));
    CascadeMux I__2836 (
            .O(N__19565),
            .I(\b2v_inst11.dutycycle_RNITSFK3Z0Z_9_cascade_ ));
    CascadeMux I__2835 (
            .O(N__19562),
            .I(N__19559));
    InMux I__2834 (
            .O(N__19559),
            .I(N__19556));
    LocalMux I__2833 (
            .O(N__19556),
            .I(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_9 ));
    InMux I__2832 (
            .O(N__19553),
            .I(N__19550));
    LocalMux I__2831 (
            .O(N__19550),
            .I(\b2v_inst20.un4_counter_4_and ));
    InMux I__2830 (
            .O(N__19547),
            .I(N__19544));
    LocalMux I__2829 (
            .O(N__19544),
            .I(\b2v_inst20.un4_counter_5_and ));
    InMux I__2828 (
            .O(N__19541),
            .I(bfn_5_5_0_));
    InMux I__2827 (
            .O(N__19538),
            .I(N__19534));
    InMux I__2826 (
            .O(N__19537),
            .I(N__19531));
    LocalMux I__2825 (
            .O(N__19534),
            .I(\b2v_inst11.un1_dutycycle_53_axb_11_1 ));
    LocalMux I__2824 (
            .O(N__19531),
            .I(\b2v_inst11.un1_dutycycle_53_axb_11_1 ));
    CascadeMux I__2823 (
            .O(N__19526),
            .I(\b2v_inst11.un1_dutycycle_53_39_0_1_0_cascade_ ));
    CascadeMux I__2822 (
            .O(N__19523),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_ ));
    InMux I__2821 (
            .O(N__19520),
            .I(N__19516));
    InMux I__2820 (
            .O(N__19519),
            .I(N__19513));
    LocalMux I__2819 (
            .O(N__19516),
            .I(N__19510));
    LocalMux I__2818 (
            .O(N__19513),
            .I(N__19507));
    Span4Mux_h I__2817 (
            .O(N__19510),
            .I(N__19504));
    Span4Mux_v I__2816 (
            .O(N__19507),
            .I(N__19501));
    Odrv4 I__2815 (
            .O(N__19504),
            .I(\b2v_inst16.curr_state_2_0 ));
    Odrv4 I__2814 (
            .O(N__19501),
            .I(\b2v_inst16.curr_state_2_0 ));
    InMux I__2813 (
            .O(N__19496),
            .I(N__19493));
    LocalMux I__2812 (
            .O(N__19493),
            .I(\b2v_inst20.un4_counter_2_and ));
    InMux I__2811 (
            .O(N__19490),
            .I(N__19487));
    LocalMux I__2810 (
            .O(N__19487),
            .I(\b2v_inst20.un4_counter_3_and ));
    InMux I__2809 (
            .O(N__19484),
            .I(N__19476));
    InMux I__2808 (
            .O(N__19483),
            .I(N__19476));
    InMux I__2807 (
            .O(N__19482),
            .I(N__19471));
    InMux I__2806 (
            .O(N__19481),
            .I(N__19471));
    LocalMux I__2805 (
            .O(N__19476),
            .I(N_411));
    LocalMux I__2804 (
            .O(N__19471),
            .I(N_411));
    CascadeMux I__2803 (
            .O(N__19466),
            .I(\b2v_inst200.m6_i_0_cascade_ ));
    InMux I__2802 (
            .O(N__19463),
            .I(N__19458));
    InMux I__2801 (
            .O(N__19462),
            .I(N__19455));
    InMux I__2800 (
            .O(N__19461),
            .I(N__19452));
    LocalMux I__2799 (
            .O(N__19458),
            .I(N__19447));
    LocalMux I__2798 (
            .O(N__19455),
            .I(N__19447));
    LocalMux I__2797 (
            .O(N__19452),
            .I(N__19442));
    Span4Mux_h I__2796 (
            .O(N__19447),
            .I(N__19434));
    InMux I__2795 (
            .O(N__19446),
            .I(N__19429));
    InMux I__2794 (
            .O(N__19445),
            .I(N__19429));
    Span12Mux_s5_v I__2793 (
            .O(N__19442),
            .I(N__19426));
    InMux I__2792 (
            .O(N__19441),
            .I(N__19423));
    InMux I__2791 (
            .O(N__19440),
            .I(N__19418));
    InMux I__2790 (
            .O(N__19439),
            .I(N__19418));
    InMux I__2789 (
            .O(N__19438),
            .I(N__19413));
    InMux I__2788 (
            .O(N__19437),
            .I(N__19413));
    Span4Mux_v I__2787 (
            .O(N__19434),
            .I(N__19408));
    LocalMux I__2786 (
            .O(N__19429),
            .I(N__19408));
    Odrv12 I__2785 (
            .O(N__19426),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    LocalMux I__2784 (
            .O(N__19423),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    LocalMux I__2783 (
            .O(N__19418),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    LocalMux I__2782 (
            .O(N__19413),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    Odrv4 I__2781 (
            .O(N__19408),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    InMux I__2780 (
            .O(N__19397),
            .I(N__19394));
    LocalMux I__2779 (
            .O(N__19394),
            .I(\b2v_inst200.curr_state_3_0 ));
    InMux I__2778 (
            .O(N__19391),
            .I(N__19388));
    LocalMux I__2777 (
            .O(N__19388),
            .I(\b2v_inst200.curr_stateZ0Z_2 ));
    CascadeMux I__2776 (
            .O(N__19385),
            .I(\b2v_inst200.i4_mux_cascade_ ));
    CascadeMux I__2775 (
            .O(N__19382),
            .I(\b2v_inst200.curr_state_i_2_cascade_ ));
    IoInMux I__2774 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__2773 (
            .O(N__19376),
            .I(N__19373));
    IoSpan4Mux I__2772 (
            .O(N__19373),
            .I(N__19370));
    Span4Mux_s0_h I__2771 (
            .O(N__19370),
            .I(N__19367));
    Span4Mux_h I__2770 (
            .O(N__19367),
            .I(N__19364));
    Odrv4 I__2769 (
            .O(N__19364),
            .I(hda_sdo_atp));
    InMux I__2768 (
            .O(N__19361),
            .I(N__19357));
    InMux I__2767 (
            .O(N__19360),
            .I(N__19354));
    LocalMux I__2766 (
            .O(N__19357),
            .I(\b2v_inst200.N_3031_i ));
    LocalMux I__2765 (
            .O(N__19354),
            .I(\b2v_inst200.N_3031_i ));
    CascadeMux I__2764 (
            .O(N__19349),
            .I(N__19345));
    InMux I__2763 (
            .O(N__19348),
            .I(N__19337));
    InMux I__2762 (
            .O(N__19345),
            .I(N__19337));
    InMux I__2761 (
            .O(N__19344),
            .I(N__19337));
    LocalMux I__2760 (
            .O(N__19337),
            .I(\b2v_inst200.N_205 ));
    InMux I__2759 (
            .O(N__19334),
            .I(N__19325));
    InMux I__2758 (
            .O(N__19333),
            .I(N__19325));
    InMux I__2757 (
            .O(N__19332),
            .I(N__19325));
    LocalMux I__2756 (
            .O(N__19325),
            .I(\b2v_inst200.curr_state_i_2 ));
    CascadeMux I__2755 (
            .O(N__19322),
            .I(\b2v_inst200.N_205_cascade_ ));
    InMux I__2754 (
            .O(N__19319),
            .I(N__19316));
    LocalMux I__2753 (
            .O(N__19316),
            .I(\b2v_inst200.HDA_SDO_ATP_0 ));
    InMux I__2752 (
            .O(N__19313),
            .I(N__19305));
    InMux I__2751 (
            .O(N__19312),
            .I(N__19305));
    InMux I__2750 (
            .O(N__19311),
            .I(N__19300));
    InMux I__2749 (
            .O(N__19310),
            .I(N__19300));
    LocalMux I__2748 (
            .O(N__19305),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    LocalMux I__2747 (
            .O(N__19300),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    CascadeMux I__2746 (
            .O(N__19295),
            .I(N__19291));
    InMux I__2745 (
            .O(N__19294),
            .I(N__19287));
    InMux I__2744 (
            .O(N__19291),
            .I(N__19284));
    InMux I__2743 (
            .O(N__19290),
            .I(N__19281));
    LocalMux I__2742 (
            .O(N__19287),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    LocalMux I__2741 (
            .O(N__19284),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    LocalMux I__2740 (
            .O(N__19281),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    CascadeMux I__2739 (
            .O(N__19274),
            .I(N__19268));
    CascadeMux I__2738 (
            .O(N__19273),
            .I(N__19265));
    InMux I__2737 (
            .O(N__19272),
            .I(N__19258));
    InMux I__2736 (
            .O(N__19271),
            .I(N__19258));
    InMux I__2735 (
            .O(N__19268),
            .I(N__19258));
    InMux I__2734 (
            .O(N__19265),
            .I(N__19255));
    LocalMux I__2733 (
            .O(N__19258),
            .I(\b2v_inst200.N_282 ));
    LocalMux I__2732 (
            .O(N__19255),
            .I(\b2v_inst200.N_282 ));
    InMux I__2731 (
            .O(N__19250),
            .I(N__19247));
    LocalMux I__2730 (
            .O(N__19247),
            .I(\b2v_inst200.curr_state_3_1 ));
    CascadeMux I__2729 (
            .O(N__19244),
            .I(N__19240));
    CascadeMux I__2728 (
            .O(N__19243),
            .I(N__19236));
    InMux I__2727 (
            .O(N__19240),
            .I(N__19229));
    InMux I__2726 (
            .O(N__19239),
            .I(N__19229));
    InMux I__2725 (
            .O(N__19236),
            .I(N__19229));
    LocalMux I__2724 (
            .O(N__19229),
            .I(G_2814));
    InMux I__2723 (
            .O(N__19226),
            .I(\b2v_inst11.mult1_un166_sum_cry_5 ));
    CascadeMux I__2722 (
            .O(N__19223),
            .I(N__19220));
    InMux I__2721 (
            .O(N__19220),
            .I(N__19217));
    LocalMux I__2720 (
            .O(N__19217),
            .I(N__19214));
    Odrv12 I__2719 (
            .O(N__19214),
            .I(\b2v_inst11.un85_clk_100khz_0 ));
    CascadeMux I__2718 (
            .O(N__19211),
            .I(\b2v_inst200.N_58_cascade_ ));
    CascadeMux I__2717 (
            .O(N__19208),
            .I(\b2v_inst200.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__2716 (
            .O(N__19205),
            .I(\b2v_inst200.curr_stateZ0Z_1_cascade_ ));
    InMux I__2715 (
            .O(N__19202),
            .I(N__19199));
    LocalMux I__2714 (
            .O(N__19199),
            .I(\b2v_inst200.N_56 ));
    CascadeMux I__2713 (
            .O(N__19196),
            .I(N__19193));
    InMux I__2712 (
            .O(N__19193),
            .I(N__19190));
    LocalMux I__2711 (
            .O(N__19190),
            .I(N__19187));
    Span4Mux_h I__2710 (
            .O(N__19187),
            .I(N__19184));
    Odrv4 I__2709 (
            .O(N__19184),
            .I(gpio_fpga_soc_1));
    InMux I__2708 (
            .O(N__19181),
            .I(N__19178));
    LocalMux I__2707 (
            .O(N__19178),
            .I(\b2v_inst200.m6_i_0 ));
    CascadeMux I__2706 (
            .O(N__19175),
            .I(N__19170));
    InMux I__2705 (
            .O(N__19174),
            .I(N__19166));
    InMux I__2704 (
            .O(N__19173),
            .I(N__19161));
    InMux I__2703 (
            .O(N__19170),
            .I(N__19161));
    InMux I__2702 (
            .O(N__19169),
            .I(N__19158));
    LocalMux I__2701 (
            .O(N__19166),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__2700 (
            .O(N__19161),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__2699 (
            .O(N__19158),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    CascadeMux I__2698 (
            .O(N__19151),
            .I(N__19148));
    InMux I__2697 (
            .O(N__19148),
            .I(N__19145));
    LocalMux I__2696 (
            .O(N__19145),
            .I(\b2v_inst11.mult1_un110_sum_cry_5_s ));
    InMux I__2695 (
            .O(N__19142),
            .I(\b2v_inst11.mult1_un117_sum_cry_5 ));
    InMux I__2694 (
            .O(N__19139),
            .I(N__19136));
    LocalMux I__2693 (
            .O(N__19136),
            .I(\b2v_inst11.mult1_un110_sum_cry_6_s ));
    CascadeMux I__2692 (
            .O(N__19133),
            .I(N__19129));
    CascadeMux I__2691 (
            .O(N__19132),
            .I(N__19125));
    InMux I__2690 (
            .O(N__19129),
            .I(N__19118));
    InMux I__2689 (
            .O(N__19128),
            .I(N__19118));
    InMux I__2688 (
            .O(N__19125),
            .I(N__19118));
    LocalMux I__2687 (
            .O(N__19118),
            .I(\b2v_inst11.mult1_un110_sum_i_0_8 ));
    InMux I__2686 (
            .O(N__19115),
            .I(\b2v_inst11.mult1_un117_sum_cry_6 ));
    CascadeMux I__2685 (
            .O(N__19112),
            .I(N__19109));
    InMux I__2684 (
            .O(N__19109),
            .I(N__19106));
    LocalMux I__2683 (
            .O(N__19106),
            .I(\b2v_inst11.mult1_un117_sum_axb_8 ));
    InMux I__2682 (
            .O(N__19103),
            .I(\b2v_inst11.mult1_un117_sum_cry_7 ));
    CascadeMux I__2681 (
            .O(N__19100),
            .I(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ));
    InMux I__2680 (
            .O(N__19097),
            .I(N__19094));
    LocalMux I__2679 (
            .O(N__19094),
            .I(N__19091));
    Span4Mux_v I__2678 (
            .O(N__19091),
            .I(N__19088));
    Odrv4 I__2677 (
            .O(N__19088),
            .I(\b2v_inst11.mult1_un103_sum_cry_4_s ));
    InMux I__2676 (
            .O(N__19085),
            .I(\b2v_inst11.mult1_un110_sum_cry_4 ));
    CascadeMux I__2675 (
            .O(N__19082),
            .I(N__19079));
    InMux I__2674 (
            .O(N__19079),
            .I(N__19076));
    LocalMux I__2673 (
            .O(N__19076),
            .I(N__19073));
    Span4Mux_v I__2672 (
            .O(N__19073),
            .I(N__19070));
    Odrv4 I__2671 (
            .O(N__19070),
            .I(\b2v_inst11.mult1_un103_sum_cry_5_s ));
    InMux I__2670 (
            .O(N__19067),
            .I(\b2v_inst11.mult1_un110_sum_cry_5 ));
    InMux I__2669 (
            .O(N__19064),
            .I(N__19061));
    LocalMux I__2668 (
            .O(N__19061),
            .I(N__19058));
    Span4Mux_h I__2667 (
            .O(N__19058),
            .I(N__19055));
    Odrv4 I__2666 (
            .O(N__19055),
            .I(\b2v_inst11.mult1_un103_sum_cry_6_s ));
    CascadeMux I__2665 (
            .O(N__19052),
            .I(N__19048));
    CascadeMux I__2664 (
            .O(N__19051),
            .I(N__19044));
    InMux I__2663 (
            .O(N__19048),
            .I(N__19037));
    InMux I__2662 (
            .O(N__19047),
            .I(N__19037));
    InMux I__2661 (
            .O(N__19044),
            .I(N__19037));
    LocalMux I__2660 (
            .O(N__19037),
            .I(\b2v_inst11.mult1_un103_sum_i_0_8 ));
    InMux I__2659 (
            .O(N__19034),
            .I(\b2v_inst11.mult1_un110_sum_cry_6 ));
    CascadeMux I__2658 (
            .O(N__19031),
            .I(N__19028));
    InMux I__2657 (
            .O(N__19028),
            .I(N__19025));
    LocalMux I__2656 (
            .O(N__19025),
            .I(N__19022));
    Span4Mux_h I__2655 (
            .O(N__19022),
            .I(N__19019));
    Odrv4 I__2654 (
            .O(N__19019),
            .I(\b2v_inst11.mult1_un110_sum_axb_8 ));
    InMux I__2653 (
            .O(N__19016),
            .I(\b2v_inst11.mult1_un110_sum_cry_7 ));
    CascadeMux I__2652 (
            .O(N__19013),
            .I(\b2v_inst11.mult1_un110_sum_s_8_cascade_ ));
    InMux I__2651 (
            .O(N__19010),
            .I(\b2v_inst11.mult1_un117_sum_cry_2 ));
    CascadeMux I__2650 (
            .O(N__19007),
            .I(N__19004));
    InMux I__2649 (
            .O(N__19004),
            .I(N__19001));
    LocalMux I__2648 (
            .O(N__19001),
            .I(\b2v_inst11.mult1_un110_sum_cry_3_s ));
    InMux I__2647 (
            .O(N__18998),
            .I(\b2v_inst11.mult1_un117_sum_cry_3 ));
    InMux I__2646 (
            .O(N__18995),
            .I(N__18992));
    LocalMux I__2645 (
            .O(N__18992),
            .I(\b2v_inst11.mult1_un110_sum_cry_4_s ));
    InMux I__2644 (
            .O(N__18989),
            .I(\b2v_inst11.mult1_un117_sum_cry_4 ));
    InMux I__2643 (
            .O(N__18986),
            .I(N__18983));
    LocalMux I__2642 (
            .O(N__18983),
            .I(N__18980));
    Odrv4 I__2641 (
            .O(N__18980),
            .I(\b2v_inst11.mult1_un68_sum_i_8 ));
    InMux I__2640 (
            .O(N__18977),
            .I(N__18974));
    LocalMux I__2639 (
            .O(N__18974),
            .I(N__18971));
    Span12Mux_s10_h I__2638 (
            .O(N__18971),
            .I(N__18966));
    InMux I__2637 (
            .O(N__18970),
            .I(N__18963));
    InMux I__2636 (
            .O(N__18969),
            .I(N__18960));
    Odrv12 I__2635 (
            .O(N__18966),
            .I(\b2v_inst11.countZ0Z_14 ));
    LocalMux I__2634 (
            .O(N__18963),
            .I(\b2v_inst11.countZ0Z_14 ));
    LocalMux I__2633 (
            .O(N__18960),
            .I(\b2v_inst11.countZ0Z_14 ));
    CascadeMux I__2632 (
            .O(N__18953),
            .I(N__18950));
    InMux I__2631 (
            .O(N__18950),
            .I(N__18947));
    LocalMux I__2630 (
            .O(N__18947),
            .I(N__18944));
    Odrv4 I__2629 (
            .O(N__18944),
            .I(\b2v_inst11.N_5994_i ));
    InMux I__2628 (
            .O(N__18941),
            .I(N__18938));
    LocalMux I__2627 (
            .O(N__18938),
            .I(N__18935));
    Span4Mux_h I__2626 (
            .O(N__18935),
            .I(N__18930));
    InMux I__2625 (
            .O(N__18934),
            .I(N__18927));
    InMux I__2624 (
            .O(N__18933),
            .I(N__18924));
    Odrv4 I__2623 (
            .O(N__18930),
            .I(\b2v_inst11.countZ0Z_15 ));
    LocalMux I__2622 (
            .O(N__18927),
            .I(\b2v_inst11.countZ0Z_15 ));
    LocalMux I__2621 (
            .O(N__18924),
            .I(\b2v_inst11.countZ0Z_15 ));
    InMux I__2620 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__2619 (
            .O(N__18914),
            .I(N__18911));
    Odrv4 I__2618 (
            .O(N__18911),
            .I(\b2v_inst11.mult1_un61_sum_i_8 ));
    CascadeMux I__2617 (
            .O(N__18908),
            .I(N__18905));
    InMux I__2616 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__2615 (
            .O(N__18902),
            .I(\b2v_inst11.N_5995_i ));
    InMux I__2614 (
            .O(N__18899),
            .I(bfn_4_13_0_));
    InMux I__2613 (
            .O(N__18896),
            .I(N__18893));
    LocalMux I__2612 (
            .O(N__18893),
            .I(\b2v_inst11.mult1_un110_sum_i_8 ));
    InMux I__2611 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__2610 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_v I__2609 (
            .O(N__18884),
            .I(N__18881));
    Odrv4 I__2608 (
            .O(N__18881),
            .I(\b2v_inst11.mult1_un103_sum_i ));
    InMux I__2607 (
            .O(N__18878),
            .I(\b2v_inst11.mult1_un110_sum_cry_2 ));
    CascadeMux I__2606 (
            .O(N__18875),
            .I(N__18872));
    InMux I__2605 (
            .O(N__18872),
            .I(N__18869));
    LocalMux I__2604 (
            .O(N__18869),
            .I(N__18866));
    Span4Mux_h I__2603 (
            .O(N__18866),
            .I(N__18863));
    Odrv4 I__2602 (
            .O(N__18863),
            .I(\b2v_inst11.mult1_un103_sum_cry_3_s ));
    InMux I__2601 (
            .O(N__18860),
            .I(\b2v_inst11.mult1_un110_sum_cry_3 ));
    InMux I__2600 (
            .O(N__18857),
            .I(N__18854));
    LocalMux I__2599 (
            .O(N__18854),
            .I(N__18851));
    Span4Mux_h I__2598 (
            .O(N__18851),
            .I(N__18848));
    Span4Mux_v I__2597 (
            .O(N__18848),
            .I(N__18843));
    InMux I__2596 (
            .O(N__18847),
            .I(N__18840));
    InMux I__2595 (
            .O(N__18846),
            .I(N__18837));
    Odrv4 I__2594 (
            .O(N__18843),
            .I(\b2v_inst11.countZ0Z_6 ));
    LocalMux I__2593 (
            .O(N__18840),
            .I(\b2v_inst11.countZ0Z_6 ));
    LocalMux I__2592 (
            .O(N__18837),
            .I(\b2v_inst11.countZ0Z_6 ));
    InMux I__2591 (
            .O(N__18830),
            .I(N__18827));
    LocalMux I__2590 (
            .O(N__18827),
            .I(\b2v_inst11.N_5986_i ));
    InMux I__2589 (
            .O(N__18824),
            .I(N__18821));
    LocalMux I__2588 (
            .O(N__18821),
            .I(N__18818));
    Span4Mux_v I__2587 (
            .O(N__18818),
            .I(N__18815));
    Span4Mux_v I__2586 (
            .O(N__18815),
            .I(N__18810));
    InMux I__2585 (
            .O(N__18814),
            .I(N__18807));
    InMux I__2584 (
            .O(N__18813),
            .I(N__18804));
    Odrv4 I__2583 (
            .O(N__18810),
            .I(\b2v_inst11.countZ0Z_7 ));
    LocalMux I__2582 (
            .O(N__18807),
            .I(\b2v_inst11.countZ0Z_7 ));
    LocalMux I__2581 (
            .O(N__18804),
            .I(\b2v_inst11.countZ0Z_7 ));
    InMux I__2580 (
            .O(N__18797),
            .I(N__18794));
    LocalMux I__2579 (
            .O(N__18794),
            .I(\b2v_inst11.N_5987_i ));
    InMux I__2578 (
            .O(N__18791),
            .I(N__18788));
    LocalMux I__2577 (
            .O(N__18788),
            .I(N__18783));
    InMux I__2576 (
            .O(N__18787),
            .I(N__18780));
    InMux I__2575 (
            .O(N__18786),
            .I(N__18777));
    Span4Mux_v I__2574 (
            .O(N__18783),
            .I(N__18774));
    LocalMux I__2573 (
            .O(N__18780),
            .I(N__18771));
    LocalMux I__2572 (
            .O(N__18777),
            .I(N__18768));
    Odrv4 I__2571 (
            .O(N__18774),
            .I(\b2v_inst11.countZ0Z_8 ));
    Odrv4 I__2570 (
            .O(N__18771),
            .I(\b2v_inst11.countZ0Z_8 ));
    Odrv4 I__2569 (
            .O(N__18768),
            .I(\b2v_inst11.countZ0Z_8 ));
    CascadeMux I__2568 (
            .O(N__18761),
            .I(N__18758));
    InMux I__2567 (
            .O(N__18758),
            .I(N__18755));
    LocalMux I__2566 (
            .O(N__18755),
            .I(\b2v_inst11.N_5988_i ));
    InMux I__2565 (
            .O(N__18752),
            .I(N__18749));
    LocalMux I__2564 (
            .O(N__18749),
            .I(N__18744));
    InMux I__2563 (
            .O(N__18748),
            .I(N__18741));
    InMux I__2562 (
            .O(N__18747),
            .I(N__18738));
    Span4Mux_h I__2561 (
            .O(N__18744),
            .I(N__18731));
    LocalMux I__2560 (
            .O(N__18741),
            .I(N__18731));
    LocalMux I__2559 (
            .O(N__18738),
            .I(N__18731));
    Odrv4 I__2558 (
            .O(N__18731),
            .I(\b2v_inst11.countZ0Z_9 ));
    CascadeMux I__2557 (
            .O(N__18728),
            .I(N__18725));
    InMux I__2556 (
            .O(N__18725),
            .I(N__18722));
    LocalMux I__2555 (
            .O(N__18722),
            .I(\b2v_inst11.N_5989_i ));
    InMux I__2554 (
            .O(N__18719),
            .I(N__18716));
    LocalMux I__2553 (
            .O(N__18716),
            .I(N__18713));
    Span4Mux_h I__2552 (
            .O(N__18713),
            .I(N__18710));
    Odrv4 I__2551 (
            .O(N__18710),
            .I(\b2v_inst11.mult1_un96_sum_i_8 ));
    InMux I__2550 (
            .O(N__18707),
            .I(N__18704));
    LocalMux I__2549 (
            .O(N__18704),
            .I(N__18700));
    InMux I__2548 (
            .O(N__18703),
            .I(N__18696));
    Span4Mux_h I__2547 (
            .O(N__18700),
            .I(N__18693));
    InMux I__2546 (
            .O(N__18699),
            .I(N__18690));
    LocalMux I__2545 (
            .O(N__18696),
            .I(N__18687));
    Span4Mux_s0_h I__2544 (
            .O(N__18693),
            .I(N__18682));
    LocalMux I__2543 (
            .O(N__18690),
            .I(N__18682));
    Odrv4 I__2542 (
            .O(N__18687),
            .I(\b2v_inst11.countZ0Z_10 ));
    Odrv4 I__2541 (
            .O(N__18682),
            .I(\b2v_inst11.countZ0Z_10 ));
    CascadeMux I__2540 (
            .O(N__18677),
            .I(N__18674));
    InMux I__2539 (
            .O(N__18674),
            .I(N__18671));
    LocalMux I__2538 (
            .O(N__18671),
            .I(\b2v_inst11.N_5990_i ));
    InMux I__2537 (
            .O(N__18668),
            .I(N__18665));
    LocalMux I__2536 (
            .O(N__18665),
            .I(N__18662));
    Odrv4 I__2535 (
            .O(N__18662),
            .I(\b2v_inst11.mult1_un89_sum_i_8 ));
    InMux I__2534 (
            .O(N__18659),
            .I(N__18655));
    InMux I__2533 (
            .O(N__18658),
            .I(N__18652));
    LocalMux I__2532 (
            .O(N__18655),
            .I(N__18648));
    LocalMux I__2531 (
            .O(N__18652),
            .I(N__18645));
    InMux I__2530 (
            .O(N__18651),
            .I(N__18642));
    Span4Mux_s3_v I__2529 (
            .O(N__18648),
            .I(N__18639));
    Span4Mux_h I__2528 (
            .O(N__18645),
            .I(N__18634));
    LocalMux I__2527 (
            .O(N__18642),
            .I(N__18634));
    Odrv4 I__2526 (
            .O(N__18639),
            .I(\b2v_inst11.countZ0Z_11 ));
    Odrv4 I__2525 (
            .O(N__18634),
            .I(\b2v_inst11.countZ0Z_11 ));
    CascadeMux I__2524 (
            .O(N__18629),
            .I(N__18626));
    InMux I__2523 (
            .O(N__18626),
            .I(N__18623));
    LocalMux I__2522 (
            .O(N__18623),
            .I(\b2v_inst11.N_5991_i ));
    InMux I__2521 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__2520 (
            .O(N__18617),
            .I(N__18612));
    CascadeMux I__2519 (
            .O(N__18616),
            .I(N__18609));
    InMux I__2518 (
            .O(N__18615),
            .I(N__18606));
    Span4Mux_v I__2517 (
            .O(N__18612),
            .I(N__18603));
    InMux I__2516 (
            .O(N__18609),
            .I(N__18600));
    LocalMux I__2515 (
            .O(N__18606),
            .I(N__18597));
    Odrv4 I__2514 (
            .O(N__18603),
            .I(\b2v_inst11.countZ0Z_12 ));
    LocalMux I__2513 (
            .O(N__18600),
            .I(\b2v_inst11.countZ0Z_12 ));
    Odrv4 I__2512 (
            .O(N__18597),
            .I(\b2v_inst11.countZ0Z_12 ));
    InMux I__2511 (
            .O(N__18590),
            .I(N__18587));
    LocalMux I__2510 (
            .O(N__18587),
            .I(N__18584));
    Span4Mux_h I__2509 (
            .O(N__18584),
            .I(N__18581));
    Odrv4 I__2508 (
            .O(N__18581),
            .I(\b2v_inst11.mult1_un82_sum_i_8 ));
    CascadeMux I__2507 (
            .O(N__18578),
            .I(N__18575));
    InMux I__2506 (
            .O(N__18575),
            .I(N__18572));
    LocalMux I__2505 (
            .O(N__18572),
            .I(\b2v_inst11.N_5992_i ));
    InMux I__2504 (
            .O(N__18569),
            .I(N__18566));
    LocalMux I__2503 (
            .O(N__18566),
            .I(N__18563));
    Span4Mux_h I__2502 (
            .O(N__18563),
            .I(N__18560));
    Odrv4 I__2501 (
            .O(N__18560),
            .I(\b2v_inst11.mult1_un75_sum_i_8 ));
    InMux I__2500 (
            .O(N__18557),
            .I(N__18553));
    InMux I__2499 (
            .O(N__18556),
            .I(N__18550));
    LocalMux I__2498 (
            .O(N__18553),
            .I(N__18547));
    LocalMux I__2497 (
            .O(N__18550),
            .I(N__18544));
    Span4Mux_v I__2496 (
            .O(N__18547),
            .I(N__18538));
    Span4Mux_s2_v I__2495 (
            .O(N__18544),
            .I(N__18538));
    InMux I__2494 (
            .O(N__18543),
            .I(N__18535));
    Odrv4 I__2493 (
            .O(N__18538),
            .I(\b2v_inst11.countZ0Z_13 ));
    LocalMux I__2492 (
            .O(N__18535),
            .I(\b2v_inst11.countZ0Z_13 ));
    CascadeMux I__2491 (
            .O(N__18530),
            .I(N__18527));
    InMux I__2490 (
            .O(N__18527),
            .I(N__18524));
    LocalMux I__2489 (
            .O(N__18524),
            .I(\b2v_inst11.N_5993_i ));
    InMux I__2488 (
            .O(N__18521),
            .I(N__18518));
    LocalMux I__2487 (
            .O(N__18518),
            .I(N__18515));
    Odrv12 I__2486 (
            .O(N__18515),
            .I(\b2v_inst11.mult1_un75_sum_i ));
    InMux I__2485 (
            .O(N__18512),
            .I(N__18509));
    LocalMux I__2484 (
            .O(N__18509),
            .I(N__18505));
    CascadeMux I__2483 (
            .O(N__18508),
            .I(N__18501));
    Span4Mux_h I__2482 (
            .O(N__18505),
            .I(N__18497));
    InMux I__2481 (
            .O(N__18504),
            .I(N__18492));
    InMux I__2480 (
            .O(N__18501),
            .I(N__18492));
    InMux I__2479 (
            .O(N__18500),
            .I(N__18489));
    Odrv4 I__2478 (
            .O(N__18497),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__2477 (
            .O(N__18492),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__2476 (
            .O(N__18489),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    InMux I__2475 (
            .O(N__18482),
            .I(N__18479));
    LocalMux I__2474 (
            .O(N__18479),
            .I(N__18475));
    InMux I__2473 (
            .O(N__18478),
            .I(N__18468));
    Span4Mux_v I__2472 (
            .O(N__18475),
            .I(N__18465));
    InMux I__2471 (
            .O(N__18474),
            .I(N__18462));
    InMux I__2470 (
            .O(N__18473),
            .I(N__18455));
    InMux I__2469 (
            .O(N__18472),
            .I(N__18455));
    InMux I__2468 (
            .O(N__18471),
            .I(N__18455));
    LocalMux I__2467 (
            .O(N__18468),
            .I(N__18452));
    Odrv4 I__2466 (
            .O(N__18465),
            .I(\b2v_inst11.countZ0Z_0 ));
    LocalMux I__2465 (
            .O(N__18462),
            .I(\b2v_inst11.countZ0Z_0 ));
    LocalMux I__2464 (
            .O(N__18455),
            .I(\b2v_inst11.countZ0Z_0 ));
    Odrv4 I__2463 (
            .O(N__18452),
            .I(\b2v_inst11.countZ0Z_0 ));
    InMux I__2462 (
            .O(N__18443),
            .I(N__18440));
    LocalMux I__2461 (
            .O(N__18440),
            .I(\b2v_inst11.N_5980_i ));
    InMux I__2460 (
            .O(N__18437),
            .I(N__18434));
    LocalMux I__2459 (
            .O(N__18434),
            .I(N__18429));
    CascadeMux I__2458 (
            .O(N__18433),
            .I(N__18426));
    InMux I__2457 (
            .O(N__18432),
            .I(N__18423));
    Span4Mux_v I__2456 (
            .O(N__18429),
            .I(N__18420));
    InMux I__2455 (
            .O(N__18426),
            .I(N__18417));
    LocalMux I__2454 (
            .O(N__18423),
            .I(N__18414));
    Odrv4 I__2453 (
            .O(N__18420),
            .I(\b2v_inst11.countZ0Z_1 ));
    LocalMux I__2452 (
            .O(N__18417),
            .I(\b2v_inst11.countZ0Z_1 ));
    Odrv4 I__2451 (
            .O(N__18414),
            .I(\b2v_inst11.countZ0Z_1 ));
    InMux I__2450 (
            .O(N__18407),
            .I(N__18404));
    LocalMux I__2449 (
            .O(N__18404),
            .I(\b2v_inst11.N_5981_i ));
    InMux I__2448 (
            .O(N__18401),
            .I(N__18398));
    LocalMux I__2447 (
            .O(N__18398),
            .I(N__18395));
    Span4Mux_v I__2446 (
            .O(N__18395),
            .I(N__18391));
    CascadeMux I__2445 (
            .O(N__18394),
            .I(N__18388));
    Span4Mux_h I__2444 (
            .O(N__18391),
            .I(N__18384));
    InMux I__2443 (
            .O(N__18388),
            .I(N__18381));
    InMux I__2442 (
            .O(N__18387),
            .I(N__18378));
    Odrv4 I__2441 (
            .O(N__18384),
            .I(\b2v_inst11.countZ0Z_2 ));
    LocalMux I__2440 (
            .O(N__18381),
            .I(\b2v_inst11.countZ0Z_2 ));
    LocalMux I__2439 (
            .O(N__18378),
            .I(\b2v_inst11.countZ0Z_2 ));
    CascadeMux I__2438 (
            .O(N__18371),
            .I(N__18368));
    InMux I__2437 (
            .O(N__18368),
            .I(N__18365));
    LocalMux I__2436 (
            .O(N__18365),
            .I(\b2v_inst11.N_5982_i ));
    InMux I__2435 (
            .O(N__18362),
            .I(N__18359));
    LocalMux I__2434 (
            .O(N__18359),
            .I(N__18355));
    CascadeMux I__2433 (
            .O(N__18358),
            .I(N__18351));
    Span4Mux_v I__2432 (
            .O(N__18355),
            .I(N__18348));
    InMux I__2431 (
            .O(N__18354),
            .I(N__18345));
    InMux I__2430 (
            .O(N__18351),
            .I(N__18342));
    Odrv4 I__2429 (
            .O(N__18348),
            .I(\b2v_inst11.countZ0Z_3 ));
    LocalMux I__2428 (
            .O(N__18345),
            .I(\b2v_inst11.countZ0Z_3 ));
    LocalMux I__2427 (
            .O(N__18342),
            .I(\b2v_inst11.countZ0Z_3 ));
    CascadeMux I__2426 (
            .O(N__18335),
            .I(N__18332));
    InMux I__2425 (
            .O(N__18332),
            .I(N__18329));
    LocalMux I__2424 (
            .O(N__18329),
            .I(\b2v_inst11.N_5983_i ));
    InMux I__2423 (
            .O(N__18326),
            .I(N__18323));
    LocalMux I__2422 (
            .O(N__18323),
            .I(N__18320));
    Span4Mux_v I__2421 (
            .O(N__18320),
            .I(N__18315));
    InMux I__2420 (
            .O(N__18319),
            .I(N__18312));
    InMux I__2419 (
            .O(N__18318),
            .I(N__18309));
    Odrv4 I__2418 (
            .O(N__18315),
            .I(\b2v_inst11.countZ0Z_4 ));
    LocalMux I__2417 (
            .O(N__18312),
            .I(\b2v_inst11.countZ0Z_4 ));
    LocalMux I__2416 (
            .O(N__18309),
            .I(\b2v_inst11.countZ0Z_4 ));
    CascadeMux I__2415 (
            .O(N__18302),
            .I(N__18299));
    InMux I__2414 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__2413 (
            .O(N__18296),
            .I(\b2v_inst11.N_5984_i ));
    InMux I__2412 (
            .O(N__18293),
            .I(N__18290));
    LocalMux I__2411 (
            .O(N__18290),
            .I(N__18287));
    Span4Mux_v I__2410 (
            .O(N__18287),
            .I(N__18282));
    InMux I__2409 (
            .O(N__18286),
            .I(N__18279));
    InMux I__2408 (
            .O(N__18285),
            .I(N__18276));
    Odrv4 I__2407 (
            .O(N__18282),
            .I(\b2v_inst11.countZ0Z_5 ));
    LocalMux I__2406 (
            .O(N__18279),
            .I(\b2v_inst11.countZ0Z_5 ));
    LocalMux I__2405 (
            .O(N__18276),
            .I(\b2v_inst11.countZ0Z_5 ));
    CascadeMux I__2404 (
            .O(N__18269),
            .I(N__18266));
    InMux I__2403 (
            .O(N__18266),
            .I(N__18263));
    LocalMux I__2402 (
            .O(N__18263),
            .I(\b2v_inst11.N_5985_i ));
    InMux I__2401 (
            .O(N__18260),
            .I(N__18257));
    LocalMux I__2400 (
            .O(N__18257),
            .I(N__18254));
    Odrv4 I__2399 (
            .O(N__18254),
            .I(\b2v_inst11.mult1_un61_sum_axb_8 ));
    InMux I__2398 (
            .O(N__18251),
            .I(\b2v_inst11.mult1_un54_sum_cry_6 ));
    InMux I__2397 (
            .O(N__18248),
            .I(\b2v_inst11.mult1_un54_sum_cry_7 ));
    CascadeMux I__2396 (
            .O(N__18245),
            .I(N__18240));
    InMux I__2395 (
            .O(N__18244),
            .I(N__18237));
    InMux I__2394 (
            .O(N__18243),
            .I(N__18232));
    InMux I__2393 (
            .O(N__18240),
            .I(N__18232));
    LocalMux I__2392 (
            .O(N__18237),
            .I(N__18228));
    LocalMux I__2391 (
            .O(N__18232),
            .I(N__18225));
    InMux I__2390 (
            .O(N__18231),
            .I(N__18222));
    Span4Mux_s3_h I__2389 (
            .O(N__18228),
            .I(N__18219));
    Odrv4 I__2388 (
            .O(N__18225),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    LocalMux I__2387 (
            .O(N__18222),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    Odrv4 I__2386 (
            .O(N__18219),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    CascadeMux I__2385 (
            .O(N__18212),
            .I(N__18209));
    InMux I__2384 (
            .O(N__18209),
            .I(N__18206));
    LocalMux I__2383 (
            .O(N__18206),
            .I(\b2v_inst11.mult1_un47_sum_l_fx_3 ));
    InMux I__2382 (
            .O(N__18203),
            .I(N__18200));
    LocalMux I__2381 (
            .O(N__18200),
            .I(N__18197));
    Span4Mux_v I__2380 (
            .O(N__18197),
            .I(N__18194));
    Odrv4 I__2379 (
            .O(N__18194),
            .I(vpp_ok));
    IoInMux I__2378 (
            .O(N__18191),
            .I(N__18188));
    LocalMux I__2377 (
            .O(N__18188),
            .I(N__18185));
    IoSpan4Mux I__2376 (
            .O(N__18185),
            .I(N__18182));
    Span4Mux_s1_h I__2375 (
            .O(N__18182),
            .I(N__18179));
    Span4Mux_v I__2374 (
            .O(N__18179),
            .I(N__18176));
    Odrv4 I__2373 (
            .O(N__18176),
            .I(vddq_en));
    InMux I__2372 (
            .O(N__18173),
            .I(N__18170));
    LocalMux I__2371 (
            .O(N__18170),
            .I(N__18167));
    Span4Mux_s3_h I__2370 (
            .O(N__18167),
            .I(N__18164));
    Odrv4 I__2369 (
            .O(N__18164),
            .I(\b2v_inst11.mult1_un54_sum_i ));
    InMux I__2368 (
            .O(N__18161),
            .I(N__18158));
    LocalMux I__2367 (
            .O(N__18158),
            .I(N__18154));
    CascadeMux I__2366 (
            .O(N__18157),
            .I(N__18150));
    Span4Mux_h I__2365 (
            .O(N__18154),
            .I(N__18146));
    InMux I__2364 (
            .O(N__18153),
            .I(N__18141));
    InMux I__2363 (
            .O(N__18150),
            .I(N__18141));
    InMux I__2362 (
            .O(N__18149),
            .I(N__18138));
    Odrv4 I__2361 (
            .O(N__18146),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__2360 (
            .O(N__18141),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__2359 (
            .O(N__18138),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    InMux I__2358 (
            .O(N__18131),
            .I(N__18128));
    LocalMux I__2357 (
            .O(N__18128),
            .I(N__18125));
    Span4Mux_s3_h I__2356 (
            .O(N__18125),
            .I(N__18122));
    Odrv4 I__2355 (
            .O(N__18122),
            .I(\b2v_inst11.mult1_un61_sum_i ));
    CascadeMux I__2354 (
            .O(N__18119),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_6_cascade_ ));
    InMux I__2353 (
            .O(N__18116),
            .I(N__18113));
    LocalMux I__2352 (
            .O(N__18113),
            .I(\b2v_inst11.dutycycle_RNI_9Z0Z_7 ));
    CascadeMux I__2351 (
            .O(N__18110),
            .I(\b2v_inst11.un1_dutycycle_53_46_0_cascade_ ));
    InMux I__2350 (
            .O(N__18107),
            .I(N__18104));
    LocalMux I__2349 (
            .O(N__18104),
            .I(N__18101));
    Odrv4 I__2348 (
            .O(N__18101),
            .I(\b2v_inst11.un1_dutycycle_53_axb_11_1_0 ));
    CascadeMux I__2347 (
            .O(N__18098),
            .I(N__18095));
    InMux I__2346 (
            .O(N__18095),
            .I(N__18092));
    LocalMux I__2345 (
            .O(N__18092),
            .I(N__18089));
    Odrv4 I__2344 (
            .O(N__18089),
            .I(\b2v_inst11.mult1_un54_sum_cry_3_s ));
    InMux I__2343 (
            .O(N__18086),
            .I(\b2v_inst11.mult1_un54_sum_cry_2 ));
    InMux I__2342 (
            .O(N__18083),
            .I(N__18080));
    LocalMux I__2341 (
            .O(N__18080),
            .I(N__18077));
    Odrv4 I__2340 (
            .O(N__18077),
            .I(\b2v_inst11.mult1_un54_sum_cry_4_s ));
    InMux I__2339 (
            .O(N__18074),
            .I(\b2v_inst11.mult1_un54_sum_cry_3 ));
    CascadeMux I__2338 (
            .O(N__18071),
            .I(N__18068));
    InMux I__2337 (
            .O(N__18068),
            .I(N__18065));
    LocalMux I__2336 (
            .O(N__18065),
            .I(N__18062));
    Odrv4 I__2335 (
            .O(N__18062),
            .I(\b2v_inst11.mult1_un54_sum_cry_5_s ));
    InMux I__2334 (
            .O(N__18059),
            .I(\b2v_inst11.mult1_un54_sum_cry_4 ));
    InMux I__2333 (
            .O(N__18056),
            .I(N__18053));
    LocalMux I__2332 (
            .O(N__18053),
            .I(N__18050));
    Odrv4 I__2331 (
            .O(N__18050),
            .I(\b2v_inst11.mult1_un54_sum_cry_6_s ));
    InMux I__2330 (
            .O(N__18047),
            .I(\b2v_inst11.mult1_un54_sum_cry_5 ));
    InMux I__2329 (
            .O(N__18044),
            .I(N__18041));
    LocalMux I__2328 (
            .O(N__18041),
            .I(\b2v_inst11.un1_dutycycle_53_55_1_tz ));
    CascadeMux I__2327 (
            .O(N__18038),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_11_cascade_ ));
    InMux I__2326 (
            .O(N__18035),
            .I(N__18032));
    LocalMux I__2325 (
            .O(N__18032),
            .I(\b2v_inst11.un1_dutycycle_53_50_a0_1 ));
    CascadeMux I__2324 (
            .O(N__18029),
            .I(\b2v_inst11.un1_dutycycle_53_50_a0_1_cascade_ ));
    CascadeMux I__2323 (
            .O(N__18026),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_6_cascade_ ));
    CascadeMux I__2322 (
            .O(N__18023),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_12_cascade_ ));
    InMux I__2321 (
            .O(N__18020),
            .I(N__18017));
    LocalMux I__2320 (
            .O(N__18017),
            .I(\b2v_inst11.un1_dutycycle_53_4_1 ));
    InMux I__2319 (
            .O(N__18014),
            .I(N__18011));
    LocalMux I__2318 (
            .O(N__18011),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_12 ));
    CascadeMux I__2317 (
            .O(N__18008),
            .I(\b2v_inst11.un1_dutycycle_53_4_1_cascade_ ));
    InMux I__2316 (
            .O(N__18005),
            .I(N__17999));
    InMux I__2315 (
            .O(N__18004),
            .I(N__17999));
    LocalMux I__2314 (
            .O(N__17999),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_8 ));
    InMux I__2313 (
            .O(N__17996),
            .I(N__17993));
    LocalMux I__2312 (
            .O(N__17993),
            .I(N__17990));
    Span4Mux_h I__2311 (
            .O(N__17990),
            .I(N__17987));
    Odrv4 I__2310 (
            .O(N__17987),
            .I(\b2v_inst16.curr_state_2_1 ));
    InMux I__2309 (
            .O(N__17984),
            .I(N__17981));
    LocalMux I__2308 (
            .O(N__17981),
            .I(N__17978));
    Span4Mux_v I__2307 (
            .O(N__17978),
            .I(N__17975));
    Odrv4 I__2306 (
            .O(N__17975),
            .I(\b2v_inst16.curr_state_7_0_1 ));
    CascadeMux I__2305 (
            .O(N__17972),
            .I(\b2v_inst11.un1_dutycycle_53_44_0_2_cascade_ ));
    InMux I__2304 (
            .O(N__17969),
            .I(N__17966));
    LocalMux I__2303 (
            .O(N__17966),
            .I(\b2v_inst11.un2_count_clk_17_0_a2_1_4 ));
    CascadeMux I__2302 (
            .O(N__17963),
            .I(\b2v_inst11.N_355_cascade_ ));
    InMux I__2301 (
            .O(N__17960),
            .I(N__17954));
    InMux I__2300 (
            .O(N__17959),
            .I(N__17954));
    LocalMux I__2299 (
            .O(N__17954),
            .I(N__17951));
    Odrv4 I__2298 (
            .O(N__17951),
            .I(\b2v_inst16.count_rst_1 ));
    InMux I__2297 (
            .O(N__17948),
            .I(N__17945));
    LocalMux I__2296 (
            .O(N__17945),
            .I(\b2v_inst16.count_4_12 ));
    CascadeMux I__2295 (
            .O(N__17942),
            .I(N__17938));
    InMux I__2294 (
            .O(N__17941),
            .I(N__17935));
    InMux I__2293 (
            .O(N__17938),
            .I(N__17932));
    LocalMux I__2292 (
            .O(N__17935),
            .I(N__17929));
    LocalMux I__2291 (
            .O(N__17932),
            .I(\b2v_inst16.countZ0Z_13 ));
    Odrv4 I__2290 (
            .O(N__17929),
            .I(\b2v_inst16.countZ0Z_13 ));
    InMux I__2289 (
            .O(N__17924),
            .I(N__17918));
    InMux I__2288 (
            .O(N__17923),
            .I(N__17918));
    LocalMux I__2287 (
            .O(N__17918),
            .I(N__17915));
    Odrv4 I__2286 (
            .O(N__17915),
            .I(\b2v_inst16.count_rst_2 ));
    InMux I__2285 (
            .O(N__17912),
            .I(N__17909));
    LocalMux I__2284 (
            .O(N__17909),
            .I(\b2v_inst16.count_4_13 ));
    SRMux I__2283 (
            .O(N__17906),
            .I(N__17900));
    SRMux I__2282 (
            .O(N__17905),
            .I(N__17896));
    SRMux I__2281 (
            .O(N__17904),
            .I(N__17893));
    SRMux I__2280 (
            .O(N__17903),
            .I(N__17889));
    LocalMux I__2279 (
            .O(N__17900),
            .I(N__17885));
    SRMux I__2278 (
            .O(N__17899),
            .I(N__17882));
    LocalMux I__2277 (
            .O(N__17896),
            .I(N__17877));
    LocalMux I__2276 (
            .O(N__17893),
            .I(N__17877));
    SRMux I__2275 (
            .O(N__17892),
            .I(N__17874));
    LocalMux I__2274 (
            .O(N__17889),
            .I(N__17871));
    SRMux I__2273 (
            .O(N__17888),
            .I(N__17868));
    Span4Mux_v I__2272 (
            .O(N__17885),
            .I(N__17863));
    LocalMux I__2271 (
            .O(N__17882),
            .I(N__17863));
    Span4Mux_v I__2270 (
            .O(N__17877),
            .I(N__17860));
    LocalMux I__2269 (
            .O(N__17874),
            .I(N__17857));
    Span4Mux_v I__2268 (
            .O(N__17871),
            .I(N__17852));
    LocalMux I__2267 (
            .O(N__17868),
            .I(N__17852));
    Span4Mux_h I__2266 (
            .O(N__17863),
            .I(N__17849));
    Odrv4 I__2265 (
            .O(N__17860),
            .I(\b2v_inst16.N_3079_i ));
    Odrv4 I__2264 (
            .O(N__17857),
            .I(\b2v_inst16.N_3079_i ));
    Odrv4 I__2263 (
            .O(N__17852),
            .I(\b2v_inst16.N_3079_i ));
    Odrv4 I__2262 (
            .O(N__17849),
            .I(\b2v_inst16.N_3079_i ));
    InMux I__2261 (
            .O(N__17840),
            .I(N__17837));
    LocalMux I__2260 (
            .O(N__17837),
            .I(N__17834));
    Span4Mux_h I__2259 (
            .O(N__17834),
            .I(N__17831));
    Odrv4 I__2258 (
            .O(N__17831),
            .I(\b2v_inst16.count_4_3 ));
    InMux I__2257 (
            .O(N__17828),
            .I(N__17825));
    LocalMux I__2256 (
            .O(N__17825),
            .I(\b2v_inst16.count_rst_8 ));
    InMux I__2255 (
            .O(N__17822),
            .I(N__17818));
    InMux I__2254 (
            .O(N__17821),
            .I(N__17815));
    LocalMux I__2253 (
            .O(N__17818),
            .I(N__17811));
    LocalMux I__2252 (
            .O(N__17815),
            .I(N__17808));
    InMux I__2251 (
            .O(N__17814),
            .I(N__17804));
    Span4Mux_s3_h I__2250 (
            .O(N__17811),
            .I(N__17801));
    Span4Mux_s3_h I__2249 (
            .O(N__17808),
            .I(N__17798));
    InMux I__2248 (
            .O(N__17807),
            .I(N__17795));
    LocalMux I__2247 (
            .O(N__17804),
            .I(\b2v_inst16.countZ0Z_3 ));
    Odrv4 I__2246 (
            .O(N__17801),
            .I(\b2v_inst16.countZ0Z_3 ));
    Odrv4 I__2245 (
            .O(N__17798),
            .I(\b2v_inst16.countZ0Z_3 ));
    LocalMux I__2244 (
            .O(N__17795),
            .I(\b2v_inst16.countZ0Z_3 ));
    InMux I__2243 (
            .O(N__17786),
            .I(N__17780));
    InMux I__2242 (
            .O(N__17785),
            .I(N__17780));
    LocalMux I__2241 (
            .O(N__17780),
            .I(\b2v_inst11.dutycycleZ1Z_7 ));
    CascadeMux I__2240 (
            .O(N__17777),
            .I(\b2v_inst11.dutycycleZ1Z_3_cascade_ ));
    CascadeMux I__2239 (
            .O(N__17774),
            .I(\b2v_inst11.un1_dutycycle_53_axb_7_1_cascade_ ));
    IoInMux I__2238 (
            .O(N__17771),
            .I(N__17768));
    LocalMux I__2237 (
            .O(N__17768),
            .I(N__17765));
    Span4Mux_s3_h I__2236 (
            .O(N__17765),
            .I(N__17762));
    Span4Mux_h I__2235 (
            .O(N__17762),
            .I(N__17759));
    Span4Mux_v I__2234 (
            .O(N__17759),
            .I(N__17756));
    Span4Mux_v I__2233 (
            .O(N__17756),
            .I(N__17753));
    Odrv4 I__2232 (
            .O(N__17753),
            .I(vpp_en));
    InMux I__2231 (
            .O(N__17750),
            .I(N__17747));
    LocalMux I__2230 (
            .O(N__17747),
            .I(\b2v_inst16.delayed_vddq_pwrgd_eZ0Z_0 ));
    InMux I__2229 (
            .O(N__17744),
            .I(N__17738));
    CEMux I__2228 (
            .O(N__17743),
            .I(N__17738));
    LocalMux I__2227 (
            .O(N__17738),
            .I(N__17735));
    Odrv4 I__2226 (
            .O(N__17735),
            .I(\b2v_inst16.delayed_vddq_pwrgd_en ));
    CascadeMux I__2225 (
            .O(N__17732),
            .I(N__17718));
    CascadeMux I__2224 (
            .O(N__17731),
            .I(N__17705));
    CascadeMux I__2223 (
            .O(N__17730),
            .I(N__17701));
    InMux I__2222 (
            .O(N__17729),
            .I(N__17695));
    InMux I__2221 (
            .O(N__17728),
            .I(N__17692));
    InMux I__2220 (
            .O(N__17727),
            .I(N__17683));
    InMux I__2219 (
            .O(N__17726),
            .I(N__17683));
    InMux I__2218 (
            .O(N__17725),
            .I(N__17683));
    InMux I__2217 (
            .O(N__17724),
            .I(N__17683));
    InMux I__2216 (
            .O(N__17723),
            .I(N__17675));
    InMux I__2215 (
            .O(N__17722),
            .I(N__17675));
    InMux I__2214 (
            .O(N__17721),
            .I(N__17675));
    InMux I__2213 (
            .O(N__17718),
            .I(N__17662));
    InMux I__2212 (
            .O(N__17717),
            .I(N__17662));
    InMux I__2211 (
            .O(N__17716),
            .I(N__17662));
    InMux I__2210 (
            .O(N__17715),
            .I(N__17662));
    InMux I__2209 (
            .O(N__17714),
            .I(N__17662));
    InMux I__2208 (
            .O(N__17713),
            .I(N__17662));
    InMux I__2207 (
            .O(N__17712),
            .I(N__17653));
    InMux I__2206 (
            .O(N__17711),
            .I(N__17653));
    InMux I__2205 (
            .O(N__17710),
            .I(N__17653));
    InMux I__2204 (
            .O(N__17709),
            .I(N__17653));
    InMux I__2203 (
            .O(N__17708),
            .I(N__17642));
    InMux I__2202 (
            .O(N__17705),
            .I(N__17642));
    InMux I__2201 (
            .O(N__17704),
            .I(N__17642));
    InMux I__2200 (
            .O(N__17701),
            .I(N__17642));
    InMux I__2199 (
            .O(N__17700),
            .I(N__17642));
    InMux I__2198 (
            .O(N__17699),
            .I(N__17639));
    InMux I__2197 (
            .O(N__17698),
            .I(N__17636));
    LocalMux I__2196 (
            .O(N__17695),
            .I(N__17633));
    LocalMux I__2195 (
            .O(N__17692),
            .I(N__17628));
    LocalMux I__2194 (
            .O(N__17683),
            .I(N__17628));
    InMux I__2193 (
            .O(N__17682),
            .I(N__17625));
    LocalMux I__2192 (
            .O(N__17675),
            .I(N__17620));
    LocalMux I__2191 (
            .O(N__17662),
            .I(N__17620));
    LocalMux I__2190 (
            .O(N__17653),
            .I(N__17615));
    LocalMux I__2189 (
            .O(N__17642),
            .I(N__17615));
    LocalMux I__2188 (
            .O(N__17639),
            .I(N__17611));
    LocalMux I__2187 (
            .O(N__17636),
            .I(N__17608));
    Span4Mux_s2_v I__2186 (
            .O(N__17633),
            .I(N__17601));
    Span4Mux_v I__2185 (
            .O(N__17628),
            .I(N__17601));
    LocalMux I__2184 (
            .O(N__17625),
            .I(N__17601));
    Span4Mux_s3_h I__2183 (
            .O(N__17620),
            .I(N__17598));
    Span4Mux_s3_h I__2182 (
            .O(N__17615),
            .I(N__17595));
    InMux I__2181 (
            .O(N__17614),
            .I(N__17592));
    Odrv12 I__2180 (
            .O(N__17611),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__2179 (
            .O(N__17608),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__2178 (
            .O(N__17601),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__2177 (
            .O(N__17598),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__2176 (
            .O(N__17595),
            .I(\b2v_inst16.N_26 ));
    LocalMux I__2175 (
            .O(N__17592),
            .I(\b2v_inst16.N_26 ));
    CascadeMux I__2174 (
            .O(N__17579),
            .I(N__17572));
    InMux I__2173 (
            .O(N__17578),
            .I(N__17561));
    InMux I__2172 (
            .O(N__17577),
            .I(N__17550));
    InMux I__2171 (
            .O(N__17576),
            .I(N__17550));
    InMux I__2170 (
            .O(N__17575),
            .I(N__17550));
    InMux I__2169 (
            .O(N__17572),
            .I(N__17550));
    InMux I__2168 (
            .O(N__17571),
            .I(N__17550));
    InMux I__2167 (
            .O(N__17570),
            .I(N__17547));
    InMux I__2166 (
            .O(N__17569),
            .I(N__17544));
    InMux I__2165 (
            .O(N__17568),
            .I(N__17532));
    InMux I__2164 (
            .O(N__17567),
            .I(N__17532));
    InMux I__2163 (
            .O(N__17566),
            .I(N__17532));
    InMux I__2162 (
            .O(N__17565),
            .I(N__17532));
    InMux I__2161 (
            .O(N__17564),
            .I(N__17529));
    LocalMux I__2160 (
            .O(N__17561),
            .I(N__17524));
    LocalMux I__2159 (
            .O(N__17550),
            .I(N__17524));
    LocalMux I__2158 (
            .O(N__17547),
            .I(N__17519));
    LocalMux I__2157 (
            .O(N__17544),
            .I(N__17519));
    InMux I__2156 (
            .O(N__17543),
            .I(N__17516));
    InMux I__2155 (
            .O(N__17542),
            .I(N__17511));
    InMux I__2154 (
            .O(N__17541),
            .I(N__17511));
    LocalMux I__2153 (
            .O(N__17532),
            .I(N__17508));
    LocalMux I__2152 (
            .O(N__17529),
            .I(N__17503));
    Span4Mux_s0_v I__2151 (
            .O(N__17524),
            .I(N__17503));
    Span12Mux_s2_v I__2150 (
            .O(N__17519),
            .I(N__17500));
    LocalMux I__2149 (
            .O(N__17516),
            .I(\b2v_inst16.N_416 ));
    LocalMux I__2148 (
            .O(N__17511),
            .I(\b2v_inst16.N_416 ));
    Odrv4 I__2147 (
            .O(N__17508),
            .I(\b2v_inst16.N_416 ));
    Odrv4 I__2146 (
            .O(N__17503),
            .I(\b2v_inst16.N_416 ));
    Odrv12 I__2145 (
            .O(N__17500),
            .I(\b2v_inst16.N_416 ));
    CascadeMux I__2144 (
            .O(N__17489),
            .I(N__17485));
    InMux I__2143 (
            .O(N__17488),
            .I(N__17482));
    InMux I__2142 (
            .O(N__17485),
            .I(N__17479));
    LocalMux I__2141 (
            .O(N__17482),
            .I(N__17476));
    LocalMux I__2140 (
            .O(N__17479),
            .I(N__17473));
    Odrv4 I__2139 (
            .O(N__17476),
            .I(\b2v_inst16.un4_count_1_cry_2_THRU_CO ));
    Odrv4 I__2138 (
            .O(N__17473),
            .I(\b2v_inst16.un4_count_1_cry_2_THRU_CO ));
    CascadeMux I__2137 (
            .O(N__17468),
            .I(\b2v_inst16.N_26_cascade_ ));
    InMux I__2136 (
            .O(N__17465),
            .I(N__17462));
    LocalMux I__2135 (
            .O(N__17462),
            .I(N__17459));
    Span4Mux_s3_h I__2134 (
            .O(N__17459),
            .I(N__17456));
    Odrv4 I__2133 (
            .O(N__17456),
            .I(\b2v_inst16.count_4_i_a3_10_0 ));
    InMux I__2132 (
            .O(N__17453),
            .I(N__17449));
    InMux I__2131 (
            .O(N__17452),
            .I(N__17446));
    LocalMux I__2130 (
            .O(N__17449),
            .I(N__17443));
    LocalMux I__2129 (
            .O(N__17446),
            .I(\b2v_inst16.countZ0Z_14 ));
    Odrv4 I__2128 (
            .O(N__17443),
            .I(\b2v_inst16.countZ0Z_14 ));
    InMux I__2127 (
            .O(N__17438),
            .I(N__17432));
    InMux I__2126 (
            .O(N__17437),
            .I(N__17432));
    LocalMux I__2125 (
            .O(N__17432),
            .I(N__17429));
    Odrv12 I__2124 (
            .O(N__17429),
            .I(\b2v_inst16.count_rst_3 ));
    InMux I__2123 (
            .O(N__17426),
            .I(N__17423));
    LocalMux I__2122 (
            .O(N__17423),
            .I(\b2v_inst16.count_4_14 ));
    InMux I__2121 (
            .O(N__17420),
            .I(N__17416));
    InMux I__2120 (
            .O(N__17419),
            .I(N__17413));
    LocalMux I__2119 (
            .O(N__17416),
            .I(N__17410));
    LocalMux I__2118 (
            .O(N__17413),
            .I(\b2v_inst16.countZ0Z_12 ));
    Odrv4 I__2117 (
            .O(N__17410),
            .I(\b2v_inst16.countZ0Z_12 ));
    CascadeMux I__2116 (
            .O(N__17405),
            .I(N__17402));
    InMux I__2115 (
            .O(N__17402),
            .I(N__17396));
    InMux I__2114 (
            .O(N__17401),
            .I(N__17396));
    LocalMux I__2113 (
            .O(N__17396),
            .I(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ));
    InMux I__2112 (
            .O(N__17393),
            .I(N__17390));
    LocalMux I__2111 (
            .O(N__17390),
            .I(\b2v_inst11.count_0_15 ));
    CascadeMux I__2110 (
            .O(N__17387),
            .I(N__17384));
    InMux I__2109 (
            .O(N__17384),
            .I(N__17378));
    InMux I__2108 (
            .O(N__17383),
            .I(N__17378));
    LocalMux I__2107 (
            .O(N__17378),
            .I(\b2v_inst11.count_1_7 ));
    InMux I__2106 (
            .O(N__17375),
            .I(N__17372));
    LocalMux I__2105 (
            .O(N__17372),
            .I(\b2v_inst11.count_0_7 ));
    IoInMux I__2104 (
            .O(N__17369),
            .I(N__17366));
    LocalMux I__2103 (
            .O(N__17366),
            .I(N__17363));
    Span4Mux_s3_h I__2102 (
            .O(N__17363),
            .I(N__17360));
    Sp12to4 I__2101 (
            .O(N__17360),
            .I(N__17357));
    Odrv12 I__2100 (
            .O(N__17357),
            .I(\b2v_inst200.count_enZ0 ));
    IoInMux I__2099 (
            .O(N__17354),
            .I(N__17351));
    LocalMux I__2098 (
            .O(N__17351),
            .I(N__17348));
    IoSpan4Mux I__2097 (
            .O(N__17348),
            .I(N__17345));
    Span4Mux_s0_h I__2096 (
            .O(N__17345),
            .I(N__17341));
    IoInMux I__2095 (
            .O(N__17344),
            .I(N__17338));
    Sp12to4 I__2094 (
            .O(N__17341),
            .I(N__17334));
    LocalMux I__2093 (
            .O(N__17338),
            .I(N__17331));
    IoInMux I__2092 (
            .O(N__17337),
            .I(N__17328));
    Span12Mux_s8_h I__2091 (
            .O(N__17334),
            .I(N__17325));
    IoSpan4Mux I__2090 (
            .O(N__17331),
            .I(N__17322));
    LocalMux I__2089 (
            .O(N__17328),
            .I(N__17319));
    Odrv12 I__2088 (
            .O(N__17325),
            .I(pch_pwrok));
    Odrv4 I__2087 (
            .O(N__17322),
            .I(pch_pwrok));
    Odrv12 I__2086 (
            .O(N__17319),
            .I(pch_pwrok));
    CascadeMux I__2085 (
            .O(N__17312),
            .I(\b2v_inst11.un79_clk_100khzlt6_cascade_ ));
    CascadeMux I__2084 (
            .O(N__17309),
            .I(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ));
    CascadeMux I__2083 (
            .O(N__17306),
            .I(\b2v_inst11.un79_clk_100khzlto15_7_cascade_ ));
    InMux I__2082 (
            .O(N__17303),
            .I(N__17300));
    LocalMux I__2081 (
            .O(N__17300),
            .I(\b2v_inst11.un79_clk_100khzlto15_3 ));
    CascadeMux I__2080 (
            .O(N__17297),
            .I(\b2v_inst11.count_RNIZ0Z_8_cascade_ ));
    InMux I__2079 (
            .O(N__17294),
            .I(N__17288));
    InMux I__2078 (
            .O(N__17293),
            .I(N__17288));
    LocalMux I__2077 (
            .O(N__17288),
            .I(N__17285));
    Odrv4 I__2076 (
            .O(N__17285),
            .I(\b2v_inst11.N_8 ));
    InMux I__2075 (
            .O(N__17282),
            .I(N__17276));
    InMux I__2074 (
            .O(N__17281),
            .I(N__17276));
    LocalMux I__2073 (
            .O(N__17276),
            .I(\b2v_inst11.count_1_14 ));
    InMux I__2072 (
            .O(N__17273),
            .I(N__17270));
    LocalMux I__2071 (
            .O(N__17270),
            .I(\b2v_inst11.count_0_14 ));
    CascadeMux I__2070 (
            .O(N__17267),
            .I(N__17264));
    InMux I__2069 (
            .O(N__17264),
            .I(N__17258));
    InMux I__2068 (
            .O(N__17263),
            .I(N__17258));
    LocalMux I__2067 (
            .O(N__17258),
            .I(\b2v_inst11.count_1_6 ));
    InMux I__2066 (
            .O(N__17255),
            .I(N__17252));
    LocalMux I__2065 (
            .O(N__17252),
            .I(\b2v_inst11.count_0_6 ));
    CascadeMux I__2064 (
            .O(N__17249),
            .I(N__17246));
    InMux I__2063 (
            .O(N__17246),
            .I(N__17240));
    InMux I__2062 (
            .O(N__17245),
            .I(N__17240));
    LocalMux I__2061 (
            .O(N__17240),
            .I(\b2v_inst11.count_1_3 ));
    InMux I__2060 (
            .O(N__17237),
            .I(N__17234));
    LocalMux I__2059 (
            .O(N__17234),
            .I(\b2v_inst11.count_0_3 ));
    InMux I__2058 (
            .O(N__17231),
            .I(N__17225));
    InMux I__2057 (
            .O(N__17230),
            .I(N__17225));
    LocalMux I__2056 (
            .O(N__17225),
            .I(N__17222));
    Odrv4 I__2055 (
            .O(N__17222),
            .I(\b2v_inst11.count_1_13 ));
    InMux I__2054 (
            .O(N__17219),
            .I(N__17216));
    LocalMux I__2053 (
            .O(N__17216),
            .I(\b2v_inst11.count_0_13 ));
    CascadeMux I__2052 (
            .O(N__17213),
            .I(N__17210));
    InMux I__2051 (
            .O(N__17210),
            .I(N__17204));
    InMux I__2050 (
            .O(N__17209),
            .I(N__17204));
    LocalMux I__2049 (
            .O(N__17204),
            .I(\b2v_inst11.count_1_4 ));
    InMux I__2048 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__2047 (
            .O(N__17198),
            .I(\b2v_inst11.count_0_4 ));
    CascadeMux I__2046 (
            .O(N__17195),
            .I(N__17192));
    InMux I__2045 (
            .O(N__17192),
            .I(N__17186));
    InMux I__2044 (
            .O(N__17191),
            .I(N__17186));
    LocalMux I__2043 (
            .O(N__17186),
            .I(\b2v_inst11.count_1_5 ));
    InMux I__2042 (
            .O(N__17183),
            .I(N__17180));
    LocalMux I__2041 (
            .O(N__17180),
            .I(\b2v_inst11.count_0_5 ));
    SRMux I__2040 (
            .O(N__17177),
            .I(N__17174));
    LocalMux I__2039 (
            .O(N__17174),
            .I(N__17171));
    Odrv12 I__2038 (
            .O(N__17171),
            .I(\b2v_inst11.pwm_out_1_sqmuxa ));
    IoInMux I__2037 (
            .O(N__17168),
            .I(N__17165));
    LocalMux I__2036 (
            .O(N__17165),
            .I(N__17162));
    Odrv12 I__2035 (
            .O(N__17162),
            .I(pwrbtn_led));
    CascadeMux I__2034 (
            .O(N__17159),
            .I(\b2v_inst11.curr_state_3_0_cascade_ ));
    CascadeMux I__2033 (
            .O(N__17156),
            .I(\b2v_inst11.curr_stateZ0Z_0_cascade_ ));
    InMux I__2032 (
            .O(N__17153),
            .I(N__17132));
    InMux I__2031 (
            .O(N__17152),
            .I(N__17132));
    InMux I__2030 (
            .O(N__17151),
            .I(N__17132));
    InMux I__2029 (
            .O(N__17150),
            .I(N__17123));
    InMux I__2028 (
            .O(N__17149),
            .I(N__17123));
    InMux I__2027 (
            .O(N__17148),
            .I(N__17123));
    InMux I__2026 (
            .O(N__17147),
            .I(N__17123));
    InMux I__2025 (
            .O(N__17146),
            .I(N__17114));
    InMux I__2024 (
            .O(N__17145),
            .I(N__17114));
    InMux I__2023 (
            .O(N__17144),
            .I(N__17114));
    InMux I__2022 (
            .O(N__17143),
            .I(N__17114));
    CascadeMux I__2021 (
            .O(N__17142),
            .I(N__17110));
    InMux I__2020 (
            .O(N__17141),
            .I(N__17102));
    InMux I__2019 (
            .O(N__17140),
            .I(N__17102));
    InMux I__2018 (
            .O(N__17139),
            .I(N__17102));
    LocalMux I__2017 (
            .O(N__17132),
            .I(N__17095));
    LocalMux I__2016 (
            .O(N__17123),
            .I(N__17095));
    LocalMux I__2015 (
            .O(N__17114),
            .I(N__17095));
    InMux I__2014 (
            .O(N__17113),
            .I(N__17088));
    InMux I__2013 (
            .O(N__17110),
            .I(N__17088));
    InMux I__2012 (
            .O(N__17109),
            .I(N__17088));
    LocalMux I__2011 (
            .O(N__17102),
            .I(N__17085));
    Span4Mux_s2_v I__2010 (
            .O(N__17095),
            .I(N__17082));
    LocalMux I__2009 (
            .O(N__17088),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    Odrv4 I__2008 (
            .O(N__17085),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    Odrv4 I__2007 (
            .O(N__17082),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    CascadeMux I__2006 (
            .O(N__17075),
            .I(\b2v_inst11.count_0_sqmuxa_i_cascade_ ));
    CascadeMux I__2005 (
            .O(N__17072),
            .I(\b2v_inst11.count_1_0_cascade_ ));
    InMux I__2004 (
            .O(N__17069),
            .I(N__17066));
    LocalMux I__2003 (
            .O(N__17066),
            .I(\b2v_inst11.count_0_0 ));
    InMux I__2002 (
            .O(N__17063),
            .I(N__17057));
    InMux I__2001 (
            .O(N__17062),
            .I(N__17057));
    LocalMux I__2000 (
            .O(N__17057),
            .I(\b2v_inst11.pwm_outZ0 ));
    CascadeMux I__1999 (
            .O(N__17054),
            .I(N__17050));
    CascadeMux I__1998 (
            .O(N__17053),
            .I(N__17047));
    InMux I__1997 (
            .O(N__17050),
            .I(N__17042));
    InMux I__1996 (
            .O(N__17047),
            .I(N__17042));
    LocalMux I__1995 (
            .O(N__17042),
            .I(\b2v_inst11.g0_i_o3_0 ));
    InMux I__1994 (
            .O(N__17039),
            .I(\b2v_inst11.mult1_un103_sum_cry_2 ));
    CascadeMux I__1993 (
            .O(N__17036),
            .I(N__17033));
    InMux I__1992 (
            .O(N__17033),
            .I(N__17030));
    LocalMux I__1991 (
            .O(N__17030),
            .I(\b2v_inst11.mult1_un96_sum_cry_3_s ));
    InMux I__1990 (
            .O(N__17027),
            .I(\b2v_inst11.mult1_un103_sum_cry_3 ));
    InMux I__1989 (
            .O(N__17024),
            .I(N__17021));
    LocalMux I__1988 (
            .O(N__17021),
            .I(\b2v_inst11.mult1_un96_sum_cry_4_s ));
    InMux I__1987 (
            .O(N__17018),
            .I(\b2v_inst11.mult1_un103_sum_cry_4 ));
    CascadeMux I__1986 (
            .O(N__17015),
            .I(N__17010));
    InMux I__1985 (
            .O(N__17014),
            .I(N__17006));
    InMux I__1984 (
            .O(N__17013),
            .I(N__17001));
    InMux I__1983 (
            .O(N__17010),
            .I(N__17001));
    InMux I__1982 (
            .O(N__17009),
            .I(N__16998));
    LocalMux I__1981 (
            .O(N__17006),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    LocalMux I__1980 (
            .O(N__17001),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    LocalMux I__1979 (
            .O(N__16998),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    CascadeMux I__1978 (
            .O(N__16991),
            .I(N__16988));
    InMux I__1977 (
            .O(N__16988),
            .I(N__16985));
    LocalMux I__1976 (
            .O(N__16985),
            .I(\b2v_inst11.mult1_un96_sum_cry_5_s ));
    InMux I__1975 (
            .O(N__16982),
            .I(\b2v_inst11.mult1_un103_sum_cry_5 ));
    InMux I__1974 (
            .O(N__16979),
            .I(N__16976));
    LocalMux I__1973 (
            .O(N__16976),
            .I(\b2v_inst11.mult1_un96_sum_cry_6_s ));
    CascadeMux I__1972 (
            .O(N__16973),
            .I(N__16969));
    CascadeMux I__1971 (
            .O(N__16972),
            .I(N__16965));
    InMux I__1970 (
            .O(N__16969),
            .I(N__16958));
    InMux I__1969 (
            .O(N__16968),
            .I(N__16958));
    InMux I__1968 (
            .O(N__16965),
            .I(N__16958));
    LocalMux I__1967 (
            .O(N__16958),
            .I(\b2v_inst11.mult1_un96_sum_i_0_8 ));
    InMux I__1966 (
            .O(N__16955),
            .I(\b2v_inst11.mult1_un103_sum_cry_6 ));
    CascadeMux I__1965 (
            .O(N__16952),
            .I(N__16949));
    InMux I__1964 (
            .O(N__16949),
            .I(N__16946));
    LocalMux I__1963 (
            .O(N__16946),
            .I(\b2v_inst11.mult1_un103_sum_axb_8 ));
    InMux I__1962 (
            .O(N__16943),
            .I(\b2v_inst11.mult1_un103_sum_cry_7 ));
    CascadeMux I__1961 (
            .O(N__16940),
            .I(N__16935));
    InMux I__1960 (
            .O(N__16939),
            .I(N__16931));
    InMux I__1959 (
            .O(N__16938),
            .I(N__16926));
    InMux I__1958 (
            .O(N__16935),
            .I(N__16926));
    InMux I__1957 (
            .O(N__16934),
            .I(N__16923));
    LocalMux I__1956 (
            .O(N__16931),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__1955 (
            .O(N__16926),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__1954 (
            .O(N__16923),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    InMux I__1953 (
            .O(N__16916),
            .I(N__16913));
    LocalMux I__1952 (
            .O(N__16913),
            .I(\b2v_inst11.mult1_un75_sum_cry_6_s ));
    CascadeMux I__1951 (
            .O(N__16910),
            .I(N__16906));
    CascadeMux I__1950 (
            .O(N__16909),
            .I(N__16902));
    InMux I__1949 (
            .O(N__16906),
            .I(N__16895));
    InMux I__1948 (
            .O(N__16905),
            .I(N__16895));
    InMux I__1947 (
            .O(N__16902),
            .I(N__16895));
    LocalMux I__1946 (
            .O(N__16895),
            .I(\b2v_inst11.mult1_un75_sum_i_0_8 ));
    CascadeMux I__1945 (
            .O(N__16892),
            .I(N__16889));
    InMux I__1944 (
            .O(N__16889),
            .I(N__16886));
    LocalMux I__1943 (
            .O(N__16886),
            .I(\b2v_inst11.mult1_un89_sum_axb_8 ));
    InMux I__1942 (
            .O(N__16883),
            .I(\b2v_inst11.mult1_un82_sum_cry_6 ));
    CascadeMux I__1941 (
            .O(N__16880),
            .I(N__16877));
    InMux I__1940 (
            .O(N__16877),
            .I(N__16874));
    LocalMux I__1939 (
            .O(N__16874),
            .I(\b2v_inst11.mult1_un82_sum_axb_8 ));
    InMux I__1938 (
            .O(N__16871),
            .I(\b2v_inst11.mult1_un82_sum_cry_7 ));
    CascadeMux I__1937 (
            .O(N__16868),
            .I(N__16864));
    CascadeMux I__1936 (
            .O(N__16867),
            .I(N__16860));
    InMux I__1935 (
            .O(N__16864),
            .I(N__16853));
    InMux I__1934 (
            .O(N__16863),
            .I(N__16853));
    InMux I__1933 (
            .O(N__16860),
            .I(N__16853));
    LocalMux I__1932 (
            .O(N__16853),
            .I(\b2v_inst11.mult1_un54_sum_i_8 ));
    CascadeMux I__1931 (
            .O(N__16850),
            .I(N__16845));
    InMux I__1930 (
            .O(N__16849),
            .I(N__16841));
    InMux I__1929 (
            .O(N__16848),
            .I(N__16836));
    InMux I__1928 (
            .O(N__16845),
            .I(N__16836));
    InMux I__1927 (
            .O(N__16844),
            .I(N__16833));
    LocalMux I__1926 (
            .O(N__16841),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__1925 (
            .O(N__16836),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__1924 (
            .O(N__16833),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    InMux I__1923 (
            .O(N__16826),
            .I(N__16823));
    LocalMux I__1922 (
            .O(N__16823),
            .I(\b2v_inst11.mult1_un68_sum_i ));
    InMux I__1921 (
            .O(N__16820),
            .I(N__16817));
    LocalMux I__1920 (
            .O(N__16817),
            .I(\b2v_inst11.mult1_un82_sum_i ));
    InMux I__1919 (
            .O(N__16814),
            .I(N__16811));
    LocalMux I__1918 (
            .O(N__16811),
            .I(N__16808));
    Span4Mux_s1_h I__1917 (
            .O(N__16808),
            .I(N__16805));
    Odrv4 I__1916 (
            .O(N__16805),
            .I(\b2v_inst11.mult1_un89_sum_i ));
    CascadeMux I__1915 (
            .O(N__16802),
            .I(N__16798));
    CascadeMux I__1914 (
            .O(N__16801),
            .I(N__16794));
    InMux I__1913 (
            .O(N__16798),
            .I(N__16787));
    InMux I__1912 (
            .O(N__16797),
            .I(N__16787));
    InMux I__1911 (
            .O(N__16794),
            .I(N__16787));
    LocalMux I__1910 (
            .O(N__16787),
            .I(\b2v_inst11.mult1_un82_sum_i_0_8 ));
    CascadeMux I__1909 (
            .O(N__16784),
            .I(N__16780));
    InMux I__1908 (
            .O(N__16783),
            .I(N__16772));
    InMux I__1907 (
            .O(N__16780),
            .I(N__16772));
    InMux I__1906 (
            .O(N__16779),
            .I(N__16769));
    InMux I__1905 (
            .O(N__16778),
            .I(N__16764));
    InMux I__1904 (
            .O(N__16777),
            .I(N__16764));
    LocalMux I__1903 (
            .O(N__16772),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__1902 (
            .O(N__16769),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__1901 (
            .O(N__16764),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    CascadeMux I__1900 (
            .O(N__16757),
            .I(N__16754));
    InMux I__1899 (
            .O(N__16754),
            .I(N__16751));
    LocalMux I__1898 (
            .O(N__16751),
            .I(\b2v_inst11.mult1_un68_sum_axb_8 ));
    InMux I__1897 (
            .O(N__16748),
            .I(\b2v_inst11.mult1_un61_sum_cry_6 ));
    InMux I__1896 (
            .O(N__16745),
            .I(\b2v_inst11.mult1_un61_sum_cry_7 ));
    CascadeMux I__1895 (
            .O(N__16742),
            .I(\b2v_inst11.mult1_un61_sum_s_8_cascade_ ));
    CascadeMux I__1894 (
            .O(N__16739),
            .I(N__16735));
    CascadeMux I__1893 (
            .O(N__16738),
            .I(N__16731));
    InMux I__1892 (
            .O(N__16735),
            .I(N__16724));
    InMux I__1891 (
            .O(N__16734),
            .I(N__16724));
    InMux I__1890 (
            .O(N__16731),
            .I(N__16724));
    LocalMux I__1889 (
            .O(N__16724),
            .I(\b2v_inst11.mult1_un61_sum_i_0_8 ));
    CascadeMux I__1888 (
            .O(N__16721),
            .I(N__16718));
    InMux I__1887 (
            .O(N__16718),
            .I(N__16715));
    LocalMux I__1886 (
            .O(N__16715),
            .I(\b2v_inst11.mult1_un82_sum_cry_3_s ));
    InMux I__1885 (
            .O(N__16712),
            .I(\b2v_inst11.mult1_un82_sum_cry_2 ));
    CascadeMux I__1884 (
            .O(N__16709),
            .I(N__16706));
    InMux I__1883 (
            .O(N__16706),
            .I(N__16703));
    LocalMux I__1882 (
            .O(N__16703),
            .I(\b2v_inst11.mult1_un75_sum_cry_3_s ));
    InMux I__1881 (
            .O(N__16700),
            .I(N__16697));
    LocalMux I__1880 (
            .O(N__16697),
            .I(\b2v_inst11.mult1_un82_sum_cry_4_s ));
    InMux I__1879 (
            .O(N__16694),
            .I(\b2v_inst11.mult1_un82_sum_cry_3 ));
    InMux I__1878 (
            .O(N__16691),
            .I(N__16688));
    LocalMux I__1877 (
            .O(N__16688),
            .I(\b2v_inst11.mult1_un75_sum_cry_4_s ));
    CascadeMux I__1876 (
            .O(N__16685),
            .I(N__16682));
    InMux I__1875 (
            .O(N__16682),
            .I(N__16679));
    LocalMux I__1874 (
            .O(N__16679),
            .I(\b2v_inst11.mult1_un82_sum_cry_5_s ));
    InMux I__1873 (
            .O(N__16676),
            .I(\b2v_inst11.mult1_un82_sum_cry_4 ));
    CascadeMux I__1872 (
            .O(N__16673),
            .I(N__16670));
    InMux I__1871 (
            .O(N__16670),
            .I(N__16667));
    LocalMux I__1870 (
            .O(N__16667),
            .I(\b2v_inst11.mult1_un75_sum_cry_5_s ));
    InMux I__1869 (
            .O(N__16664),
            .I(N__16661));
    LocalMux I__1868 (
            .O(N__16661),
            .I(\b2v_inst11.mult1_un82_sum_cry_6_s ));
    InMux I__1867 (
            .O(N__16658),
            .I(\b2v_inst11.mult1_un82_sum_cry_5 ));
    InMux I__1866 (
            .O(N__16655),
            .I(N__16649));
    InMux I__1865 (
            .O(N__16654),
            .I(N__16649));
    LocalMux I__1864 (
            .O(N__16649),
            .I(\b2v_inst200.count_3_13 ));
    InMux I__1863 (
            .O(N__16646),
            .I(N__16637));
    InMux I__1862 (
            .O(N__16645),
            .I(N__16637));
    InMux I__1861 (
            .O(N__16644),
            .I(N__16637));
    LocalMux I__1860 (
            .O(N__16637),
            .I(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ));
    InMux I__1859 (
            .O(N__16634),
            .I(N__16631));
    LocalMux I__1858 (
            .O(N__16631),
            .I(\b2v_inst200.un2_count_1_axb_13 ));
    InMux I__1857 (
            .O(N__16628),
            .I(N__16625));
    LocalMux I__1856 (
            .O(N__16625),
            .I(N__16622));
    Span4Mux_v I__1855 (
            .O(N__16622),
            .I(N__16617));
    InMux I__1854 (
            .O(N__16621),
            .I(N__16612));
    InMux I__1853 (
            .O(N__16620),
            .I(N__16612));
    Odrv4 I__1852 (
            .O(N__16617),
            .I(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ));
    LocalMux I__1851 (
            .O(N__16612),
            .I(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ));
    InMux I__1850 (
            .O(N__16607),
            .I(N__16603));
    InMux I__1849 (
            .O(N__16606),
            .I(N__16600));
    LocalMux I__1848 (
            .O(N__16603),
            .I(\b2v_inst200.count_3_5 ));
    LocalMux I__1847 (
            .O(N__16600),
            .I(\b2v_inst200.count_3_5 ));
    CascadeMux I__1846 (
            .O(N__16595),
            .I(N__16592));
    InMux I__1845 (
            .O(N__16592),
            .I(N__16588));
    CascadeMux I__1844 (
            .O(N__16591),
            .I(N__16585));
    LocalMux I__1843 (
            .O(N__16588),
            .I(N__16582));
    InMux I__1842 (
            .O(N__16585),
            .I(N__16579));
    Odrv12 I__1841 (
            .O(N__16582),
            .I(\b2v_inst200.countZ0Z_7 ));
    LocalMux I__1840 (
            .O(N__16579),
            .I(\b2v_inst200.countZ0Z_7 ));
    InMux I__1839 (
            .O(N__16574),
            .I(N__16540));
    InMux I__1838 (
            .O(N__16573),
            .I(N__16540));
    InMux I__1837 (
            .O(N__16572),
            .I(N__16540));
    InMux I__1836 (
            .O(N__16571),
            .I(N__16540));
    InMux I__1835 (
            .O(N__16570),
            .I(N__16529));
    InMux I__1834 (
            .O(N__16569),
            .I(N__16529));
    InMux I__1833 (
            .O(N__16568),
            .I(N__16529));
    InMux I__1832 (
            .O(N__16567),
            .I(N__16529));
    InMux I__1831 (
            .O(N__16566),
            .I(N__16529));
    InMux I__1830 (
            .O(N__16565),
            .I(N__16524));
    InMux I__1829 (
            .O(N__16564),
            .I(N__16524));
    InMux I__1828 (
            .O(N__16563),
            .I(N__16515));
    InMux I__1827 (
            .O(N__16562),
            .I(N__16515));
    InMux I__1826 (
            .O(N__16561),
            .I(N__16515));
    InMux I__1825 (
            .O(N__16560),
            .I(N__16515));
    InMux I__1824 (
            .O(N__16559),
            .I(N__16502));
    InMux I__1823 (
            .O(N__16558),
            .I(N__16502));
    InMux I__1822 (
            .O(N__16557),
            .I(N__16502));
    InMux I__1821 (
            .O(N__16556),
            .I(N__16502));
    InMux I__1820 (
            .O(N__16555),
            .I(N__16502));
    InMux I__1819 (
            .O(N__16554),
            .I(N__16502));
    InMux I__1818 (
            .O(N__16553),
            .I(N__16491));
    InMux I__1817 (
            .O(N__16552),
            .I(N__16491));
    InMux I__1816 (
            .O(N__16551),
            .I(N__16491));
    InMux I__1815 (
            .O(N__16550),
            .I(N__16491));
    InMux I__1814 (
            .O(N__16549),
            .I(N__16491));
    LocalMux I__1813 (
            .O(N__16540),
            .I(N__16482));
    LocalMux I__1812 (
            .O(N__16529),
            .I(N__16479));
    LocalMux I__1811 (
            .O(N__16524),
            .I(N__16476));
    LocalMux I__1810 (
            .O(N__16515),
            .I(N__16473));
    LocalMux I__1809 (
            .O(N__16502),
            .I(N__16470));
    LocalMux I__1808 (
            .O(N__16491),
            .I(N__16467));
    CEMux I__1807 (
            .O(N__16490),
            .I(N__16442));
    CEMux I__1806 (
            .O(N__16489),
            .I(N__16442));
    CEMux I__1805 (
            .O(N__16488),
            .I(N__16442));
    CEMux I__1804 (
            .O(N__16487),
            .I(N__16442));
    CEMux I__1803 (
            .O(N__16486),
            .I(N__16442));
    CEMux I__1802 (
            .O(N__16485),
            .I(N__16442));
    Glb2LocalMux I__1801 (
            .O(N__16482),
            .I(N__16442));
    Glb2LocalMux I__1800 (
            .O(N__16479),
            .I(N__16442));
    Glb2LocalMux I__1799 (
            .O(N__16476),
            .I(N__16442));
    Glb2LocalMux I__1798 (
            .O(N__16473),
            .I(N__16442));
    Glb2LocalMux I__1797 (
            .O(N__16470),
            .I(N__16442));
    Glb2LocalMux I__1796 (
            .O(N__16467),
            .I(N__16442));
    GlobalMux I__1795 (
            .O(N__16442),
            .I(N__16439));
    gio2CtrlBuf I__1794 (
            .O(N__16439),
            .I(\b2v_inst200.count_en_g ));
    InMux I__1793 (
            .O(N__16436),
            .I(N__16433));
    LocalMux I__1792 (
            .O(N__16433),
            .I(\b2v_inst200.un25_clk_100khz_3 ));
    CascadeMux I__1791 (
            .O(N__16430),
            .I(N__16427));
    InMux I__1790 (
            .O(N__16427),
            .I(N__16424));
    LocalMux I__1789 (
            .O(N__16424),
            .I(\b2v_inst11.mult1_un61_sum_cry_3_s ));
    InMux I__1788 (
            .O(N__16421),
            .I(\b2v_inst11.mult1_un61_sum_cry_2 ));
    InMux I__1787 (
            .O(N__16418),
            .I(N__16415));
    LocalMux I__1786 (
            .O(N__16415),
            .I(\b2v_inst11.mult1_un61_sum_cry_4_s ));
    InMux I__1785 (
            .O(N__16412),
            .I(\b2v_inst11.mult1_un61_sum_cry_3 ));
    CascadeMux I__1784 (
            .O(N__16409),
            .I(N__16406));
    InMux I__1783 (
            .O(N__16406),
            .I(N__16403));
    LocalMux I__1782 (
            .O(N__16403),
            .I(\b2v_inst11.mult1_un61_sum_cry_5_s ));
    InMux I__1781 (
            .O(N__16400),
            .I(\b2v_inst11.mult1_un61_sum_cry_4 ));
    InMux I__1780 (
            .O(N__16397),
            .I(N__16394));
    LocalMux I__1779 (
            .O(N__16394),
            .I(\b2v_inst11.mult1_un61_sum_cry_6_s ));
    InMux I__1778 (
            .O(N__16391),
            .I(\b2v_inst11.mult1_un61_sum_cry_5 ));
    InMux I__1777 (
            .O(N__16388),
            .I(N__16382));
    InMux I__1776 (
            .O(N__16387),
            .I(N__16382));
    LocalMux I__1775 (
            .O(N__16382),
            .I(\b2v_inst200.count_3_9 ));
    CascadeMux I__1774 (
            .O(N__16379),
            .I(\b2v_inst200.countZ0Z_12_cascade_ ));
    InMux I__1773 (
            .O(N__16376),
            .I(N__16367));
    InMux I__1772 (
            .O(N__16375),
            .I(N__16367));
    InMux I__1771 (
            .O(N__16374),
            .I(N__16367));
    LocalMux I__1770 (
            .O(N__16367),
            .I(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ));
    InMux I__1769 (
            .O(N__16364),
            .I(N__16361));
    LocalMux I__1768 (
            .O(N__16361),
            .I(\b2v_inst200.un2_count_1_axb_5 ));
    InMux I__1767 (
            .O(N__16358),
            .I(N__16355));
    LocalMux I__1766 (
            .O(N__16355),
            .I(N__16352));
    Odrv4 I__1765 (
            .O(N__16352),
            .I(\b2v_inst200.count_3_11 ));
    InMux I__1764 (
            .O(N__16349),
            .I(N__16346));
    LocalMux I__1763 (
            .O(N__16346),
            .I(N__16342));
    InMux I__1762 (
            .O(N__16345),
            .I(N__16339));
    Odrv4 I__1761 (
            .O(N__16342),
            .I(\b2v_inst200.count_1_11 ));
    LocalMux I__1760 (
            .O(N__16339),
            .I(\b2v_inst200.count_1_11 ));
    InMux I__1759 (
            .O(N__16334),
            .I(N__16331));
    LocalMux I__1758 (
            .O(N__16331),
            .I(N__16328));
    Span4Mux_s1_h I__1757 (
            .O(N__16328),
            .I(N__16324));
    InMux I__1756 (
            .O(N__16327),
            .I(N__16321));
    Odrv4 I__1755 (
            .O(N__16324),
            .I(\b2v_inst200.countZ0Z_11 ));
    LocalMux I__1754 (
            .O(N__16321),
            .I(\b2v_inst200.countZ0Z_11 ));
    InMux I__1753 (
            .O(N__16316),
            .I(N__16313));
    LocalMux I__1752 (
            .O(N__16313),
            .I(N__16310));
    Odrv4 I__1751 (
            .O(N__16310),
            .I(\b2v_inst200.un2_count_1_axb_3 ));
    CascadeMux I__1750 (
            .O(N__16307),
            .I(N__16304));
    InMux I__1749 (
            .O(N__16304),
            .I(N__16300));
    InMux I__1748 (
            .O(N__16303),
            .I(N__16297));
    LocalMux I__1747 (
            .O(N__16300),
            .I(N__16292));
    LocalMux I__1746 (
            .O(N__16297),
            .I(N__16292));
    Odrv4 I__1745 (
            .O(N__16292),
            .I(\b2v_inst200.countZ0Z_14 ));
    InMux I__1744 (
            .O(N__16289),
            .I(N__16286));
    LocalMux I__1743 (
            .O(N__16286),
            .I(\b2v_inst200.un25_clk_100khz_4 ));
    CascadeMux I__1742 (
            .O(N__16283),
            .I(\b2v_inst200.un25_clk_100khz_5_cascade_ ));
    InMux I__1741 (
            .O(N__16280),
            .I(N__16277));
    LocalMux I__1740 (
            .O(N__16277),
            .I(N__16274));
    Odrv4 I__1739 (
            .O(N__16274),
            .I(\b2v_inst200.un25_clk_100khz_14 ));
    InMux I__1738 (
            .O(N__16271),
            .I(N__16265));
    InMux I__1737 (
            .O(N__16270),
            .I(N__16265));
    LocalMux I__1736 (
            .O(N__16265),
            .I(\b2v_inst200.count_3_3 ));
    CascadeMux I__1735 (
            .O(N__16262),
            .I(N__16259));
    InMux I__1734 (
            .O(N__16259),
            .I(N__16256));
    LocalMux I__1733 (
            .O(N__16256),
            .I(N__16252));
    InMux I__1732 (
            .O(N__16255),
            .I(N__16249));
    Span12Mux_v I__1731 (
            .O(N__16252),
            .I(N__16246));
    LocalMux I__1730 (
            .O(N__16249),
            .I(N__16243));
    Odrv12 I__1729 (
            .O(N__16246),
            .I(\b2v_inst200.countZ0Z_4 ));
    Odrv4 I__1728 (
            .O(N__16243),
            .I(\b2v_inst200.countZ0Z_4 ));
    InMux I__1727 (
            .O(N__16238),
            .I(N__16229));
    InMux I__1726 (
            .O(N__16237),
            .I(N__16229));
    InMux I__1725 (
            .O(N__16236),
            .I(N__16229));
    LocalMux I__1724 (
            .O(N__16229),
            .I(N__16226));
    Odrv4 I__1723 (
            .O(N__16226),
            .I(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ));
    InMux I__1722 (
            .O(N__16223),
            .I(N__16220));
    LocalMux I__1721 (
            .O(N__16220),
            .I(\b2v_inst200.un25_clk_100khz_2 ));
    InMux I__1720 (
            .O(N__16217),
            .I(N__16208));
    InMux I__1719 (
            .O(N__16216),
            .I(N__16208));
    InMux I__1718 (
            .O(N__16215),
            .I(N__16208));
    LocalMux I__1717 (
            .O(N__16208),
            .I(\b2v_inst200.count_1_8 ));
    CascadeMux I__1716 (
            .O(N__16205),
            .I(N__16202));
    InMux I__1715 (
            .O(N__16202),
            .I(N__16196));
    InMux I__1714 (
            .O(N__16201),
            .I(N__16196));
    LocalMux I__1713 (
            .O(N__16196),
            .I(\b2v_inst200.count_3_8 ));
    InMux I__1712 (
            .O(N__16193),
            .I(N__16190));
    LocalMux I__1711 (
            .O(N__16190),
            .I(\b2v_inst200.un2_count_1_axb_8 ));
    InMux I__1710 (
            .O(N__16187),
            .I(N__16184));
    LocalMux I__1709 (
            .O(N__16184),
            .I(\b2v_inst200.un2_count_1_axb_15 ));
    InMux I__1708 (
            .O(N__16181),
            .I(N__16175));
    InMux I__1707 (
            .O(N__16180),
            .I(N__16175));
    LocalMux I__1706 (
            .O(N__16175),
            .I(\b2v_inst200.count_3_15 ));
    CascadeMux I__1705 (
            .O(N__16172),
            .I(N__16167));
    InMux I__1704 (
            .O(N__16171),
            .I(N__16160));
    InMux I__1703 (
            .O(N__16170),
            .I(N__16160));
    InMux I__1702 (
            .O(N__16167),
            .I(N__16160));
    LocalMux I__1701 (
            .O(N__16160),
            .I(\b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71 ));
    CascadeMux I__1700 (
            .O(N__16157),
            .I(N__16153));
    CascadeMux I__1699 (
            .O(N__16156),
            .I(N__16150));
    InMux I__1698 (
            .O(N__16153),
            .I(N__16147));
    InMux I__1697 (
            .O(N__16150),
            .I(N__16144));
    LocalMux I__1696 (
            .O(N__16147),
            .I(\b2v_inst200.countZ0Z_6 ));
    LocalMux I__1695 (
            .O(N__16144),
            .I(\b2v_inst200.countZ0Z_6 ));
    InMux I__1694 (
            .O(N__16139),
            .I(N__16136));
    LocalMux I__1693 (
            .O(N__16136),
            .I(\b2v_inst200.un25_clk_100khz_7 ));
    InMux I__1692 (
            .O(N__16133),
            .I(N__16130));
    LocalMux I__1691 (
            .O(N__16130),
            .I(N__16127));
    Span4Mux_v I__1690 (
            .O(N__16127),
            .I(N__16124));
    Odrv4 I__1689 (
            .O(N__16124),
            .I(\b2v_inst200.un25_clk_100khz_13 ));
    CascadeMux I__1688 (
            .O(N__16121),
            .I(\b2v_inst200.un25_clk_100khz_6_cascade_ ));
    CascadeMux I__1687 (
            .O(N__16118),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_ ));
    InMux I__1686 (
            .O(N__16115),
            .I(N__16111));
    CascadeMux I__1685 (
            .O(N__16114),
            .I(N__16107));
    LocalMux I__1684 (
            .O(N__16111),
            .I(N__16101));
    InMux I__1683 (
            .O(N__16110),
            .I(N__16098));
    InMux I__1682 (
            .O(N__16107),
            .I(N__16095));
    InMux I__1681 (
            .O(N__16106),
            .I(N__16088));
    InMux I__1680 (
            .O(N__16105),
            .I(N__16088));
    InMux I__1679 (
            .O(N__16104),
            .I(N__16088));
    Odrv4 I__1678 (
            .O(N__16101),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__1677 (
            .O(N__16098),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__1676 (
            .O(N__16095),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__1675 (
            .O(N__16088),
            .I(\b2v_inst200.countZ0Z_0 ));
    InMux I__1674 (
            .O(N__16079),
            .I(N__16076));
    LocalMux I__1673 (
            .O(N__16076),
            .I(\b2v_inst200.count_3_0 ));
    InMux I__1672 (
            .O(N__16073),
            .I(N__16070));
    LocalMux I__1671 (
            .O(N__16070),
            .I(\b2v_inst200.un2_count_1_axb_9 ));
    InMux I__1670 (
            .O(N__16067),
            .I(N__16064));
    LocalMux I__1669 (
            .O(N__16064),
            .I(\b2v_inst200.count_3_12 ));
    InMux I__1668 (
            .O(N__16061),
            .I(N__16055));
    InMux I__1667 (
            .O(N__16060),
            .I(N__16055));
    LocalMux I__1666 (
            .O(N__16055),
            .I(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ));
    InMux I__1665 (
            .O(N__16052),
            .I(N__16049));
    LocalMux I__1664 (
            .O(N__16049),
            .I(\b2v_inst200.countZ0Z_12 ));
    InMux I__1663 (
            .O(N__16046),
            .I(N__16043));
    LocalMux I__1662 (
            .O(N__16043),
            .I(\b2v_inst200.count_3_6 ));
    InMux I__1661 (
            .O(N__16040),
            .I(N__16036));
    InMux I__1660 (
            .O(N__16039),
            .I(N__16033));
    LocalMux I__1659 (
            .O(N__16036),
            .I(\b2v_inst200.count_1_6 ));
    LocalMux I__1658 (
            .O(N__16033),
            .I(\b2v_inst200.count_1_6 ));
    InMux I__1657 (
            .O(N__16028),
            .I(N__16025));
    LocalMux I__1656 (
            .O(N__16025),
            .I(\b2v_inst200.count_3_7 ));
    InMux I__1655 (
            .O(N__16022),
            .I(N__16018));
    InMux I__1654 (
            .O(N__16021),
            .I(N__16015));
    LocalMux I__1653 (
            .O(N__16018),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    LocalMux I__1652 (
            .O(N__16015),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    InMux I__1651 (
            .O(N__16010),
            .I(N__16007));
    LocalMux I__1650 (
            .O(N__16007),
            .I(N__16004));
    Span4Mux_h I__1649 (
            .O(N__16004),
            .I(N__16001));
    Odrv4 I__1648 (
            .O(N__16001),
            .I(\b2v_inst200.count_0_17 ));
    InMux I__1647 (
            .O(N__15998),
            .I(N__15995));
    LocalMux I__1646 (
            .O(N__15995),
            .I(N__15991));
    InMux I__1645 (
            .O(N__15994),
            .I(N__15988));
    Span4Mux_h I__1644 (
            .O(N__15991),
            .I(N__15985));
    LocalMux I__1643 (
            .O(N__15988),
            .I(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ));
    Odrv4 I__1642 (
            .O(N__15985),
            .I(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ));
    InMux I__1641 (
            .O(N__15980),
            .I(N__15977));
    LocalMux I__1640 (
            .O(N__15977),
            .I(N__15973));
    InMux I__1639 (
            .O(N__15976),
            .I(N__15970));
    Odrv4 I__1638 (
            .O(N__15973),
            .I(\b2v_inst200.countZ0Z_17 ));
    LocalMux I__1637 (
            .O(N__15970),
            .I(\b2v_inst200.countZ0Z_17 ));
    CascadeMux I__1636 (
            .O(N__15965),
            .I(N__15961));
    InMux I__1635 (
            .O(N__15964),
            .I(N__15958));
    InMux I__1634 (
            .O(N__15961),
            .I(N__15955));
    LocalMux I__1633 (
            .O(N__15958),
            .I(N__15950));
    LocalMux I__1632 (
            .O(N__15955),
            .I(N__15950));
    Odrv4 I__1631 (
            .O(N__15950),
            .I(\b2v_inst200.count_1_10 ));
    InMux I__1630 (
            .O(N__15947),
            .I(N__15944));
    LocalMux I__1629 (
            .O(N__15944),
            .I(N__15941));
    Odrv4 I__1628 (
            .O(N__15941),
            .I(\b2v_inst200.count_3_10 ));
    InMux I__1627 (
            .O(N__15938),
            .I(N__15935));
    LocalMux I__1626 (
            .O(N__15935),
            .I(N__15932));
    Odrv4 I__1625 (
            .O(N__15932),
            .I(\b2v_inst200.count_1_0 ));
    CascadeMux I__1624 (
            .O(N__15929),
            .I(N__15926));
    InMux I__1623 (
            .O(N__15926),
            .I(N__15922));
    InMux I__1622 (
            .O(N__15925),
            .I(N__15919));
    LocalMux I__1621 (
            .O(N__15922),
            .I(N__15916));
    LocalMux I__1620 (
            .O(N__15919),
            .I(\b2v_inst200.countZ0Z_10 ));
    Odrv4 I__1619 (
            .O(N__15916),
            .I(\b2v_inst200.countZ0Z_10 ));
    InMux I__1618 (
            .O(N__15911),
            .I(N__15906));
    InMux I__1617 (
            .O(N__15910),
            .I(N__15901));
    InMux I__1616 (
            .O(N__15909),
            .I(N__15901));
    LocalMux I__1615 (
            .O(N__15906),
            .I(N__15898));
    LocalMux I__1614 (
            .O(N__15901),
            .I(\b2v_inst16.countZ0Z_11 ));
    Odrv4 I__1613 (
            .O(N__15898),
            .I(\b2v_inst16.countZ0Z_11 ));
    InMux I__1612 (
            .O(N__15893),
            .I(N__15887));
    InMux I__1611 (
            .O(N__15892),
            .I(N__15887));
    LocalMux I__1610 (
            .O(N__15887),
            .I(N__15884));
    Odrv4 I__1609 (
            .O(N__15884),
            .I(\b2v_inst16.un4_count_1_cry_10_THRU_CO ));
    InMux I__1608 (
            .O(N__15881),
            .I(\b2v_inst16.un4_count_1_cry_10 ));
    InMux I__1607 (
            .O(N__15878),
            .I(\b2v_inst16.un4_count_1_cry_11 ));
    InMux I__1606 (
            .O(N__15875),
            .I(\b2v_inst16.un4_count_1_cry_12 ));
    InMux I__1605 (
            .O(N__15872),
            .I(\b2v_inst16.un4_count_1_cry_13 ));
    InMux I__1604 (
            .O(N__15869),
            .I(N__15866));
    LocalMux I__1603 (
            .O(N__15866),
            .I(N__15862));
    InMux I__1602 (
            .O(N__15865),
            .I(N__15859));
    Odrv4 I__1601 (
            .O(N__15862),
            .I(\b2v_inst16.countZ0Z_15 ));
    LocalMux I__1600 (
            .O(N__15859),
            .I(\b2v_inst16.countZ0Z_15 ));
    InMux I__1599 (
            .O(N__15854),
            .I(\b2v_inst16.un4_count_1_cry_14 ));
    InMux I__1598 (
            .O(N__15851),
            .I(N__15847));
    InMux I__1597 (
            .O(N__15850),
            .I(N__15844));
    LocalMux I__1596 (
            .O(N__15847),
            .I(\b2v_inst16.count_rst_4 ));
    LocalMux I__1595 (
            .O(N__15844),
            .I(\b2v_inst16.count_rst_4 ));
    InMux I__1594 (
            .O(N__15839),
            .I(N__15836));
    LocalMux I__1593 (
            .O(N__15836),
            .I(\b2v_inst200.count_3_14 ));
    InMux I__1592 (
            .O(N__15833),
            .I(N__15829));
    InMux I__1591 (
            .O(N__15832),
            .I(N__15826));
    LocalMux I__1590 (
            .O(N__15829),
            .I(N__15821));
    LocalMux I__1589 (
            .O(N__15826),
            .I(N__15821));
    Odrv4 I__1588 (
            .O(N__15821),
            .I(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ));
    InMux I__1587 (
            .O(N__15818),
            .I(\b2v_inst16.un4_count_1_cry_1 ));
    InMux I__1586 (
            .O(N__15815),
            .I(\b2v_inst16.un4_count_1_cry_2 ));
    CascadeMux I__1585 (
            .O(N__15812),
            .I(N__15809));
    InMux I__1584 (
            .O(N__15809),
            .I(N__15804));
    InMux I__1583 (
            .O(N__15808),
            .I(N__15801));
    InMux I__1582 (
            .O(N__15807),
            .I(N__15798));
    LocalMux I__1581 (
            .O(N__15804),
            .I(N__15795));
    LocalMux I__1580 (
            .O(N__15801),
            .I(N__15790));
    LocalMux I__1579 (
            .O(N__15798),
            .I(N__15790));
    Odrv4 I__1578 (
            .O(N__15795),
            .I(\b2v_inst16.countZ0Z_4 ));
    Odrv4 I__1577 (
            .O(N__15790),
            .I(\b2v_inst16.countZ0Z_4 ));
    InMux I__1576 (
            .O(N__15785),
            .I(N__15779));
    InMux I__1575 (
            .O(N__15784),
            .I(N__15779));
    LocalMux I__1574 (
            .O(N__15779),
            .I(N__15776));
    Odrv4 I__1573 (
            .O(N__15776),
            .I(\b2v_inst16.un4_count_1_cry_3_THRU_CO ));
    InMux I__1572 (
            .O(N__15773),
            .I(\b2v_inst16.un4_count_1_cry_3 ));
    InMux I__1571 (
            .O(N__15770),
            .I(N__15765));
    InMux I__1570 (
            .O(N__15769),
            .I(N__15762));
    InMux I__1569 (
            .O(N__15768),
            .I(N__15759));
    LocalMux I__1568 (
            .O(N__15765),
            .I(N__15756));
    LocalMux I__1567 (
            .O(N__15762),
            .I(\b2v_inst16.countZ0Z_5 ));
    LocalMux I__1566 (
            .O(N__15759),
            .I(\b2v_inst16.countZ0Z_5 ));
    Odrv4 I__1565 (
            .O(N__15756),
            .I(\b2v_inst16.countZ0Z_5 ));
    InMux I__1564 (
            .O(N__15749),
            .I(N__15743));
    InMux I__1563 (
            .O(N__15748),
            .I(N__15743));
    LocalMux I__1562 (
            .O(N__15743),
            .I(N__15740));
    Odrv4 I__1561 (
            .O(N__15740),
            .I(\b2v_inst16.un4_count_1_cry_4_THRU_CO ));
    InMux I__1560 (
            .O(N__15737),
            .I(\b2v_inst16.un4_count_1_cry_4 ));
    InMux I__1559 (
            .O(N__15734),
            .I(N__15730));
    InMux I__1558 (
            .O(N__15733),
            .I(N__15727));
    LocalMux I__1557 (
            .O(N__15730),
            .I(\b2v_inst16.countZ0Z_6 ));
    LocalMux I__1556 (
            .O(N__15727),
            .I(\b2v_inst16.countZ0Z_6 ));
    InMux I__1555 (
            .O(N__15722),
            .I(N__15716));
    InMux I__1554 (
            .O(N__15721),
            .I(N__15716));
    LocalMux I__1553 (
            .O(N__15716),
            .I(\b2v_inst16.count_rst_11 ));
    InMux I__1552 (
            .O(N__15713),
            .I(\b2v_inst16.un4_count_1_cry_5 ));
    CascadeMux I__1551 (
            .O(N__15710),
            .I(N__15705));
    InMux I__1550 (
            .O(N__15709),
            .I(N__15701));
    InMux I__1549 (
            .O(N__15708),
            .I(N__15698));
    InMux I__1548 (
            .O(N__15705),
            .I(N__15695));
    InMux I__1547 (
            .O(N__15704),
            .I(N__15692));
    LocalMux I__1546 (
            .O(N__15701),
            .I(N__15689));
    LocalMux I__1545 (
            .O(N__15698),
            .I(\b2v_inst16.countZ0Z_7 ));
    LocalMux I__1544 (
            .O(N__15695),
            .I(\b2v_inst16.countZ0Z_7 ));
    LocalMux I__1543 (
            .O(N__15692),
            .I(\b2v_inst16.countZ0Z_7 ));
    Odrv4 I__1542 (
            .O(N__15689),
            .I(\b2v_inst16.countZ0Z_7 ));
    InMux I__1541 (
            .O(N__15680),
            .I(N__15676));
    InMux I__1540 (
            .O(N__15679),
            .I(N__15673));
    LocalMux I__1539 (
            .O(N__15676),
            .I(N__15668));
    LocalMux I__1538 (
            .O(N__15673),
            .I(N__15668));
    Odrv4 I__1537 (
            .O(N__15668),
            .I(\b2v_inst16.un4_count_1_cry_6_THRU_CO ));
    InMux I__1536 (
            .O(N__15665),
            .I(\b2v_inst16.un4_count_1_cry_6 ));
    CascadeMux I__1535 (
            .O(N__15662),
            .I(N__15658));
    InMux I__1534 (
            .O(N__15661),
            .I(N__15653));
    InMux I__1533 (
            .O(N__15658),
            .I(N__15650));
    InMux I__1532 (
            .O(N__15657),
            .I(N__15645));
    InMux I__1531 (
            .O(N__15656),
            .I(N__15645));
    LocalMux I__1530 (
            .O(N__15653),
            .I(N__15642));
    LocalMux I__1529 (
            .O(N__15650),
            .I(\b2v_inst16.countZ0Z_8 ));
    LocalMux I__1528 (
            .O(N__15645),
            .I(\b2v_inst16.countZ0Z_8 ));
    Odrv4 I__1527 (
            .O(N__15642),
            .I(\b2v_inst16.countZ0Z_8 ));
    CascadeMux I__1526 (
            .O(N__15635),
            .I(N__15631));
    InMux I__1525 (
            .O(N__15634),
            .I(N__15628));
    InMux I__1524 (
            .O(N__15631),
            .I(N__15625));
    LocalMux I__1523 (
            .O(N__15628),
            .I(N__15622));
    LocalMux I__1522 (
            .O(N__15625),
            .I(\b2v_inst16.un4_count_1_cry_7_THRU_CO ));
    Odrv4 I__1521 (
            .O(N__15622),
            .I(\b2v_inst16.un4_count_1_cry_7_THRU_CO ));
    InMux I__1520 (
            .O(N__15617),
            .I(\b2v_inst16.un4_count_1_cry_7 ));
    InMux I__1519 (
            .O(N__15614),
            .I(N__15609));
    InMux I__1518 (
            .O(N__15613),
            .I(N__15606));
    InMux I__1517 (
            .O(N__15612),
            .I(N__15603));
    LocalMux I__1516 (
            .O(N__15609),
            .I(N__15598));
    LocalMux I__1515 (
            .O(N__15606),
            .I(N__15598));
    LocalMux I__1514 (
            .O(N__15603),
            .I(\b2v_inst16.countZ0Z_9 ));
    Odrv4 I__1513 (
            .O(N__15598),
            .I(\b2v_inst16.countZ0Z_9 ));
    CascadeMux I__1512 (
            .O(N__15593),
            .I(N__15589));
    InMux I__1511 (
            .O(N__15592),
            .I(N__15586));
    InMux I__1510 (
            .O(N__15589),
            .I(N__15583));
    LocalMux I__1509 (
            .O(N__15586),
            .I(N__15578));
    LocalMux I__1508 (
            .O(N__15583),
            .I(N__15578));
    Span4Mux_s1_h I__1507 (
            .O(N__15578),
            .I(N__15575));
    Odrv4 I__1506 (
            .O(N__15575),
            .I(\b2v_inst16.un4_count_1_cry_8_THRU_CO ));
    InMux I__1505 (
            .O(N__15572),
            .I(bfn_2_4_0_));
    InMux I__1504 (
            .O(N__15569),
            .I(\b2v_inst16.un4_count_1_cry_9 ));
    CascadeMux I__1503 (
            .O(N__15566),
            .I(\b2v_inst16.countZ0Z_2_cascade_ ));
    InMux I__1502 (
            .O(N__15563),
            .I(N__15560));
    LocalMux I__1501 (
            .O(N__15560),
            .I(\b2v_inst16.count_4_i_a3_8_0 ));
    CascadeMux I__1500 (
            .O(N__15557),
            .I(\b2v_inst16.count_4_i_a3_9_0_cascade_ ));
    InMux I__1499 (
            .O(N__15554),
            .I(N__15551));
    LocalMux I__1498 (
            .O(N__15551),
            .I(\b2v_inst16.count_4_i_a3_7_0 ));
    InMux I__1497 (
            .O(N__15548),
            .I(N__15545));
    LocalMux I__1496 (
            .O(N__15545),
            .I(\b2v_inst16.count_rst_5 ));
    CascadeMux I__1495 (
            .O(N__15542),
            .I(\b2v_inst16.countZ0Z_0_cascade_ ));
    InMux I__1494 (
            .O(N__15539),
            .I(N__15534));
    InMux I__1493 (
            .O(N__15538),
            .I(N__15531));
    InMux I__1492 (
            .O(N__15537),
            .I(N__15528));
    LocalMux I__1491 (
            .O(N__15534),
            .I(\b2v_inst16.N_414 ));
    LocalMux I__1490 (
            .O(N__15531),
            .I(\b2v_inst16.N_414 ));
    LocalMux I__1489 (
            .O(N__15528),
            .I(\b2v_inst16.N_414 ));
    InMux I__1488 (
            .O(N__15521),
            .I(N__15518));
    LocalMux I__1487 (
            .O(N__15518),
            .I(\b2v_inst16.count_4_0 ));
    CascadeMux I__1486 (
            .O(N__15515),
            .I(N__15512));
    InMux I__1485 (
            .O(N__15512),
            .I(N__15506));
    InMux I__1484 (
            .O(N__15511),
            .I(N__15506));
    LocalMux I__1483 (
            .O(N__15506),
            .I(\b2v_inst16.count_4_2 ));
    InMux I__1482 (
            .O(N__15503),
            .I(N__15494));
    InMux I__1481 (
            .O(N__15502),
            .I(N__15494));
    InMux I__1480 (
            .O(N__15501),
            .I(N__15491));
    InMux I__1479 (
            .O(N__15500),
            .I(N__15486));
    InMux I__1478 (
            .O(N__15499),
            .I(N__15486));
    LocalMux I__1477 (
            .O(N__15494),
            .I(\b2v_inst16.countZ0Z_0 ));
    LocalMux I__1476 (
            .O(N__15491),
            .I(\b2v_inst16.countZ0Z_0 ));
    LocalMux I__1475 (
            .O(N__15486),
            .I(\b2v_inst16.countZ0Z_0 ));
    CascadeMux I__1474 (
            .O(N__15479),
            .I(N__15474));
    InMux I__1473 (
            .O(N__15478),
            .I(N__15469));
    InMux I__1472 (
            .O(N__15477),
            .I(N__15469));
    InMux I__1471 (
            .O(N__15474),
            .I(N__15466));
    LocalMux I__1470 (
            .O(N__15469),
            .I(\b2v_inst16.countZ0Z_1 ));
    LocalMux I__1469 (
            .O(N__15466),
            .I(\b2v_inst16.countZ0Z_1 ));
    CascadeMux I__1468 (
            .O(N__15461),
            .I(N__15458));
    InMux I__1467 (
            .O(N__15458),
            .I(N__15455));
    LocalMux I__1466 (
            .O(N__15455),
            .I(\b2v_inst16.un4_count_1_axb_2 ));
    CascadeMux I__1465 (
            .O(N__15452),
            .I(N__15448));
    InMux I__1464 (
            .O(N__15451),
            .I(N__15440));
    InMux I__1463 (
            .O(N__15448),
            .I(N__15440));
    InMux I__1462 (
            .O(N__15447),
            .I(N__15440));
    LocalMux I__1461 (
            .O(N__15440),
            .I(\b2v_inst16.un4_count_1_cry_1_c_RNIAGMEZ0 ));
    InMux I__1460 (
            .O(N__15437),
            .I(\b2v_inst11.un1_count_cry_14 ));
    CascadeMux I__1459 (
            .O(N__15434),
            .I(\b2v_inst16.count_rst_9_cascade_ ));
    CascadeMux I__1458 (
            .O(N__15431),
            .I(\b2v_inst16.countZ0Z_4_cascade_ ));
    InMux I__1457 (
            .O(N__15428),
            .I(N__15425));
    LocalMux I__1456 (
            .O(N__15425),
            .I(\b2v_inst16.count_4_4 ));
    CascadeMux I__1455 (
            .O(N__15422),
            .I(\b2v_inst16.count_rst_10_cascade_ ));
    CascadeMux I__1454 (
            .O(N__15419),
            .I(\b2v_inst16.countZ0Z_5_cascade_ ));
    InMux I__1453 (
            .O(N__15416),
            .I(N__15413));
    LocalMux I__1452 (
            .O(N__15413),
            .I(\b2v_inst16.count_4_5 ));
    InMux I__1451 (
            .O(N__15410),
            .I(N__15407));
    LocalMux I__1450 (
            .O(N__15407),
            .I(\b2v_inst16.count_4_7 ));
    InMux I__1449 (
            .O(N__15404),
            .I(\b2v_inst11.un1_count_cry_6 ));
    CascadeMux I__1448 (
            .O(N__15401),
            .I(N__15398));
    InMux I__1447 (
            .O(N__15398),
            .I(N__15392));
    InMux I__1446 (
            .O(N__15397),
            .I(N__15392));
    LocalMux I__1445 (
            .O(N__15392),
            .I(N__15389));
    Odrv4 I__1444 (
            .O(N__15389),
            .I(\b2v_inst11.count_1_8 ));
    InMux I__1443 (
            .O(N__15386),
            .I(\b2v_inst11.un1_count_cry_7 ));
    CascadeMux I__1442 (
            .O(N__15383),
            .I(N__15380));
    InMux I__1441 (
            .O(N__15380),
            .I(N__15374));
    InMux I__1440 (
            .O(N__15379),
            .I(N__15374));
    LocalMux I__1439 (
            .O(N__15374),
            .I(N__15371));
    Odrv4 I__1438 (
            .O(N__15371),
            .I(\b2v_inst11.count_1_9 ));
    InMux I__1437 (
            .O(N__15368),
            .I(bfn_1_16_0_));
    InMux I__1436 (
            .O(N__15365),
            .I(N__15359));
    InMux I__1435 (
            .O(N__15364),
            .I(N__15359));
    LocalMux I__1434 (
            .O(N__15359),
            .I(N__15356));
    Odrv4 I__1433 (
            .O(N__15356),
            .I(\b2v_inst11.count_1_10 ));
    InMux I__1432 (
            .O(N__15353),
            .I(\b2v_inst11.un1_count_cry_9 ));
    InMux I__1431 (
            .O(N__15350),
            .I(N__15344));
    InMux I__1430 (
            .O(N__15349),
            .I(N__15344));
    LocalMux I__1429 (
            .O(N__15344),
            .I(N__15341));
    Odrv4 I__1428 (
            .O(N__15341),
            .I(\b2v_inst11.count_1_11 ));
    InMux I__1427 (
            .O(N__15338),
            .I(\b2v_inst11.un1_count_cry_10 ));
    InMux I__1426 (
            .O(N__15335),
            .I(N__15329));
    InMux I__1425 (
            .O(N__15334),
            .I(N__15329));
    LocalMux I__1424 (
            .O(N__15329),
            .I(N__15326));
    Odrv4 I__1423 (
            .O(N__15326),
            .I(\b2v_inst11.count_1_12 ));
    InMux I__1422 (
            .O(N__15323),
            .I(\b2v_inst11.un1_count_cry_11 ));
    InMux I__1421 (
            .O(N__15320),
            .I(\b2v_inst11.un1_count_cry_12 ));
    InMux I__1420 (
            .O(N__15317),
            .I(\b2v_inst11.un1_count_cry_13 ));
    InMux I__1419 (
            .O(N__15314),
            .I(N__15311));
    LocalMux I__1418 (
            .O(N__15311),
            .I(\b2v_inst11.count_0_2 ));
    InMux I__1417 (
            .O(N__15308),
            .I(N__15305));
    LocalMux I__1416 (
            .O(N__15305),
            .I(\b2v_inst11.count_0_12 ));
    CascadeMux I__1415 (
            .O(N__15302),
            .I(N__15298));
    InMux I__1414 (
            .O(N__15301),
            .I(N__15293));
    InMux I__1413 (
            .O(N__15298),
            .I(N__15293));
    LocalMux I__1412 (
            .O(N__15293),
            .I(\b2v_inst11.count_1_2 ));
    InMux I__1411 (
            .O(N__15290),
            .I(\b2v_inst11.un1_count_cry_1_cZ0 ));
    InMux I__1410 (
            .O(N__15287),
            .I(\b2v_inst11.un1_count_cry_2 ));
    InMux I__1409 (
            .O(N__15284),
            .I(\b2v_inst11.un1_count_cry_3 ));
    InMux I__1408 (
            .O(N__15281),
            .I(\b2v_inst11.un1_count_cry_4 ));
    InMux I__1407 (
            .O(N__15278),
            .I(\b2v_inst11.un1_count_cry_5 ));
    InMux I__1406 (
            .O(N__15275),
            .I(N__15272));
    LocalMux I__1405 (
            .O(N__15272),
            .I(\b2v_inst11.count_0_9 ));
    InMux I__1404 (
            .O(N__15269),
            .I(N__15266));
    LocalMux I__1403 (
            .O(N__15266),
            .I(\b2v_inst11.count_0_10 ));
    InMux I__1402 (
            .O(N__15263),
            .I(N__15260));
    LocalMux I__1401 (
            .O(N__15260),
            .I(\b2v_inst11.count_0_11 ));
    CascadeMux I__1400 (
            .O(N__15257),
            .I(\b2v_inst11.count_1_1_cascade_ ));
    CascadeMux I__1399 (
            .O(N__15254),
            .I(\b2v_inst11.countZ0Z_1_cascade_ ));
    InMux I__1398 (
            .O(N__15251),
            .I(N__15248));
    LocalMux I__1397 (
            .O(N__15248),
            .I(\b2v_inst11.count_0_1 ));
    CascadeMux I__1396 (
            .O(N__15245),
            .I(N__15242));
    InMux I__1395 (
            .O(N__15242),
            .I(N__15239));
    LocalMux I__1394 (
            .O(N__15239),
            .I(\b2v_inst11.mult1_un89_sum_cry_3_s ));
    InMux I__1393 (
            .O(N__15236),
            .I(\b2v_inst11.mult1_un96_sum_cry_3 ));
    InMux I__1392 (
            .O(N__15233),
            .I(N__15230));
    LocalMux I__1391 (
            .O(N__15230),
            .I(\b2v_inst11.mult1_un89_sum_cry_4_s ));
    InMux I__1390 (
            .O(N__15227),
            .I(\b2v_inst11.mult1_un96_sum_cry_4 ));
    CascadeMux I__1389 (
            .O(N__15224),
            .I(N__15221));
    InMux I__1388 (
            .O(N__15221),
            .I(N__15218));
    LocalMux I__1387 (
            .O(N__15218),
            .I(\b2v_inst11.mult1_un89_sum_cry_5_s ));
    InMux I__1386 (
            .O(N__15215),
            .I(\b2v_inst11.mult1_un96_sum_cry_5 ));
    InMux I__1385 (
            .O(N__15212),
            .I(N__15209));
    LocalMux I__1384 (
            .O(N__15209),
            .I(\b2v_inst11.mult1_un89_sum_cry_6_s ));
    CascadeMux I__1383 (
            .O(N__15206),
            .I(N__15202));
    CascadeMux I__1382 (
            .O(N__15205),
            .I(N__15198));
    InMux I__1381 (
            .O(N__15202),
            .I(N__15191));
    InMux I__1380 (
            .O(N__15201),
            .I(N__15191));
    InMux I__1379 (
            .O(N__15198),
            .I(N__15191));
    LocalMux I__1378 (
            .O(N__15191),
            .I(\b2v_inst11.mult1_un89_sum_i_0_8 ));
    InMux I__1377 (
            .O(N__15188),
            .I(\b2v_inst11.mult1_un96_sum_cry_6 ));
    CascadeMux I__1376 (
            .O(N__15185),
            .I(N__15182));
    InMux I__1375 (
            .O(N__15182),
            .I(N__15179));
    LocalMux I__1374 (
            .O(N__15179),
            .I(\b2v_inst11.mult1_un96_sum_axb_8 ));
    InMux I__1373 (
            .O(N__15176),
            .I(\b2v_inst11.mult1_un96_sum_cry_7 ));
    CascadeMux I__1372 (
            .O(N__15173),
            .I(\b2v_inst11.mult1_un96_sum_s_8_cascade_ ));
    InMux I__1371 (
            .O(N__15170),
            .I(N__15167));
    LocalMux I__1370 (
            .O(N__15167),
            .I(\b2v_inst11.count_0_8 ));
    InMux I__1369 (
            .O(N__15164),
            .I(\b2v_inst11.mult1_un89_sum_cry_2 ));
    InMux I__1368 (
            .O(N__15161),
            .I(\b2v_inst11.mult1_un89_sum_cry_3 ));
    InMux I__1367 (
            .O(N__15158),
            .I(\b2v_inst11.mult1_un89_sum_cry_4 ));
    InMux I__1366 (
            .O(N__15155),
            .I(\b2v_inst11.mult1_un89_sum_cry_5 ));
    InMux I__1365 (
            .O(N__15152),
            .I(\b2v_inst11.mult1_un89_sum_cry_6 ));
    InMux I__1364 (
            .O(N__15149),
            .I(\b2v_inst11.mult1_un89_sum_cry_7 ));
    CascadeMux I__1363 (
            .O(N__15146),
            .I(\b2v_inst11.mult1_un89_sum_s_8_cascade_ ));
    InMux I__1362 (
            .O(N__15143),
            .I(\b2v_inst11.mult1_un96_sum_cry_2 ));
    InMux I__1361 (
            .O(N__15140),
            .I(\b2v_inst11.mult1_un75_sum_cry_2 ));
    CascadeMux I__1360 (
            .O(N__15137),
            .I(N__15134));
    InMux I__1359 (
            .O(N__15134),
            .I(N__15131));
    LocalMux I__1358 (
            .O(N__15131),
            .I(\b2v_inst11.mult1_un68_sum_cry_3_s ));
    InMux I__1357 (
            .O(N__15128),
            .I(\b2v_inst11.mult1_un75_sum_cry_3 ));
    InMux I__1356 (
            .O(N__15125),
            .I(N__15122));
    LocalMux I__1355 (
            .O(N__15122),
            .I(\b2v_inst11.mult1_un68_sum_cry_4_s ));
    InMux I__1354 (
            .O(N__15119),
            .I(\b2v_inst11.mult1_un75_sum_cry_4 ));
    CascadeMux I__1353 (
            .O(N__15116),
            .I(N__15113));
    InMux I__1352 (
            .O(N__15113),
            .I(N__15110));
    LocalMux I__1351 (
            .O(N__15110),
            .I(\b2v_inst11.mult1_un68_sum_cry_5_s ));
    InMux I__1350 (
            .O(N__15107),
            .I(\b2v_inst11.mult1_un75_sum_cry_5 ));
    InMux I__1349 (
            .O(N__15104),
            .I(N__15101));
    LocalMux I__1348 (
            .O(N__15101),
            .I(\b2v_inst11.mult1_un68_sum_cry_6_s ));
    CascadeMux I__1347 (
            .O(N__15098),
            .I(N__15094));
    CascadeMux I__1346 (
            .O(N__15097),
            .I(N__15090));
    InMux I__1345 (
            .O(N__15094),
            .I(N__15083));
    InMux I__1344 (
            .O(N__15093),
            .I(N__15083));
    InMux I__1343 (
            .O(N__15090),
            .I(N__15083));
    LocalMux I__1342 (
            .O(N__15083),
            .I(\b2v_inst11.mult1_un68_sum_i_0_8 ));
    InMux I__1341 (
            .O(N__15080),
            .I(\b2v_inst11.mult1_un75_sum_cry_6 ));
    CascadeMux I__1340 (
            .O(N__15077),
            .I(N__15074));
    InMux I__1339 (
            .O(N__15074),
            .I(N__15071));
    LocalMux I__1338 (
            .O(N__15071),
            .I(\b2v_inst11.mult1_un75_sum_axb_8 ));
    InMux I__1337 (
            .O(N__15068),
            .I(\b2v_inst11.mult1_un75_sum_cry_7 ));
    CascadeMux I__1336 (
            .O(N__15065),
            .I(\b2v_inst11.mult1_un75_sum_s_8_cascade_ ));
    InMux I__1335 (
            .O(N__15062),
            .I(\b2v_inst11.mult1_un68_sum_cry_2 ));
    InMux I__1334 (
            .O(N__15059),
            .I(\b2v_inst11.mult1_un68_sum_cry_3 ));
    InMux I__1333 (
            .O(N__15056),
            .I(\b2v_inst11.mult1_un68_sum_cry_4 ));
    InMux I__1332 (
            .O(N__15053),
            .I(\b2v_inst11.mult1_un68_sum_cry_5 ));
    InMux I__1331 (
            .O(N__15050),
            .I(\b2v_inst11.mult1_un68_sum_cry_6 ));
    InMux I__1330 (
            .O(N__15047),
            .I(\b2v_inst11.mult1_un68_sum_cry_7 ));
    CascadeMux I__1329 (
            .O(N__15044),
            .I(\b2v_inst11.mult1_un68_sum_s_8_cascade_ ));
    InMux I__1328 (
            .O(N__15041),
            .I(\b2v_inst200.un2_count_1_cry_9 ));
    InMux I__1327 (
            .O(N__15038),
            .I(\b2v_inst200.un2_count_1_cry_10 ));
    InMux I__1326 (
            .O(N__15035),
            .I(\b2v_inst200.un2_count_1_cry_11 ));
    InMux I__1325 (
            .O(N__15032),
            .I(\b2v_inst200.un2_count_1_cry_12 ));
    InMux I__1324 (
            .O(N__15029),
            .I(\b2v_inst200.un2_count_1_cry_13 ));
    InMux I__1323 (
            .O(N__15026),
            .I(\b2v_inst200.un2_count_1_cry_14 ));
    CascadeMux I__1322 (
            .O(N__15023),
            .I(N__15020));
    InMux I__1321 (
            .O(N__15020),
            .I(N__15017));
    LocalMux I__1320 (
            .O(N__15017),
            .I(N__15014));
    Odrv12 I__1319 (
            .O(N__15014),
            .I(\b2v_inst200.un2_count_1_axb_16 ));
    InMux I__1318 (
            .O(N__15011),
            .I(N__15002));
    InMux I__1317 (
            .O(N__15010),
            .I(N__15002));
    InMux I__1316 (
            .O(N__15009),
            .I(N__15002));
    LocalMux I__1315 (
            .O(N__15002),
            .I(N__14999));
    Odrv12 I__1314 (
            .O(N__14999),
            .I(\b2v_inst200.count_1_16 ));
    InMux I__1313 (
            .O(N__14996),
            .I(\b2v_inst200.un2_count_1_cry_15 ));
    InMux I__1312 (
            .O(N__14993),
            .I(bfn_1_8_0_));
    InMux I__1311 (
            .O(N__14990),
            .I(N__14986));
    InMux I__1310 (
            .O(N__14989),
            .I(N__14983));
    LocalMux I__1309 (
            .O(N__14986),
            .I(N__14980));
    LocalMux I__1308 (
            .O(N__14983),
            .I(\b2v_inst200.un2_count_1_axb_1 ));
    Odrv4 I__1307 (
            .O(N__14980),
            .I(\b2v_inst200.un2_count_1_axb_1 ));
    InMux I__1306 (
            .O(N__14975),
            .I(N__14971));
    InMux I__1305 (
            .O(N__14974),
            .I(N__14968));
    LocalMux I__1304 (
            .O(N__14971),
            .I(N__14965));
    LocalMux I__1303 (
            .O(N__14968),
            .I(\b2v_inst200.countZ0Z_2 ));
    Odrv4 I__1302 (
            .O(N__14965),
            .I(\b2v_inst200.countZ0Z_2 ));
    InMux I__1301 (
            .O(N__14960),
            .I(N__14956));
    InMux I__1300 (
            .O(N__14959),
            .I(N__14953));
    LocalMux I__1299 (
            .O(N__14956),
            .I(N__14950));
    LocalMux I__1298 (
            .O(N__14953),
            .I(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ));
    Odrv4 I__1297 (
            .O(N__14950),
            .I(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ));
    InMux I__1296 (
            .O(N__14945),
            .I(\b2v_inst200.un2_count_1_cry_1 ));
    InMux I__1295 (
            .O(N__14942),
            .I(\b2v_inst200.un2_count_1_cry_2 ));
    InMux I__1294 (
            .O(N__14939),
            .I(N__14935));
    InMux I__1293 (
            .O(N__14938),
            .I(N__14932));
    LocalMux I__1292 (
            .O(N__14935),
            .I(N__14929));
    LocalMux I__1291 (
            .O(N__14932),
            .I(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ));
    Odrv4 I__1290 (
            .O(N__14929),
            .I(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ));
    InMux I__1289 (
            .O(N__14924),
            .I(\b2v_inst200.un2_count_1_cry_3 ));
    InMux I__1288 (
            .O(N__14921),
            .I(\b2v_inst200.un2_count_1_cry_4 ));
    InMux I__1287 (
            .O(N__14918),
            .I(\b2v_inst200.un2_count_1_cry_5_cZ0 ));
    InMux I__1286 (
            .O(N__14915),
            .I(\b2v_inst200.un2_count_1_cry_6 ));
    InMux I__1285 (
            .O(N__14912),
            .I(\b2v_inst200.un2_count_1_cry_7 ));
    InMux I__1284 (
            .O(N__14909),
            .I(bfn_1_7_0_));
    CascadeMux I__1283 (
            .O(N__14906),
            .I(\b2v_inst200.count_RNIZ0Z_1_cascade_ ));
    CascadeMux I__1282 (
            .O(N__14903),
            .I(\b2v_inst200.un2_count_1_axb_1_cascade_ ));
    CascadeMux I__1281 (
            .O(N__14900),
            .I(N__14897));
    InMux I__1280 (
            .O(N__14897),
            .I(N__14893));
    InMux I__1279 (
            .O(N__14896),
            .I(N__14890));
    LocalMux I__1278 (
            .O(N__14893),
            .I(\b2v_inst200.count_3_1 ));
    LocalMux I__1277 (
            .O(N__14890),
            .I(\b2v_inst200.count_3_1 ));
    InMux I__1276 (
            .O(N__14885),
            .I(N__14882));
    LocalMux I__1275 (
            .O(N__14882),
            .I(N__14879));
    Odrv4 I__1274 (
            .O(N__14879),
            .I(\b2v_inst200.count_3_2 ));
    InMux I__1273 (
            .O(N__14876),
            .I(N__14873));
    LocalMux I__1272 (
            .O(N__14873),
            .I(N__14870));
    Odrv4 I__1271 (
            .O(N__14870),
            .I(\b2v_inst200.count_3_4 ));
    CascadeMux I__1270 (
            .O(N__14867),
            .I(\b2v_inst200.un25_clk_100khz_1_cascade_ ));
    CascadeMux I__1269 (
            .O(N__14864),
            .I(N__14861));
    InMux I__1268 (
            .O(N__14861),
            .I(N__14857));
    InMux I__1267 (
            .O(N__14860),
            .I(N__14854));
    LocalMux I__1266 (
            .O(N__14857),
            .I(\b2v_inst200.countZ0Z_16 ));
    LocalMux I__1265 (
            .O(N__14854),
            .I(\b2v_inst200.countZ0Z_16 ));
    InMux I__1264 (
            .O(N__14849),
            .I(N__14846));
    LocalMux I__1263 (
            .O(N__14846),
            .I(\b2v_inst200.un25_clk_100khz_0 ));
    InMux I__1262 (
            .O(N__14843),
            .I(N__14840));
    LocalMux I__1261 (
            .O(N__14840),
            .I(\b2v_inst200.count_RNIZ0Z_1 ));
    CascadeMux I__1260 (
            .O(N__14837),
            .I(\b2v_inst16.countZ0Z_1_cascade_ ));
    InMux I__1259 (
            .O(N__14834),
            .I(N__14831));
    LocalMux I__1258 (
            .O(N__14831),
            .I(\b2v_inst16.count_4_1 ));
    InMux I__1257 (
            .O(N__14828),
            .I(N__14825));
    LocalMux I__1256 (
            .O(N__14825),
            .I(\b2v_inst16.count_4_11 ));
    CascadeMux I__1255 (
            .O(N__14822),
            .I(\b2v_inst16.count_rst_0_cascade_ ));
    CascadeMux I__1254 (
            .O(N__14819),
            .I(\b2v_inst16.countZ0Z_11_cascade_ ));
    InMux I__1253 (
            .O(N__14816),
            .I(N__14813));
    LocalMux I__1252 (
            .O(N__14813),
            .I(\b2v_inst16.count_4_8 ));
    InMux I__1251 (
            .O(N__14810),
            .I(N__14807));
    LocalMux I__1250 (
            .O(N__14807),
            .I(\b2v_inst16.count_4_6 ));
    InMux I__1249 (
            .O(N__14804),
            .I(N__14801));
    LocalMux I__1248 (
            .O(N__14801),
            .I(\b2v_inst16.count_4_15 ));
    CascadeMux I__1247 (
            .O(N__14798),
            .I(\b2v_inst16.count_rst_12_cascade_ ));
    CascadeMux I__1246 (
            .O(N__14795),
            .I(\b2v_inst16.count_rst_13_cascade_ ));
    CascadeMux I__1245 (
            .O(N__14792),
            .I(\b2v_inst16.count_rst_14_cascade_ ));
    CascadeMux I__1244 (
            .O(N__14789),
            .I(\b2v_inst16.countZ0Z_9_cascade_ ));
    InMux I__1243 (
            .O(N__14786),
            .I(N__14783));
    LocalMux I__1242 (
            .O(N__14783),
            .I(\b2v_inst16.count_4_9 ));
    CascadeMux I__1241 (
            .O(N__14780),
            .I(\b2v_inst16.count_rst_6_cascade_ ));
    defparam IN_MUX_bfv_11_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_1_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(\b2v_inst6.un2_count_1_cry_8 ),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(\b2v_inst5.un2_count_1_cry_7 ),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(\b2v_inst36.un2_count_1_cry_7 ),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_8 ),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_16 ),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(b2v_inst20_un4_counter_7),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_8 ),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_16 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_24 ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(\b2v_inst16.un4_count_1_cry_8 ),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\b2v_inst11.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_94_cry_7 ),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\b2v_inst11.un1_count_cry_8 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\b2v_inst11.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    ICE_GB \b2v_inst200.count_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__17369),
            .GLOBALBUFFEROUTPUT(\b2v_inst200.count_en_g ));
    ICE_GB N_606_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__31250),
            .GLOBALBUFFEROUTPUT(N_606_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_1_0 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_1_0 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_1_0  (
            .in0(N__15679),
            .in1(N__17721),
            .in2(N__15710),
            .in3(N__17565),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_1_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_1_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst16.count_RNINJ2K1_7_LC_1_1_1  (
            .in0(N__15410),
            .in1(_gnd_net_),
            .in2(N__14798),
            .in3(N__20093),
            .lcout(\b2v_inst16.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_1_2 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_1_2 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_1_2  (
            .in0(N__15634),
            .in1(N__17722),
            .in2(N__15662),
            .in3(N__17566),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3  (
            .in0(_gnd_net_),
            .in1(N__14816),
            .in2(N__14795),
            .in3(N__20094),
            .lcout(\b2v_inst16.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_1_4 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_1_4 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_1_4  (
            .in0(N__15612),
            .in1(N__17723),
            .in2(N__15593),
            .in3(N__17567),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_1_1_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_1_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNIRP4K1_9_LC_1_1_5  (
            .in0(_gnd_net_),
            .in1(N__14786),
            .in2(N__14792),
            .in3(N__20095),
            .lcout(\b2v_inst16.countZ0Z_9 ),
            .ltout(\b2v_inst16.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_9_LC_1_1_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_9_LC_1_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_9_LC_1_1_6 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst16.count_9_LC_1_1_6  (
            .in0(N__17729),
            .in1(N__17568),
            .in2(N__14789),
            .in3(N__15592),
            .lcout(\b2v_inst16.count_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36421),
            .ce(N__20108),
            .sr(N__17888));
    defparam \b2v_inst16.count_11_LC_1_2_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_11_LC_1_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_11_LC_1_2_0 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst16.count_11_LC_1_2_0  (
            .in0(N__17542),
            .in1(N__15893),
            .in2(N__17731),
            .in3(N__15909),
            .lcout(\b2v_inst16.count_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36469),
            .ce(N__20096),
            .sr(N__17906));
    defparam \b2v_inst16.count_RNI_1_LC_1_2_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_1_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_1_LC_1_2_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst16.count_RNI_1_LC_1_2_1  (
            .in0(N__15478),
            .in1(N__17700),
            .in2(_gnd_net_),
            .in3(N__15499),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI2J651_1_LC_1_2_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI2J651_1_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI2J651_1_LC_1_2_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNI2J651_1_LC_1_2_2  (
            .in0(_gnd_net_),
            .in1(N__14834),
            .in2(N__14780),
            .in3(N__20085),
            .lcout(\b2v_inst16.countZ0Z_1 ),
            .ltout(\b2v_inst16.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_1_LC_1_2_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_1_LC_1_2_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_1_LC_1_2_3 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \b2v_inst16.count_1_LC_1_2_3  (
            .in0(_gnd_net_),
            .in1(N__17704),
            .in2(N__14837),
            .in3(N__15500),
            .lcout(\b2v_inst16.count_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36469),
            .ce(N__20096),
            .sr(N__17906));
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_2_4 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_2_4 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_2_4  (
            .in0(N__17541),
            .in1(N__15892),
            .in2(N__17730),
            .in3(N__15910),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIDGU31_11_LC_1_2_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIDGU31_11_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIDGU31_11_LC_1_2_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \b2v_inst16.count_RNIDGU31_11_LC_1_2_5  (
            .in0(N__20086),
            .in1(N__14828),
            .in2(N__14822),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.countZ0Z_11 ),
            .ltout(\b2v_inst16.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_11_LC_1_2_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_11_LC_1_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_11_LC_1_2_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst16.count_RNI_11_LC_1_2_6  (
            .in0(N__15657),
            .in1(N__15614),
            .in2(N__14819),
            .in3(N__15477),
            .lcout(\b2v_inst16.count_4_i_a3_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_8_LC_1_2_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_8_LC_1_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_8_LC_1_2_7 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst16.count_8_LC_1_2_7  (
            .in0(N__17543),
            .in1(N__15656),
            .in2(N__15635),
            .in3(N__17708),
            .lcout(\b2v_inst16.count_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36469),
            .ce(N__20096),
            .sr(N__17906));
    defparam \b2v_inst16.count_RNILG1K1_6_LC_1_3_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILG1K1_6_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILG1K1_6_LC_1_3_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNILG1K1_6_LC_1_3_0  (
            .in0(N__20089),
            .in1(N__14810),
            .in2(_gnd_net_),
            .in3(N__15721),
            .lcout(\b2v_inst16.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_6_LC_1_3_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_6_LC_1_3_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_6_LC_1_3_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_6_LC_1_3_1  (
            .in0(N__15722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36422),
            .ce(N__20104),
            .sr(N__17903));
    defparam \b2v_inst16.count_RNILS241_15_LC_1_3_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILS241_15_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILS241_15_LC_1_3_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst16.count_RNILS241_15_LC_1_3_2  (
            .in0(N__20105),
            .in1(N__15851),
            .in2(_gnd_net_),
            .in3(N__14804),
            .lcout(\b2v_inst16.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_15_LC_1_3_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_15_LC_1_3_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_15_LC_1_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_15_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15850),
            .lcout(\b2v_inst16.count_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36422),
            .ce(N__20104),
            .sr(N__17903));
    defparam \b2v_inst16.count_RNI_0_0_LC_1_3_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_0_0_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_0_0_LC_1_3_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst16.count_RNI_0_0_LC_1_3_4  (
            .in0(N__15502),
            .in1(N__17699),
            .in2(_gnd_net_),
            .in3(N__15538),
            .lcout(\b2v_inst16.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_0_LC_1_3_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_0_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_0_LC_1_3_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst16.count_RNI_0_LC_1_3_5  (
            .in0(_gnd_net_),
            .in1(N__15537),
            .in2(_gnd_net_),
            .in3(N__15503),
            .lcout(\b2v_inst16.N_416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI1QV41_2_LC_1_3_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_1_3_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNI1QV41_2_LC_1_3_6  (
            .in0(N__14885),
            .in1(N__16564),
            .in2(_gnd_net_),
            .in3(N__14960),
            .lcout(\b2v_inst200.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50251_4_LC_1_3_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50251_4_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50251_4_LC_1_3_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNI50251_4_LC_1_3_7  (
            .in0(N__16565),
            .in1(N__14876),
            .in2(_gnd_net_),
            .in3(N__14939),
            .lcout(\b2v_inst200.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9S71_16_LC_1_4_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_1_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNIB9S71_16_LC_1_4_0  (
            .in0(N__15009),
            .in1(N__14860),
            .in2(_gnd_net_),
            .in3(N__16561),
            .lcout(\b2v_inst200.un2_count_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_16_LC_1_4_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_16_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_16_LC_1_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_16_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15011),
            .lcout(\b2v_inst200.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36401),
            .ce(N__16485),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNID13N_0_1_LC_1_4_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNID13N_0_1_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNID13N_0_1_LC_1_4_2 .LUT_INIT=16'b0000000001000111;
    LogicCell40 \b2v_inst200.count_RNID13N_0_1_LC_1_4_2  (
            .in0(N__14843),
            .in1(N__16563),
            .in2(N__14900),
            .in3(N__14974),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIOAVU1_1_LC_1_4_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIOAVU1_1_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIOAVU1_1_LC_1_4_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst200.count_RNIOAVU1_1_LC_1_4_3  (
            .in0(N__14849),
            .in1(N__16334),
            .in2(N__14867),
            .in3(N__16105),
            .lcout(\b2v_inst200.un25_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9S71_0_16_LC_1_4_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9S71_0_16_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9S71_0_16_LC_1_4_4 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \b2v_inst200.count_RNIB9S71_0_16_LC_1_4_4  (
            .in0(N__15010),
            .in1(N__15976),
            .in2(N__14864),
            .in3(N__16562),
            .lcout(\b2v_inst200.un25_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_1_LC_1_4_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_1_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_1_LC_1_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst200.count_RNI_1_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(N__16104),
            .in2(_gnd_net_),
            .in3(N__14989),
            .lcout(\b2v_inst200.count_RNIZ0Z_1 ),
            .ltout(\b2v_inst200.count_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNID13N_1_LC_1_4_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNID13N_1_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNID13N_1_LC_1_4_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst200.count_RNID13N_1_LC_1_4_6  (
            .in0(_gnd_net_),
            .in1(N__14896),
            .in2(N__14906),
            .in3(N__16560),
            .lcout(\b2v_inst200.un2_count_1_axb_1 ),
            .ltout(\b2v_inst200.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_1_LC_1_4_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_1_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_1_LC_1_4_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst200.count_1_LC_1_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14903),
            .in3(N__16106),
            .lcout(\b2v_inst200.count_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36401),
            .ce(N__16485),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_11_LC_1_5_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_11_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_11_LC_1_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_11_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16349),
            .lcout(\b2v_inst200.count_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36490),
            .ce(N__16488),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_14_LC_1_5_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_14_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_14_LC_1_5_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst200.count_14_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(N__15833),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36490),
            .ce(N__16488),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_2_LC_1_5_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_2_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_2_LC_1_5_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst200.count_2_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(N__14959),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36490),
            .ce(N__16488),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_4_LC_1_5_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_4_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_4_LC_1_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_4_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14938),
            .lcout(\b2v_inst200.count_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36490),
            .ce(N__16488),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_6_LC_1_5_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_6_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_6_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_6_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16040),
            .lcout(\b2v_inst200.count_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36490),
            .ce(N__16488),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_7_LC_1_5_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_7_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_7_LC_1_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_7_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16022),
            .lcout(\b2v_inst200.count_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36490),
            .ce(N__16488),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_10_LC_1_5_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_10_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_10_LC_1_5_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_10_LC_1_5_6  (
            .in0(N__15964),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36490),
            .ce(N__16488),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_1_c_LC_1_6_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_1_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_1_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_1_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__14990),
            .in2(N__16114),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_1_6_1 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_1_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__14975),
            .in2(_gnd_net_),
            .in3(N__14945),
            .lcout(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_1 ),
            .carryout(\b2v_inst200.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_1_6_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_1_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__16316),
            .in2(_gnd_net_),
            .in3(N__14942),
            .lcout(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_2 ),
            .carryout(\b2v_inst200.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_1_6_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_1_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__16255),
            .in2(_gnd_net_),
            .in3(N__14924),
            .lcout(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_3 ),
            .carryout(\b2v_inst200.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_1_6_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_1_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__16364),
            .in2(_gnd_net_),
            .in3(N__14921),
            .lcout(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_4 ),
            .carryout(\b2v_inst200.un2_count_1_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_1_6_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_1_6_5 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_1_6_5  (
            .in0(N__19437),
            .in1(_gnd_net_),
            .in2(N__16156),
            .in3(N__14918),
            .lcout(\b2v_inst200.count_1_6 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_5_cZ0 ),
            .carryout(\b2v_inst200.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_1_6_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_1_6_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16591),
            .in3(N__14915),
            .lcout(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_6 ),
            .carryout(\b2v_inst200.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_1_6_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_1_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_1_6_7  (
            .in0(N__19438),
            .in1(N__16193),
            .in2(_gnd_net_),
            .in3(N__14912),
            .lcout(\b2v_inst200.count_1_8 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_7 ),
            .carryout(\b2v_inst200.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_1_7_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_1_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__16073),
            .in2(_gnd_net_),
            .in3(N__14909),
            .lcout(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_1_7_1 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_1_7_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_1_7_1  (
            .in0(N__19439),
            .in1(_gnd_net_),
            .in2(N__15929),
            .in3(N__15041),
            .lcout(\b2v_inst200.count_1_10 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_9 ),
            .carryout(\b2v_inst200.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_1_7_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_1_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_1_7_2  (
            .in0(N__19441),
            .in1(N__16327),
            .in2(_gnd_net_),
            .in3(N__15038),
            .lcout(\b2v_inst200.count_1_11 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_10 ),
            .carryout(\b2v_inst200.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_1_7_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_1_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__16052),
            .in2(_gnd_net_),
            .in3(N__15035),
            .lcout(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_11 ),
            .carryout(\b2v_inst200.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_1_7_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_1_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__16634),
            .in2(_gnd_net_),
            .in3(N__15032),
            .lcout(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_12 ),
            .carryout(\b2v_inst200.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_1_7_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_1_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__16303),
            .in2(_gnd_net_),
            .in3(N__15029),
            .lcout(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_13 ),
            .carryout(\b2v_inst200.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_1_7_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_1_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__16187),
            .in2(_gnd_net_),
            .in3(N__15026),
            .lcout(\b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_14 ),
            .carryout(\b2v_inst200.un2_count_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_1_7_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_1_7_7 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_1_7_7  (
            .in0(N__19440),
            .in1(_gnd_net_),
            .in2(N__15023),
            .in3(N__14996),
            .lcout(\b2v_inst200.count_1_16 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_15 ),
            .carryout(\b2v_inst200.un2_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_1_8_0 .C_ON=1'b0;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_1_8_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_1_8_0  (
            .in0(N__15980),
            .in1(N__19446),
            .in2(_gnd_net_),
            .in3(N__14993),
            .lcout(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_17_LC_1_8_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_17_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_17_LC_1_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_17_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15994),
            .lcout(\b2v_inst200.count_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36542),
            .ce(N__16490),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_0_LC_1_8_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_0_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_0_LC_1_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst200.count_RNI_0_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__16115),
            .in2(_gnd_net_),
            .in3(N__19445),
            .lcout(\b2v_inst200.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21314),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_1_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_1_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__18131),
            .in2(N__16738),
            .in3(N__15062),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_1_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_1_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__16734),
            .in2(N__16430),
            .in3(N__15059),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_1_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_1_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__16418),
            .in2(N__18157),
            .in3(N__15056),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_1_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_1_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__18153),
            .in2(N__16409),
            .in3(N__15053),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_1_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_1_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_1_9_5  (
            .in0(N__18500),
            .in1(N__16397),
            .in2(N__16739),
            .in3(N__15050),
            .lcout(\b2v_inst11.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_1_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_1_9_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16757),
            .in3(N__15047),
            .lcout(\b2v_inst11.mult1_un68_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un68_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_1_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_1_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15044),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__21346),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_1_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__16826),
            .in2(N__15097),
            .in3(N__15140),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_1_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__15093),
            .in2(N__15137),
            .in3(N__15128),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_1_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__15125),
            .in2(N__18508),
            .in3(N__15119),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_1_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(N__15116),
            .in3(N__15107),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_1_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_1_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_1_10_5  (
            .in0(N__16844),
            .in1(N__15104),
            .in2(N__15098),
            .in3(N__15080),
            .lcout(\b2v_inst11.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_1_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_1_10_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15077),
            .in3(N__15068),
            .lcout(\b2v_inst11.mult1_un75_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_1_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_1_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15065),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__21419),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_11_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__16820),
            .in2(N__16801),
            .in3(N__15164),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_11_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__16797),
            .in2(N__16721),
            .in3(N__15161),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_11_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__16700),
            .in2(N__16784),
            .in3(N__15158),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_11_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__16783),
            .in2(N__16685),
            .in3(N__15155),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_11_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_11_5  (
            .in0(N__16934),
            .in1(N__16664),
            .in2(N__16802),
            .in3(N__15152),
            .lcout(\b2v_inst11.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16892),
            .in3(N__15149),
            .lcout(\b2v_inst11.mult1_un89_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un89_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15146),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__21455),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__16814),
            .in2(N__15205),
            .in3(N__15143),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__15201),
            .in2(N__15245),
            .in3(N__15236),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__15233),
            .in2(N__16940),
            .in3(N__15227),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__16938),
            .in2(N__15224),
            .in3(N__15215),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_12_5  (
            .in0(N__17009),
            .in1(N__15212),
            .in2(N__15206),
            .in3(N__15188),
            .lcout(\b2v_inst11.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15185),
            .in3(N__15176),
            .lcout(\b2v_inst11.mult1_un96_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un96_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15173),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI0AHN_8_LC_1_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_1_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNI0AHN_8_LC_1_13_0  (
            .in0(N__30732),
            .in1(N__15170),
            .in2(_gnd_net_),
            .in3(N__15397),
            .lcout(\b2v_inst11.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_8_LC_1_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_8_LC_1_13_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_8_LC_1_13_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_8_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15401),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36580),
            .ce(N__32182),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI2DIN_9_LC_1_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_1_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNI2DIN_9_LC_1_13_2  (
            .in0(N__30731),
            .in1(N__15275),
            .in2(_gnd_net_),
            .in3(N__15379),
            .lcout(\b2v_inst11.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_9_LC_1_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_9_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_9_LC_1_13_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_9_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15383),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36580),
            .ce(N__32182),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIB49T_10_LC_1_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIB49T_10_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIB49T_10_LC_1_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_RNIB49T_10_LC_1_13_4  (
            .in0(N__15365),
            .in1(N__15269),
            .in2(_gnd_net_),
            .in3(N__30733),
            .lcout(\b2v_inst11.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_10_LC_1_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_10_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_10_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_10_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15364),
            .lcout(\b2v_inst11.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36580),
            .ce(N__32182),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIK61M_11_LC_1_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIK61M_11_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIK61M_11_LC_1_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_RNIK61M_11_LC_1_13_6  (
            .in0(N__15350),
            .in1(N__15263),
            .in2(_gnd_net_),
            .in3(N__30734),
            .lcout(\b2v_inst11.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_11_LC_1_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_11_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_11_LC_1_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_11_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15349),
            .lcout(\b2v_inst11.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36580),
            .ce(N__32182),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_1_LC_1_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_1_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_1_LC_1_14_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \b2v_inst11.count_RNI_1_LC_1_14_0  (
            .in0(N__18432),
            .in1(N__18471),
            .in2(_gnd_net_),
            .in3(N__17109),
            .lcout(),
            .ltout(\b2v_inst11.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI14G9_1_LC_1_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI14G9_1_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI14G9_1_LC_1_14_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst11.count_RNI14G9_1_LC_1_14_1  (
            .in0(N__30729),
            .in1(_gnd_net_),
            .in2(N__15257),
            .in3(N__15251),
            .lcout(\b2v_inst11.countZ0Z_1 ),
            .ltout(\b2v_inst11.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_1_LC_1_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_1_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_1_LC_1_14_2 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \b2v_inst11.count_1_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__18473),
            .in2(N__15254),
            .in3(N__17113),
            .lcout(\b2v_inst11.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__32181),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_0_LC_1_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_0_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_0_LC_1_14_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst11.count_0_LC_1_14_3  (
            .in0(N__18472),
            .in1(_gnd_net_),
            .in2(N__17142),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__32181),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIKNAN_2_LC_1_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_1_14_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_RNIKNAN_2_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__15314),
            .in2(N__15302),
            .in3(N__30728),
            .lcout(\b2v_inst11.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_2_LC_1_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_2_LC_1_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_2_LC_1_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_2_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15301),
            .lcout(\b2v_inst11.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__32181),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIM92M_12_LC_1_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIM92M_12_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIM92M_12_LC_1_14_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_RNIM92M_12_LC_1_14_6  (
            .in0(N__15335),
            .in1(N__15308),
            .in2(_gnd_net_),
            .in3(N__30730),
            .lcout(\b2v_inst11.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_12_LC_1_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_12_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_12_LC_1_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_12_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15334),
            .lcout(\b2v_inst11.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__32181),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_LC_1_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_1_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__18478),
            .in2(N__18433),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\b2v_inst11.un1_count_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_15_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_15_1  (
            .in0(N__17146),
            .in1(_gnd_net_),
            .in2(N__18394),
            .in3(N__15290),
            .lcout(\b2v_inst11.count_1_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_1_cZ0 ),
            .carryout(\b2v_inst11.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_15_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_15_2  (
            .in0(N__17139),
            .in1(N__18354),
            .in2(_gnd_net_),
            .in3(N__15287),
            .lcout(\b2v_inst11.count_1_3 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_2 ),
            .carryout(\b2v_inst11.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_15_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_15_3  (
            .in0(N__17143),
            .in1(N__18319),
            .in2(_gnd_net_),
            .in3(N__15284),
            .lcout(\b2v_inst11.count_1_4 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_3 ),
            .carryout(\b2v_inst11.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_15_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_15_4  (
            .in0(N__17140),
            .in1(N__18286),
            .in2(_gnd_net_),
            .in3(N__15281),
            .lcout(\b2v_inst11.count_1_5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_4 ),
            .carryout(\b2v_inst11.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_15_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_15_5  (
            .in0(N__17144),
            .in1(N__18847),
            .in2(_gnd_net_),
            .in3(N__15278),
            .lcout(\b2v_inst11.count_1_6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_5 ),
            .carryout(\b2v_inst11.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_15_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_15_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_15_6  (
            .in0(N__17141),
            .in1(N__18814),
            .in2(_gnd_net_),
            .in3(N__15404),
            .lcout(\b2v_inst11.count_1_7 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_6 ),
            .carryout(\b2v_inst11.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_15_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_15_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_15_7  (
            .in0(N__17145),
            .in1(N__18787),
            .in2(_gnd_net_),
            .in3(N__15386),
            .lcout(\b2v_inst11.count_1_8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_7 ),
            .carryout(\b2v_inst11.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_16_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_16_0  (
            .in0(N__17147),
            .in1(N__18748),
            .in2(_gnd_net_),
            .in3(N__15368),
            .lcout(\b2v_inst11.count_1_9 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\b2v_inst11.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_16_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_16_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_16_1  (
            .in0(N__17152),
            .in1(N__18699),
            .in2(_gnd_net_),
            .in3(N__15353),
            .lcout(\b2v_inst11.count_1_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_9 ),
            .carryout(\b2v_inst11.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_16_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_16_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_16_2  (
            .in0(N__17148),
            .in1(N__18651),
            .in2(_gnd_net_),
            .in3(N__15338),
            .lcout(\b2v_inst11.count_1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_10 ),
            .carryout(\b2v_inst11.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_16_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_16_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_16_3  (
            .in0(N__17151),
            .in1(N__18615),
            .in2(_gnd_net_),
            .in3(N__15323),
            .lcout(\b2v_inst11.count_1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_11 ),
            .carryout(\b2v_inst11.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_16_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_16_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_16_4  (
            .in0(N__17149),
            .in1(N__18556),
            .in2(_gnd_net_),
            .in3(N__15320),
            .lcout(\b2v_inst11.count_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_12 ),
            .carryout(\b2v_inst11.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_16_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_16_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_16_5  (
            .in0(N__17153),
            .in1(N__18970),
            .in2(_gnd_net_),
            .in3(N__15317),
            .lcout(\b2v_inst11.count_1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_13 ),
            .carryout(\b2v_inst11.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_16_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_16_6  (
            .in0(N__17150),
            .in1(N__18934),
            .in2(_gnd_net_),
            .in3(N__15437),
            .lcout(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_1_0 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_1_0 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_1_0  (
            .in0(N__17571),
            .in1(N__15784),
            .in2(N__15812),
            .in3(N__17713),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_2_1_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_2_1_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNIHAVJ1_4_LC_2_1_1  (
            .in0(_gnd_net_),
            .in1(N__15428),
            .in2(N__15434),
            .in3(N__20087),
            .lcout(\b2v_inst16.countZ0Z_4 ),
            .ltout(\b2v_inst16.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_4_LC_2_1_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_4_LC_2_1_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_4_LC_2_1_2 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.count_4_LC_2_1_2  (
            .in0(N__17575),
            .in1(N__17716),
            .in2(N__15431),
            .in3(N__15785),
            .lcout(\b2v_inst16.count_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36420),
            .ce(N__20106),
            .sr(N__17899));
    defparam \b2v_inst16.count_3_LC_2_1_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_3_LC_2_1_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_3_LC_2_1_3 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst16.count_3_LC_2_1_3  (
            .in0(N__17715),
            .in1(N__17577),
            .in2(N__17489),
            .in3(N__17822),
            .lcout(\b2v_inst16.count_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36420),
            .ce(N__20106),
            .sr(N__17899));
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4  (
            .in0(N__15768),
            .in1(N__17714),
            .in2(N__17579),
            .in3(N__15748),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5  (
            .in0(_gnd_net_),
            .in1(N__15416),
            .in2(N__15422),
            .in3(N__20088),
            .lcout(\b2v_inst16.countZ0Z_5 ),
            .ltout(\b2v_inst16.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_5_LC_2_1_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_5_LC_2_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_5_LC_2_1_6 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.count_5_LC_2_1_6  (
            .in0(N__17576),
            .in1(N__17717),
            .in2(N__15419),
            .in3(N__15749),
            .lcout(\b2v_inst16.count_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36420),
            .ce(N__20106),
            .sr(N__17899));
    defparam \b2v_inst16.count_7_LC_2_1_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_7_LC_2_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_7_LC_2_1_7 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst16.count_7_LC_2_1_7  (
            .in0(N__17578),
            .in1(N__15704),
            .in2(N__17732),
            .in3(N__15680),
            .lcout(\b2v_inst16.count_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36420),
            .ce(N__20106),
            .sr(N__17899));
    defparam \b2v_inst16.count_2_LC_2_2_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_2_LC_2_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_2_LC_2_2_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \b2v_inst16.count_2_LC_2_2_0  (
            .in0(N__17711),
            .in1(N__15447),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36468),
            .ce(N__20038),
            .sr(N__17904));
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_2_2_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_2_2_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst16.count_RNID4TJ1_2_LC_2_2_1  (
            .in0(N__15451),
            .in1(N__17712),
            .in2(N__15515),
            .in3(N__20039),
            .lcout(),
            .ltout(\b2v_inst16.countZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNID4TJ1_2_2_LC_2_2_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNID4TJ1_2_2_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNID4TJ1_2_2_LC_2_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst16.count_RNID4TJ1_2_2_LC_2_2_2  (
            .in0(N__19958),
            .in1(N__15865),
            .in2(N__15566),
            .in3(N__15734),
            .lcout(),
            .ltout(\b2v_inst16.count_4_i_a3_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI2T6K2_13_LC_2_2_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI2T6K2_13_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI2T6K2_13_LC_2_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst16.count_RNI2T6K2_13_LC_2_2_3  (
            .in0(N__15554),
            .in1(N__15563),
            .in2(N__15557),
            .in3(N__17465),
            .lcout(\b2v_inst16.N_414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_4_LC_2_2_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_4_LC_2_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_4_LC_2_2_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst16.count_RNI_4_LC_2_2_4  (
            .in0(N__15769),
            .in1(N__15808),
            .in2(_gnd_net_),
            .in3(N__15708),
            .lcout(\b2v_inst16.count_4_i_a3_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_2_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNI1I651_0_LC_2_2_5  (
            .in0(N__15548),
            .in1(N__15521),
            .in2(_gnd_net_),
            .in3(N__20036),
            .lcout(\b2v_inst16.countZ0Z_0 ),
            .ltout(\b2v_inst16.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_0_LC_2_2_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_0_LC_2_2_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_0_LC_2_2_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \b2v_inst16.count_0_LC_2_2_6  (
            .in0(N__17710),
            .in1(_gnd_net_),
            .in2(N__15542),
            .in3(N__15539),
            .lcout(\b2v_inst16.count_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36468),
            .ce(N__20038),
            .sr(N__17904));
    defparam \b2v_inst16.count_RNID4TJ1_0_2_LC_2_2_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNID4TJ1_0_2_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNID4TJ1_0_2_LC_2_2_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \b2v_inst16.count_RNID4TJ1_0_2_LC_2_2_7  (
            .in0(N__15511),
            .in1(N__17709),
            .in2(N__15452),
            .in3(N__20037),
            .lcout(\b2v_inst16.un4_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_2_3_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_2_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_LC_2_3_0  (
            .in0(_gnd_net_),
            .in1(N__15501),
            .in2(N__15479),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_3_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_3_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15461),
            .in3(N__15818),
            .lcout(\b2v_inst16.un4_count_1_cry_1_c_RNIAGMEZ0 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_1 ),
            .carryout(\b2v_inst16.un4_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_3_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_3_2  (
            .in0(_gnd_net_),
            .in1(N__17821),
            .in2(_gnd_net_),
            .in3(N__15815),
            .lcout(\b2v_inst16.un4_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_2 ),
            .carryout(\b2v_inst16.un4_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_3_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_3_3  (
            .in0(_gnd_net_),
            .in1(N__15807),
            .in2(_gnd_net_),
            .in3(N__15773),
            .lcout(\b2v_inst16.un4_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_3 ),
            .carryout(\b2v_inst16.un4_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_3_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_3_4  (
            .in0(_gnd_net_),
            .in1(N__15770),
            .in2(_gnd_net_),
            .in3(N__15737),
            .lcout(\b2v_inst16.un4_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_4 ),
            .carryout(\b2v_inst16.un4_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_3_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_3_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_3_5  (
            .in0(N__17682),
            .in1(N__15733),
            .in2(_gnd_net_),
            .in3(N__15713),
            .lcout(\b2v_inst16.count_rst_11 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_5 ),
            .carryout(\b2v_inst16.un4_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_3_6 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_3_6  (
            .in0(_gnd_net_),
            .in1(N__15709),
            .in2(_gnd_net_),
            .in3(N__15665),
            .lcout(\b2v_inst16.un4_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_6 ),
            .carryout(\b2v_inst16.un4_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_3_7 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_3_7  (
            .in0(_gnd_net_),
            .in1(N__15661),
            .in2(_gnd_net_),
            .in3(N__15617),
            .lcout(\b2v_inst16.un4_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_7 ),
            .carryout(\b2v_inst16.un4_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_4_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(N__15613),
            .in2(_gnd_net_),
            .in3(N__15572),
            .lcout(\b2v_inst16.un4_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_4_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_4_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_4_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_4_1  (
            .in0(N__17727),
            .in1(N__19954),
            .in2(_gnd_net_),
            .in3(N__15569),
            .lcout(\b2v_inst16.count_rst ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_9 ),
            .carryout(\b2v_inst16.un4_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_4_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(N__15911),
            .in2(_gnd_net_),
            .in3(N__15881),
            .lcout(\b2v_inst16.un4_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_10 ),
            .carryout(\b2v_inst16.un4_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_4_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_4_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_4_3  (
            .in0(N__17724),
            .in1(N__17420),
            .in2(_gnd_net_),
            .in3(N__15878),
            .lcout(\b2v_inst16.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_11 ),
            .carryout(\b2v_inst16.un4_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNIHM041_LC_2_4_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNIHM041_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNIHM041_LC_2_4_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_12_c_RNIHM041_LC_2_4_4  (
            .in0(N__17728),
            .in1(N__17941),
            .in2(_gnd_net_),
            .in3(N__15875),
            .lcout(\b2v_inst16.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_12 ),
            .carryout(\b2v_inst16.un4_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_4_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_4_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_4_5  (
            .in0(N__17725),
            .in1(N__17453),
            .in2(_gnd_net_),
            .in3(N__15872),
            .lcout(\b2v_inst16.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_13 ),
            .carryout(\b2v_inst16.un4_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_4_6 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_4_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_4_6  (
            .in0(N__15869),
            .in1(N__17726),
            .in2(_gnd_net_),
            .in3(N__15854),
            .lcout(\b2v_inst16.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_10_LC_2_4_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_10_LC_2_4_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_10_LC_2_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_10_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20134),
            .lcout(\b2v_inst16.count_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36619),
            .ce(N__20103),
            .sr(N__17905));
    defparam \b2v_inst16.curr_state_1_LC_2_5_0 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_1_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_1_LC_2_5_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \b2v_inst16.curr_state_1_LC_2_5_0  (
            .in0(N__27735),
            .in1(N__17564),
            .in2(_gnd_net_),
            .in3(N__27770),
            .lcout(\b2v_inst16.curr_state_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36438),
            .ce(N__32177),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_0_LC_2_5_1 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_0_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_0_LC_2_5_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst16.curr_state_0_LC_2_5_1  (
            .in0(N__33576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27736),
            .lcout(\b2v_inst16.curr_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36438),
            .ce(N__32177),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73Q71_14_LC_2_5_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_2_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNI73Q71_14_LC_2_5_2  (
            .in0(N__16558),
            .in1(N__15839),
            .in2(_gnd_net_),
            .in3(N__15832),
            .lcout(\b2v_inst200.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI96451_6_LC_2_5_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI96451_6_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI96451_6_LC_2_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI96451_6_LC_2_5_3  (
            .in0(N__16046),
            .in1(N__16039),
            .in2(_gnd_net_),
            .in3(N__16555),
            .lcout(\b2v_inst200.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9551_7_LC_2_5_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9551_7_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9551_7_LC_2_5_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNIB9551_7_LC_2_5_4  (
            .in0(N__16556),
            .in1(N__16028),
            .in2(_gnd_net_),
            .in3(N__16021),
            .lcout(\b2v_inst200.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDCT71_17_LC_2_5_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_2_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIDCT71_17_LC_2_5_5  (
            .in0(N__16010),
            .in1(N__15998),
            .in2(_gnd_net_),
            .in3(N__16559),
            .lcout(\b2v_inst200.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_2_5_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_2_5_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst200.count_RNIOMPC1_10_LC_2_5_6  (
            .in0(N__16557),
            .in1(_gnd_net_),
            .in2(N__15965),
            .in3(N__15947),
            .lcout(\b2v_inst200.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_0_LC_2_5_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_0_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_0_LC_2_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNIC03N_0_LC_2_5_7  (
            .in0(N__16079),
            .in1(N__16554),
            .in2(_gnd_net_),
            .in3(N__15938),
            .lcout(\b2v_inst200.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_8_LC_2_6_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_8_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_8_LC_2_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_8_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16217),
            .lcout(\b2v_inst200.count_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36470),
            .ce(N__16486),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_15_LC_2_6_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_15_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_15_LC_2_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_15_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16171),
            .lcout(\b2v_inst200.count_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36470),
            .ce(N__16486),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDC651_0_8_LC_2_6_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDC651_0_8_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDC651_0_8_LC_2_6_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \b2v_inst200.count_RNIDC651_0_8_LC_2_6_2  (
            .in0(N__16573),
            .in1(N__15925),
            .in2(N__16205),
            .in3(N__16216),
            .lcout(\b2v_inst200.un25_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDC651_8_LC_2_6_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDC651_8_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDC651_8_LC_2_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNIDC651_8_LC_2_6_3  (
            .in0(N__16215),
            .in1(N__16201),
            .in2(_gnd_net_),
            .in3(N__16571),
            .lcout(\b2v_inst200.un2_count_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI2KKU_15_LC_2_6_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI2KKU_15_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI2KKU_15_LC_2_6_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst200.count_RNI2KKU_15_LC_2_6_4  (
            .in0(N__16572),
            .in1(_gnd_net_),
            .in2(N__16172),
            .in3(N__16180),
            .lcout(\b2v_inst200.un2_count_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI2KKU_0_15_LC_2_6_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI2KKU_0_15_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI2KKU_0_15_LC_2_6_5 .LUT_INIT=16'b0011000001010000;
    LogicCell40 \b2v_inst200.count_RNI2KKU_0_15_LC_2_6_5  (
            .in0(N__16181),
            .in1(N__16170),
            .in2(N__16157),
            .in3(N__16574),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI5RUP8_8_LC_2_6_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI5RUP8_8_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI5RUP8_8_LC_2_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNI5RUP8_8_LC_2_6_6  (
            .in0(N__16139),
            .in1(N__16133),
            .in2(N__16121),
            .in3(N__16280),
            .lcout(\b2v_inst200.count_RNI5RUP8Z0Z_8 ),
            .ltout(\b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_0_LC_2_6_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_0_LC_2_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_0_LC_2_6_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst200.count_0_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16118),
            .in3(N__16110),
            .lcout(\b2v_inst200.count_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36470),
            .ce(N__16486),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_12_LC_2_7_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_12_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_12_LC_2_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_12_LC_2_7_0  (
            .in0(N__16061),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36491),
            .ce(N__16487),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_9_LC_2_7_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_9_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_9_LC_2_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_9_LC_2_7_1  (
            .in0(N__16375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36491),
            .ce(N__16487),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIFF751_9_LC_2_7_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIFF751_9_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIFF751_9_LC_2_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNIFF751_9_LC_2_7_2  (
            .in0(N__16567),
            .in1(N__16387),
            .in2(_gnd_net_),
            .in3(N__16374),
            .lcout(\b2v_inst200.un2_count_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3TN71_12_LC_2_7_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_2_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI3TN71_12_LC_2_7_3  (
            .in0(N__16067),
            .in1(N__16060),
            .in2(_gnd_net_),
            .in3(N__16569),
            .lcout(\b2v_inst200.countZ0Z_12 ),
            .ltout(\b2v_inst200.countZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIFF751_0_9_LC_2_7_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIFF751_0_9_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIFF751_0_9_LC_2_7_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \b2v_inst200.count_RNIFF751_0_9_LC_2_7_4  (
            .in0(N__16570),
            .in1(N__16388),
            .in2(N__16379),
            .in3(N__16376),
            .lcout(\b2v_inst200.un25_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73351_5_LC_2_7_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73351_5_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73351_5_LC_2_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNI73351_5_LC_2_7_5  (
            .in0(N__16607),
            .in1(N__16566),
            .in2(_gnd_net_),
            .in3(N__16620),
            .lcout(\b2v_inst200.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_5_LC_2_7_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_5_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_5_LC_2_7_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_5_LC_2_7_6  (
            .in0(N__16621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36491),
            .ce(N__16487),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI1QM71_11_LC_2_7_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_2_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI1QM71_11_LC_2_7_7  (
            .in0(N__16358),
            .in1(N__16345),
            .in2(_gnd_net_),
            .in3(N__16568),
            .lcout(\b2v_inst200.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3T051_3_LC_2_8_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3T051_3_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3T051_3_LC_2_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNI3T051_3_LC_2_8_0  (
            .in0(N__16550),
            .in1(N__16270),
            .in2(_gnd_net_),
            .in3(N__16236),
            .lcout(\b2v_inst200.un2_count_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_3_LC_2_8_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_3_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_3_LC_2_8_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_3_LC_2_8_1  (
            .in0(N__16237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36531),
            .ce(N__16489),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50P71_0_13_LC_2_8_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50P71_0_13_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50P71_0_13_LC_2_8_2 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \b2v_inst200.count_RNI50P71_0_13_LC_2_8_2  (
            .in0(N__16553),
            .in1(N__16655),
            .in2(N__16307),
            .in3(N__16646),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIUF4N4_3_LC_2_8_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIUF4N4_3_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIUF4N4_3_LC_2_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNIUF4N4_3_LC_2_8_3  (
            .in0(N__16289),
            .in1(N__16223),
            .in2(N__16283),
            .in3(N__16436),
            .lcout(\b2v_inst200.un25_clk_100khz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3T051_0_3_LC_2_8_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3T051_0_3_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3T051_0_3_LC_2_8_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \b2v_inst200.count_RNI3T051_0_3_LC_2_8_4  (
            .in0(N__16552),
            .in1(N__16271),
            .in2(N__16262),
            .in3(N__16238),
            .lcout(\b2v_inst200.un25_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_13_LC_2_8_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_13_LC_2_8_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_13_LC_2_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_13_LC_2_8_5  (
            .in0(N__16645),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36531),
            .ce(N__16489),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50P71_13_LC_2_8_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50P71_13_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50P71_13_LC_2_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNI50P71_13_LC_2_8_6  (
            .in0(N__16551),
            .in1(N__16654),
            .in2(_gnd_net_),
            .in3(N__16644),
            .lcout(\b2v_inst200.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73351_0_5_LC_2_8_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73351_0_5_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73351_0_5_LC_2_8_7 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \b2v_inst200.count_RNI73351_0_5_LC_2_8_7  (
            .in0(N__16628),
            .in1(N__16606),
            .in2(N__16595),
            .in3(N__16549),
            .lcout(\b2v_inst200.un25_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_2_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_2_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__21275),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_2_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_2_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__18173),
            .in2(N__16867),
            .in3(N__16421),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_2_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_2_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__16863),
            .in2(N__18098),
            .in3(N__16412),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_2_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_2_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__18083),
            .in2(N__18245),
            .in3(N__16400),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_2_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_2_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__18243),
            .in2(N__18071),
            .in3(N__16391),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_2_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_2_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_2_9_5  (
            .in0(N__18149),
            .in1(N__18056),
            .in2(N__16868),
            .in3(N__16748),
            .lcout(\b2v_inst11.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_2_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_2_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__18260),
            .in2(_gnd_net_),
            .in3(N__16745),
            .lcout(\b2v_inst11.mult1_un61_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un61_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_2_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_2_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16742),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__21379),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__18521),
            .in2(N__16909),
            .in3(N__16712),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__16905),
            .in2(N__16709),
            .in3(N__16694),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__16691),
            .in2(N__16850),
            .in3(N__16676),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__16848),
            .in2(N__16673),
            .in3(N__16658),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_10_5  (
            .in0(N__16779),
            .in1(N__16916),
            .in2(N__16910),
            .in3(N__16883),
            .lcout(\b2v_inst11.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_10_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16880),
            .in3(N__16871),
            .lcout(\b2v_inst11.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_2_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_2_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18244),
            .lcout(\b2v_inst11.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16849),
            .lcout(\b2v_inst11.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_2_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_2_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_2_11_1  (
            .in0(N__21313),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_2_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_2_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21383),
            .lcout(\b2v_inst11.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21418),
            .lcout(\b2v_inst11.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16777),
            .lcout(\b2v_inst11.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_11_6  (
            .in0(N__16778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un82_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17014),
            .lcout(\b2v_inst11.mult1_un96_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__21496),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__20267),
            .in2(N__16972),
            .in3(N__17039),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__16968),
            .in2(N__17036),
            .in3(N__17027),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__17024),
            .in2(N__17015),
            .in3(N__17018),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__17013),
            .in2(N__16991),
            .in3(N__16982),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_12_5  (
            .in0(N__20225),
            .in1(N__16979),
            .in2(N__16973),
            .in3(N__16955),
            .lcout(\b2v_inst11.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16952),
            .in3(N__16943),
            .lcout(\b2v_inst11.mult1_un103_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16939),
            .lcout(\b2v_inst11.mult1_un89_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNI2EHH1_LC_2_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNI2EHH1_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNI2EHH1_LC_2_13_0 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \b2v_inst11.pwm_out_RNI2EHH1_LC_2_13_0  (
            .in0(N__17063),
            .in1(N__19812),
            .in2(N__17054),
            .in3(N__17294),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_2_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_2_13_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__19841),
            .in2(N__19816),
            .in3(N__19779),
            .lcout(),
            .ltout(\b2v_inst11.curr_state_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_2_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_2_13_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.curr_state_RNIJK34_0_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__19754),
            .in2(N__17159),
            .in3(N__30577),
            .lcout(\b2v_inst11.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst11.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_2_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_2_13_3 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \b2v_inst11.curr_state_RNIOCA3_0_LC_2_13_3  (
            .in0(N__30578),
            .in1(_gnd_net_),
            .in2(N__17156),
            .in3(N__19778),
            .lcout(\b2v_inst11.count_0_sqmuxa_i ),
            .ltout(\b2v_inst11.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_0_LC_2_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_0_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_0_LC_2_13_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst11.count_RNI_0_LC_2_13_4  (
            .in0(N__18474),
            .in1(_gnd_net_),
            .in2(N__17075),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst11.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI03G9_0_LC_2_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI03G9_0_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI03G9_0_LC_2_13_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst11.count_RNI03G9_0_LC_2_13_5  (
            .in0(N__30579),
            .in1(_gnd_net_),
            .in2(N__17072),
            .in3(N__17069),
            .lcout(\b2v_inst11.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_LC_2_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.pwm_out_LC_2_13_6 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \b2v_inst11.pwm_out_LC_2_13_6  (
            .in0(N__17062),
            .in1(N__19811),
            .in2(N__17053),
            .in3(N__17293),
            .lcout(\b2v_inst11.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36575),
            .ce(),
            .sr(N__17177));
    defparam \b2v_inst11.curr_state_RNIKEBL_0_LC_2_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIKEBL_0_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIKEBL_0_LC_2_13_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst11.curr_state_RNIKEBL_0_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__32223),
            .in2(_gnd_net_),
            .in3(N__19840),
            .lcout(\b2v_inst11.g0_i_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIMQBN_3_LC_2_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_2_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIMQBN_3_LC_2_14_0  (
            .in0(N__30693),
            .in1(N__17237),
            .in2(_gnd_net_),
            .in3(N__17245),
            .lcout(\b2v_inst11.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_3_LC_2_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_3_LC_2_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_3_LC_2_14_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_3_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17249),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36581),
            .ce(N__32180),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOC3M_13_LC_2_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_2_14_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \b2v_inst11.count_RNIOC3M_13_LC_2_14_2  (
            .in0(N__17231),
            .in1(N__17219),
            .in2(N__30726),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_13_LC_2_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_13_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_13_LC_2_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_13_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17230),
            .lcout(\b2v_inst11.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36581),
            .ce(N__32180),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOTCN_4_LC_2_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_2_14_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIOTCN_4_LC_2_14_4  (
            .in0(N__30692),
            .in1(N__17201),
            .in2(_gnd_net_),
            .in3(N__17209),
            .lcout(\b2v_inst11.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_4_LC_2_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_4_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_4_LC_2_14_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_4_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17213),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36581),
            .ce(N__32180),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_2_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_2_14_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIQ0EN_5_LC_2_14_6  (
            .in0(N__30694),
            .in1(N__17183),
            .in2(_gnd_net_),
            .in3(N__17191),
            .lcout(\b2v_inst11.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_5_LC_2_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_5_LC_2_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_5_LC_2_14_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_5_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17195),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36581),
            .ce(N__32180),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNO_0_LC_2_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_2_15_0 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \b2v_inst11.pwm_out_RNO_0_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__19846),
            .in2(N__19783),
            .in3(N__30700),
            .lcout(\b2v_inst11.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_2_LC_2_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_2_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_2_LC_2_15_1 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst11.count_RNI_2_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__18318),
            .in2(N__18358),
            .in3(N__18387),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlt6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_5_LC_2_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_5_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_5_LC_2_15_2 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \b2v_inst11.count_RNI_5_LC_2_15_2  (
            .in0(N__18285),
            .in1(N__18846),
            .in2(N__17312),
            .in3(N__18813),
            .lcout(\b2v_inst11.un79_clk_100khzlto15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_10_LC_2_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_10_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_10_LC_2_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_RNI_10_LC_2_15_3  (
            .in0(N__18703),
            .in1(N__18543),
            .in2(N__18616),
            .in3(N__18659),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_15_LC_2_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_15_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_15_LC_2_15_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \b2v_inst11.count_RNI_15_LC_2_15_4  (
            .in0(N__18969),
            .in1(_gnd_net_),
            .in2(N__17309),
            .in3(N__18933),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_8_LC_2_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_8_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_8_LC_2_15_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.count_RNI_8_LC_2_15_5  (
            .in0(N__18747),
            .in1(N__18786),
            .in2(N__17306),
            .in3(N__17303),
            .lcout(\b2v_inst11.count_RNIZ0Z_8 ),
            .ltout(\b2v_inst11.count_RNIZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNICRLO_0_LC_2_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNICRLO_0_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNICRLO_0_LC_2_15_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.curr_state_RNICRLO_0_LC_2_15_6  (
            .in0(N__30701),
            .in1(N__32222),
            .in2(N__17297),
            .in3(N__19845),
            .lcout(\b2v_inst11.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQF4M_14_LC_2_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_2_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_RNIQF4M_14_LC_2_16_0  (
            .in0(N__17282),
            .in1(N__17273),
            .in2(_gnd_net_),
            .in3(N__30691),
            .lcout(\b2v_inst11.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_14_LC_2_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_14_LC_2_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_14_LC_2_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_14_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17281),
            .lcout(\b2v_inst11.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36602),
            .ce(N__32179),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIS3FN_6_LC_2_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_2_16_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIS3FN_6_LC_2_16_2  (
            .in0(N__30698),
            .in1(N__17255),
            .in2(_gnd_net_),
            .in3(N__17263),
            .lcout(\b2v_inst11.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_6_LC_2_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_6_LC_2_16_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_6_LC_2_16_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_6_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17267),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36602),
            .ce(N__32179),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNISI5M_15_LC_2_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNISI5M_15_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNISI5M_15_LC_2_16_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNISI5M_15_LC_2_16_4  (
            .in0(N__17393),
            .in1(N__30690),
            .in2(_gnd_net_),
            .in3(N__17401),
            .lcout(\b2v_inst11.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_15_LC_2_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_15_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_15_LC_2_16_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_15_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17405),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36602),
            .ce(N__32179),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIU6GN_7_LC_2_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_2_16_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIU6GN_7_LC_2_16_6  (
            .in0(N__30699),
            .in1(N__17375),
            .in2(_gnd_net_),
            .in3(N__17383),
            .lcout(\b2v_inst11.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_7_LC_2_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_7_LC_2_16_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_7_LC_2_16_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_7_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17387),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36602),
            .ce(N__32179),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_4_1_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_4_1_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_4_1_3  (
            .in0(_gnd_net_),
            .in1(N__19482),
            .in2(_gnd_net_),
            .in3(N__19461),
            .lcout(\b2v_inst200.N_282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI_0_LC_4_1_4 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI_0_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI_0_LC_4_1_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst16.curr_state_RNI_0_LC_4_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17698),
            .lcout(\b2v_inst16.N_3079_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_en_LC_4_1_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_en_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_en_LC_4_1_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.count_en_LC_4_1_7  (
            .in0(_gnd_net_),
            .in1(N__19481),
            .in2(_gnd_net_),
            .in3(N__32219),
            .lcout(\b2v_inst200.count_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_4_2_1 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_4_2_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \b2v_inst16.curr_state_RNIKEBL_1_LC_4_2_1  (
            .in0(N__17614),
            .in1(N__27720),
            .in2(_gnd_net_),
            .in3(N__32220),
            .lcout(\b2v_inst16.count_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_0_LC_4_2_3 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_0_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_0_LC_4_2_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_0_LC_4_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29492),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIUCAD1_1_0_LC_4_2_4 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIUCAD1_1_0_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIUCAD1_1_0_LC_4_2_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst16.curr_state_RNIUCAD1_1_0_LC_4_2_4  (
            .in0(N__27721),
            .in1(N__17569),
            .in2(_gnd_net_),
            .in3(N__27759),
            .lcout(\b2v_inst16.curr_state_7_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.delayed_vddq_pwrgd_e_0_RNI8HF43_LC_4_3_0 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_e_0_RNI8HF43_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_e_0_RNI8HF43_LC_4_3_0 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_e_0_RNI8HF43_LC_4_3_0  (
            .in0(N__17744),
            .in1(N__17750),
            .in2(N__27734),
            .in3(N__33653),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.delayed_vddq_pwrgd_e_0_LC_4_3_1 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_e_0_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_e_0_LC_4_3_1 .LUT_INIT=16'b1100111011111111;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_e_0_LC_4_3_1  (
            .in0(N__19520),
            .in1(N__27722),
            .in2(N__30689),
            .in3(N__33578),
            .lcout(\b2v_inst16.delayed_vddq_pwrgd_eZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36208),
            .ce(N__17743),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIIRL22_0_LC_4_3_5 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIIRL22_0_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIIRL22_0_LC_4_3_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst16.curr_state_RNIIRL22_0_LC_4_3_5  (
            .in0(N__27689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32221),
            .lcout(\b2v_inst16.delayed_vddq_pwrgd_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIMPKG1_0_LC_4_3_6 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIMPKG1_0_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIMPKG1_0_LC_4_3_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \b2v_inst16.curr_state_RNIMPKG1_0_LC_4_3_6  (
            .in0(_gnd_net_),
            .in1(N__27688),
            .in2(_gnd_net_),
            .in3(N__30627),
            .lcout(\b2v_inst16.N_26 ),
            .ltout(\b2v_inst16.N_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_4_3_7 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_4_3_7 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_4_3_7  (
            .in0(N__17570),
            .in1(N__17488),
            .in2(N__17468),
            .in3(N__17814),
            .lcout(\b2v_inst16.count_rst_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNILO901_0_13_LC_4_4_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILO901_0_13_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILO901_0_13_LC_4_4_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst16.count_RNILO901_0_13_LC_4_4_0  (
            .in0(N__17419),
            .in1(N__17452),
            .in2(N__17942),
            .in3(N__17807),
            .lcout(\b2v_inst16.count_4_i_a3_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIJP141_14_LC_4_4_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIJP141_14_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIJP141_14_LC_4_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNIJP141_14_LC_4_4_1  (
            .in0(N__17426),
            .in1(N__20077),
            .in2(_gnd_net_),
            .in3(N__17437),
            .lcout(\b2v_inst16.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_14_LC_4_4_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_14_LC_4_4_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_14_LC_4_4_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_14_LC_4_4_2  (
            .in0(N__17438),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36291),
            .ce(N__20078),
            .sr(N__17892));
    defparam \b2v_inst16.count_RNIFJV31_12_LC_4_4_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIFJV31_12_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIFJV31_12_LC_4_4_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNIFJV31_12_LC_4_4_3  (
            .in0(N__17948),
            .in1(N__20075),
            .in2(_gnd_net_),
            .in3(N__17959),
            .lcout(\b2v_inst16.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_12_LC_4_4_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_12_LC_4_4_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_12_LC_4_4_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_12_LC_4_4_4  (
            .in0(N__17960),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36291),
            .ce(N__20078),
            .sr(N__17892));
    defparam \b2v_inst16.count_RNILO901_13_LC_4_4_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILO901_13_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILO901_13_LC_4_4_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNILO901_13_LC_4_4_5  (
            .in0(N__17912),
            .in1(N__20076),
            .in2(_gnd_net_),
            .in3(N__17923),
            .lcout(\b2v_inst16.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_13_LC_4_4_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_13_LC_4_4_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_13_LC_4_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_13_LC_4_4_6  (
            .in0(N__17924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36291),
            .ce(N__20078),
            .sr(N__17892));
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_4_4_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_4_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNIF7UJ1_3_LC_4_4_7  (
            .in0(N__17840),
            .in1(N__20079),
            .in2(_gnd_net_),
            .in3(N__17828),
            .lcout(\b2v_inst16.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_7_LC_4_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_7_LC_4_5_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_7_LC_4_5_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \b2v_inst11.dutycycle_7_LC_4_5_0  (
            .in0(N__33884),
            .in1(N__25346),
            .in2(N__22841),
            .in3(N__17786),
            .lcout(\b2v_inst11.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36314),
            .ce(),
            .sr(N__31031));
    defparam \b2v_inst11.dutycycle_RNIRH7VD_7_LC_4_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIRH7VD_7_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIRH7VD_7_LC_4_5_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIRH7VD_7_LC_4_5_1  (
            .in0(N__17785),
            .in1(N__33883),
            .in2(N__22840),
            .in3(N__25345),
            .lcout(\b2v_inst11.dutycycleZ1Z_3 ),
            .ltout(\b2v_inst11.dutycycleZ1Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_7_LC_4_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_7_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_7_LC_4_5_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_7_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17777),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_4_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_4_5_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_7_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__22631),
            .in2(_gnd_net_),
            .in3(N__22877),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_LC_4_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_4_5_4 .LUT_INIT=16'b1011010011010010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_LC_4_5_4  (
            .in0(N__29972),
            .in1(N__22775),
            .in2(N__17774),
            .in3(N__19715),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_4_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_4_6_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_3_LC_4_6_0  (
            .in0(N__20330),
            .in1(N__23437),
            .in2(N__30185),
            .in3(N__24629),
            .lcout(\b2v_inst11.g3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIN8NR1_1_LC_4_6_1 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIN8NR1_1_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIN8NR1_1_LC_4_6_1 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \b2v_inst16.curr_state_RNIN8NR1_1_LC_4_6_1  (
            .in0(N__17996),
            .in1(N__17984),
            .in2(_gnd_net_),
            .in3(N__30631),
            .lcout(\b2v_inst16.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_10_LC_4_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_4_6_2 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_10_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__22769),
            .in2(N__22659),
            .in3(N__23563),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_44_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_6_LC_4_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_6_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_6_LC_4_6_3 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_6_LC_4_6_3  (
            .in0(N__19538),
            .in1(N__18035),
            .in2(N__17972),
            .in3(N__29968),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_11_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_13_LC_4_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_13_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_13_LC_4_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_13_LC_4_6_4  (
            .in0(N__22635),
            .in1(N__24955),
            .in2(N__23099),
            .in3(N__23564),
            .lcout(\b2v_inst11.un2_count_clk_17_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_4_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_4_6_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_6_LC_4_6_5  (
            .in0(N__22768),
            .in1(N__25414),
            .in2(_gnd_net_),
            .in3(N__29967),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_4_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_4_6_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_3_LC_4_6_6  (
            .in0(N__25415),
            .in1(N__23436),
            .in2(_gnd_net_),
            .in3(N__24628),
            .lcout(\b2v_inst11.N_355 ),
            .ltout(\b2v_inst11.N_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_4_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_4_6_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_15_LC_4_6_7  (
            .in0(N__22770),
            .in1(N__17969),
            .in2(N__17963),
            .in3(N__24712),
            .lcout(\b2v_inst11.N_363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_4_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_4_7_0 .LUT_INIT=16'b1011111100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_8_LC_4_7_0  (
            .in0(N__24598),
            .in1(N__25422),
            .in2(N__25140),
            .in3(N__23572),
            .lcout(\b2v_inst11.un1_dutycycle_53_55_1_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_11_LC_4_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_11_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_11_LC_4_7_2 .LUT_INIT=16'b0000000101011111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_11_LC_4_7_2  (
            .in0(N__25080),
            .in1(N__22779),
            .in2(N__22658),
            .in3(N__25216),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_6Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_8_LC_4_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_8_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_8_LC_4_7_3 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_8_LC_4_7_3  (
            .in0(N__19721),
            .in1(N__18044),
            .in2(N__18038),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_4_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_4_7_4 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_10_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__24597),
            .in2(N__22657),
            .in3(N__23571),
            .lcout(\b2v_inst11.un1_dutycycle_53_50_a0_1 ),
            .ltout(\b2v_inst11.un1_dutycycle_53_50_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_4_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_4_7_5 .LUT_INIT=16'b0011000000110001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_6_LC_4_7_5  (
            .in0(N__22780),
            .in1(N__29965),
            .in2(N__18029),
            .in3(N__18116),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_6_LC_4_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_6_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_6_LC_4_7_6 .LUT_INIT=16'b1111101100000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_6_LC_4_7_6  (
            .in0(N__19636),
            .in1(N__19616),
            .in2(N__18026),
            .in3(N__24644),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_4_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_4_8_0 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_12_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(N__23573),
            .in2(N__22665),
            .in3(N__25085),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_12 ),
            .ltout(\b2v_inst11.dutycycle_RNI_1Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_6_LC_4_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_6_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_6_LC_4_8_1 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_6_LC_4_8_1  (
            .in0(N__19651),
            .in1(N__18020),
            .in2(N__18023),
            .in3(N__18005),
            .lcout(\b2v_inst11.dutycycle_RNI_8Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_4_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_4_8_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_6_LC_4_8_2  (
            .in0(N__29961),
            .in1(N__24630),
            .in2(_gnd_net_),
            .in3(N__25426),
            .lcout(\b2v_inst11.un1_dutycycle_53_4_1 ),
            .ltout(\b2v_inst11.un1_dutycycle_53_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_6_LC_4_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_6_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_6_LC_4_8_3 .LUT_INIT=16'b0000000011110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_6_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__18014),
            .in2(N__18008),
            .in3(N__18004),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_7Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_13_LC_4_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_4_8_4 .LUT_INIT=16'b1100110000111100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_13_LC_4_8_4  (
            .in0(N__24956),
            .in1(N__25086),
            .in2(N__18119),
            .in3(N__19652),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_7_LC_4_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_7_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_7_LC_4_8_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_7_LC_4_8_5  (
            .in0(N__25425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25139),
            .lcout(\b2v_inst11.dutycycle_RNI_9Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_4_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_4_8_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_11_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22666),
            .in3(N__25217),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_46_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_4_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_4_8_7 .LUT_INIT=16'b0011110011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_14_LC_4_8_7  (
            .in0(N__23091),
            .in1(N__19661),
            .in2(N__18110),
            .in3(N__18107),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21236),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19868),
            .in3(N__18086),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__19696),
            .in2(N__18212),
            .in3(N__18074),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__32052),
            .in2(N__19901),
            .in3(N__18059),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__19889),
            .in2(N__32059),
            .in3(N__18047),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_9_5  (
            .in0(N__18231),
            .in1(N__20171),
            .in2(N__19877),
            .in3(N__18251),
            .lcout(\b2v_inst11.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_6 .LUT_INIT=16'b0011000011001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__20183),
            .in2(N__20195),
            .in3(N__18248),
            .lcout(\b2v_inst11.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_9_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_9_7  (
            .in0(N__19695),
            .in1(N__19697),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un1_vddq_en_LC_4_10_0 .C_ON=1'b0;
    defparam \b2v_inst16.un1_vddq_en_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un1_vddq_en_LC_4_10_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst16.un1_vddq_en_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__33646),
            .in2(_gnd_net_),
            .in3(N__18203),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21497),
            .lcout(\b2v_inst11.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21232),
            .lcout(\b2v_inst11.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18161),
            .lcout(\b2v_inst11.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21274),
            .lcout(\b2v_inst11.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_5_LC_4_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_5_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_5_LC_4_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_5_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35182),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21347),
            .lcout(\b2v_inst11.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18512),
            .lcout(\b2v_inst11.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_4_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_4_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_4_11_0  (
            .in0(N__18482),
            .in1(N__18443),
            .in2(N__19223),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5980_i ),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_4_11_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_4_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__18407),
            .in2(N__20276),
            .in3(N__18437),
            .lcout(\b2v_inst11.N_5981_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_0 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_4_11_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_4_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__20282),
            .in2(N__18371),
            .in3(N__18401),
            .lcout(\b2v_inst11.N_5982_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_1 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_4_11_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_4_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_4_11_3  (
            .in0(N__18362),
            .in1(N__20252),
            .in2(N__18335),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5983_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_2 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_4_11_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_4_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_4_11_4  (
            .in0(N__18326),
            .in1(N__19907),
            .in2(N__18302),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5984_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_3 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_4_11_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_4_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_4_11_5  (
            .in0(N__18293),
            .in1(N__20258),
            .in2(N__18269),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5985_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_4 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_4_11_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_4_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(N__18830),
            .in2(N__20291),
            .in3(N__18857),
            .lcout(\b2v_inst11.N_5986_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_5 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_4_11_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_4_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_4_11_7  (
            .in0(N__18824),
            .in1(N__18797),
            .in2(N__19925),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5987_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_6 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_4_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_4_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__18896),
            .in2(N__18761),
            .in3(N__18791),
            .lcout(\b2v_inst11.N_5988_i ),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_4_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_4_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__20201),
            .in2(N__18728),
            .in3(N__18752),
            .lcout(\b2v_inst11.N_5989_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_8 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_4_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_4_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__18719),
            .in2(N__18677),
            .in3(N__18707),
            .lcout(\b2v_inst11.N_5990_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_9 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_4_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_4_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__18668),
            .in2(N__18629),
            .in3(N__18658),
            .lcout(\b2v_inst11.N_5991_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_10 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_4_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_4_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_4_12_4  (
            .in0(N__18620),
            .in1(N__18590),
            .in2(N__18578),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5992_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_11 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_4_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_4_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(N__18569),
            .in2(N__18530),
            .in3(N__18557),
            .lcout(\b2v_inst11.N_5993_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_12 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_4_12_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_4_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(N__18986),
            .in2(N__18953),
            .in3(N__18977),
            .lcout(\b2v_inst11.N_5994_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_13 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_4_12_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_4_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_4_12_7  (
            .in0(N__18941),
            .in1(N__18917),
            .in2(N__18908),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5995_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_14 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18899),
            .lcout(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20241),
            .lcout(\b2v_inst11.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19174),
            .lcout(\b2v_inst11.mult1_un110_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__21110),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__18890),
            .in2(N__19051),
            .in3(N__18878),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__19047),
            .in2(N__18875),
            .in3(N__18860),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__19097),
            .in2(N__20246),
            .in3(N__19085),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__20245),
            .in2(N__19082),
            .in3(N__19067),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_14_5  (
            .in0(N__19169),
            .in1(N__19064),
            .in2(N__19052),
            .in3(N__19034),
            .lcout(\b2v_inst11.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19031),
            .in3(N__19016),
            .lcout(\b2v_inst11.mult1_un110_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un110_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19013),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__21140),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__19937),
            .in2(N__19132),
            .in3(N__19010),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__19128),
            .in2(N__19007),
            .in3(N__18998),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__18995),
            .in2(N__19175),
            .in3(N__18989),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__19173),
            .in2(N__19151),
            .in3(N__19142),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_15_5  (
            .in0(N__20432),
            .in1(N__19139),
            .in2(N__19133),
            .in3(N__19115),
            .lcout(\b2v_inst11.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19112),
            .in3(N__19103),
            .lcout(\b2v_inst11.mult1_un117_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19100),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__30183),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_16_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__20498),
            .in2(N__19243),
            .in3(N__20530),
            .lcout(G_2814),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_16_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__19239),
            .in2(N__20597),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_16_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__20531),
            .in2(N__20585),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_16_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__20573),
            .in2(N__20539),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_16_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__20564),
            .in2(N__19244),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_16_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20555),
            .in3(N__19226),
            .lcout(\b2v_inst11.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_1_0 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_1_0 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_1_0  (
            .in0(N__19484),
            .in1(N__19463),
            .in2(_gnd_net_),
            .in3(N__19181),
            .lcout(),
            .ltout(\b2v_inst200.N_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNILNOU4_0_LC_5_1_1 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNILNOU4_0_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNILNOU4_0_LC_5_1_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst200.curr_state_RNILNOU4_0_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__19397),
            .in2(N__19211),
            .in3(N__30575),
            .lcout(\b2v_inst200.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_1_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_1_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19208),
            .in3(N__19361),
            .lcout(N_411),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNIMK8L4_1_LC_5_1_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNIMK8L4_1_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNIMK8L4_1_LC_5_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.curr_state_RNIMK8L4_1_LC_5_1_3  (
            .in0(N__19250),
            .in1(N__19202),
            .in2(_gnd_net_),
            .in3(N__30576),
            .lcout(\b2v_inst200.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI_1_LC_5_1_4 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI_1_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI_1_LC_5_1_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst200.curr_state_RNI_1_LC_5_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19205),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.N_3031_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_1_5 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_1_5 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_1_5  (
            .in0(N__29488),
            .in1(N__19310),
            .in2(N__19273),
            .in3(N__19294),
            .lcout(\b2v_inst200.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_1_6 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_1_6 .LUT_INIT=16'b0000010010011101;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_1_6  (
            .in0(N__19311),
            .in1(N__19290),
            .in2(N__19196),
            .in3(N__29487),
            .lcout(\b2v_inst200.m6_i_0 ),
            .ltout(\b2v_inst200.m6_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_0_LC_5_1_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_0_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_0_LC_5_1_7 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \b2v_inst200.curr_state_0_LC_5_1_7  (
            .in0(_gnd_net_),
            .in1(N__19483),
            .in2(N__19466),
            .in3(N__19462),
            .lcout(\b2v_inst200.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36209),
            .ce(N__32173),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_2_LC_5_2_1 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_2_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_2_LC_5_2_1 .LUT_INIT=16'b0000001000110011;
    LogicCell40 \b2v_inst200.curr_state_2_LC_5_2_1  (
            .in0(N__29491),
            .in1(N__19271),
            .in2(N__19349),
            .in3(N__19332),
            .lcout(\b2v_inst200.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36368),
            .ce(N__32175),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_2_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_2_2 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_2_2  (
            .in0(N__19334),
            .in1(N__19344),
            .in2(N__19274),
            .in3(N__29489),
            .lcout(),
            .ltout(\b2v_inst200.i4_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNINL8L4_2_LC_5_2_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNINL8L4_2_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNINL8L4_2_LC_5_2_3 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \b2v_inst200.curr_state_RNINL8L4_2_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__19391),
            .in2(N__19385),
            .in3(N__30632),
            .lcout(\b2v_inst200.curr_state_i_2 ),
            .ltout(\b2v_inst200.curr_state_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_2_4 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_2_4 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_2_4  (
            .in0(N__30633),
            .in1(N__19319),
            .in2(N__19382),
            .in3(N__19348),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_2_5 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_2_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst200.curr_state_RNI_0_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(N__19312),
            .in2(_gnd_net_),
            .in3(N__19360),
            .lcout(\b2v_inst200.N_205 ),
            .ltout(\b2v_inst200.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_2_6 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_2_6 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \b2v_inst200.HDA_SDO_ATP_LC_5_2_6  (
            .in0(N__19333),
            .in1(_gnd_net_),
            .in2(N__19322),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.HDA_SDO_ATP_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36368),
            .ce(N__32175),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_1_LC_5_2_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_1_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_1_LC_5_2_7 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \b2v_inst200.curr_state_1_LC_5_2_7  (
            .in0(N__29490),
            .in1(N__19313),
            .in2(N__19295),
            .in3(N__19272),
            .lcout(\b2v_inst200.curr_state_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36368),
            .ce(N__32175),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_5_3_0 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_5_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_2_c_RNO_LC_5_3_0  (
            .in0(N__20770),
            .in1(N__20611),
            .in2(N__20789),
            .in3(N__20626),
            .lcout(\b2v_inst20.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_5_3_1 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_5_3_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_3_c_RNO_LC_5_3_1  (
            .in0(N__20707),
            .in1(N__20740),
            .in2(N__20726),
            .in3(N__20755),
            .lcout(\b2v_inst20.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_5_3_2 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_5_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_4_c_RNO_LC_5_3_2  (
            .in0(N__20692),
            .in1(N__20659),
            .in2(N__20678),
            .in3(N__20911),
            .lcout(\b2v_inst20.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_5_3_3 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_5_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_5_c_RNO_LC_5_3_3  (
            .in0(N__20878),
            .in1(N__20848),
            .in2(N__20897),
            .in3(N__20863),
            .lcout(\b2v_inst20.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_5_3_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_5_3_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_0_LC_5_3_5  (
            .in0(N__28178),
            .in1(N__28130),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIUCAD1_0_LC_5_3_7 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIUCAD1_0_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIUCAD1_0_LC_5_3_7 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \b2v_inst16.curr_state_RNIUCAD1_0_LC_5_3_7  (
            .in0(N__19519),
            .in1(N__33577),
            .in2(_gnd_net_),
            .in3(N__30543),
            .lcout(\b2v_inst16.curr_state_RNIUCAD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_LC_5_4_0 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_0_c_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_LC_5_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22334),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(\b2v_inst20.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_1_c_LC_5_4_1 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_1_c_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_LC_5_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22220),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_0 ),
            .carryout(\b2v_inst20.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_LC_5_4_2 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_2_c_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_LC_5_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_2_c_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__19496),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_1 ),
            .carryout(\b2v_inst20.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_LC_5_4_3 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_3_c_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_LC_5_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_3_c_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(N__19490),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_2 ),
            .carryout(\b2v_inst20.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_LC_5_4_4 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_4_c_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_LC_5_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_4_c_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(N__19553),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_3 ),
            .carryout(\b2v_inst20.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_LC_5_4_5 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_5_c_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_LC_5_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_5_c_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(N__19547),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_4 ),
            .carryout(\b2v_inst20.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_LC_5_4_6 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_6_c_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_LC_5_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_6_c_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__19604),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_5 ),
            .carryout(\b2v_inst20.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_LC_5_4_7 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_7_c_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_LC_5_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_7_c_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__20927),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_6 ),
            .carryout(b2v_inst20_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_5_5_0.C_ON=1'b0;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_5_5_0.SEQ_MODE=4'b0000;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_5_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_5_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19541),
            .lcout(b2v_inst20_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_5_1 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_LC_5_5_1  (
            .in0(N__23545),
            .in1(N__22777),
            .in2(N__25449),
            .in3(N__24620),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_39_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_5_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_5_5_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_7_LC_5_5_2  (
            .in0(N__19537),
            .in1(N__19598),
            .in2(N__19526),
            .in3(N__22908),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_5_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_5_5_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_13_LC_5_5_3  (
            .in0(N__22642),
            .in1(N__24943),
            .in2(N__19523),
            .in3(N__22778),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_5_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_5_5_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_10_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__19610),
            .in2(_gnd_net_),
            .in3(N__22641),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_5_5_5 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_5_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_6_c_RNO_LC_5_5_5  (
            .in0(N__20833),
            .in1(N__20818),
            .in2(N__21005),
            .in3(N__20803),
            .lcout(\b2v_inst20.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_5_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_5_5_6 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_8_LC_5_5_6  (
            .in0(N__22776),
            .in1(N__23544),
            .in2(N__24631),
            .in3(N__29966),
            .lcout(\b2v_inst11.un1_dutycycle_53_39_d_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNITSFK3_10_LC_5_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITSFK3_10_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITSFK3_10_LC_5_6_0 .LUT_INIT=16'b0000001011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNITSFK3_10_LC_5_6_0  (
            .in0(N__34252),
            .in1(N__25532),
            .in2(N__25496),
            .in3(N__22646),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNITSFK3Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI9LPN6_10_LC_5_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI9LPN6_10_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI9LPN6_10_LC_5_6_1 .LUT_INIT=16'b0010001111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI9LPN6_10_LC_5_6_1  (
            .in0(N__24995),
            .in1(N__27650),
            .in2(N__19592),
            .in3(N__34812),
            .lcout(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_10 ),
            .ltout(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI3ER99_10_LC_5_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI3ER99_10_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI3ER99_10_LC_5_6_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI3ER99_10_LC_5_6_2  (
            .in0(N__31226),
            .in1(N__19576),
            .in2(N__19589),
            .in3(N__22555),
            .lcout(\b2v_inst11.dutycycleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_10_LC_5_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_10_LC_5_6_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_10_LC_5_6_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \b2v_inst11.dutycycle_10_LC_5_6_3  (
            .in0(N__22556),
            .in1(N__19586),
            .in2(N__19580),
            .in3(N__31227),
            .lcout(\b2v_inst11.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36604),
            .ce(),
            .sr(N__31043));
    defparam \b2v_inst11.dutycycle_RNIQ9K59_9_LC_5_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQ9K59_9_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQ9K59_9_LC_5_6_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIQ9K59_9_LC_5_6_4  (
            .in0(N__31225),
            .in1(N__19675),
            .in2(N__19562),
            .in3(N__22684),
            .lcout(\b2v_inst11.dutycycleZ0Z_1 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNITSFK3_9_LC_5_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITSFK3_9_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITSFK3_9_LC_5_6_5 .LUT_INIT=16'b0001111100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNITSFK3_9_LC_5_6_5  (
            .in0(N__25531),
            .in1(N__25492),
            .in2(N__19568),
            .in3(N__34251),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNITSFK3Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI9LPN6_9_LC_5_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI9LPN6_9_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI9LPN6_9_LC_5_6_6 .LUT_INIT=16'b0101010111011111;
    LogicCell40 \b2v_inst11.dutycycle_RNI9LPN6_9_LC_5_6_6  (
            .in0(N__34811),
            .in1(N__24994),
            .in2(N__19565),
            .in3(N__27646),
            .lcout(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_9 ),
            .ltout(\b2v_inst11.dutycycle_RNI9LPN6Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_9_LC_5_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_9_LC_5_6_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_9_LC_5_6_7 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.dutycycle_9_LC_5_6_7  (
            .in0(N__22685),
            .in1(N__19676),
            .in2(N__19679),
            .in3(N__31228),
            .lcout(\b2v_inst11.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36604),
            .ce(),
            .sr(N__31043));
    defparam \b2v_inst11.dutycycle_RNI_4_LC_5_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_LC_5_7_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__24608),
            .in2(_gnd_net_),
            .in3(N__22774),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_30_a1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_5_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_5_7_1 .LUT_INIT=16'b1111111100001110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_7_LC_5_7_1  (
            .in0(N__23542),
            .in1(N__22637),
            .in2(N__19664),
            .in3(N__22912),
            .lcout(\b2v_inst11.un1_dutycycle_53_44_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_5_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_5_7_2 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_13_LC_5_7_2  (
            .in0(N__25138),
            .in1(N__25081),
            .in2(N__22660),
            .in3(N__24916),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_13_LC_5_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_13_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_13_LC_5_7_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_13_LC_5_7_3  (
            .in0(N__19625),
            .in1(N__19650),
            .in2(N__19655),
            .in3(N__19637),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_6_LC_5_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_6_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_6_LC_5_7_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_6_LC_5_7_4  (
            .in0(N__25423),
            .in1(N__22773),
            .in2(N__25142),
            .in3(N__29964),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_5_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_5_7_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_4_LC_5_7_5  (
            .in0(N__22772),
            .in1(N__25134),
            .in2(N__24627),
            .in3(N__25424),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_5_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_5_7_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_8_LC_5_7_6  (
            .in0(_gnd_net_),
            .in1(N__23541),
            .in2(N__25141),
            .in3(N__22771),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_8 ),
            .ltout(\b2v_inst11.dutycycle_RNI_3Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_5_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_5_7_7 .LUT_INIT=16'b0000111100000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_11_LC_5_7_7  (
            .in0(N__20921),
            .in1(N__25215),
            .in2(N__19619),
            .in3(N__22636),
            .lcout(\b2v_inst11.un1_dutycycle_53_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_5_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_5_8_0 .LUT_INIT=16'b0000111101111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_11_LC_5_8_0  (
            .in0(N__25060),
            .in1(N__22650),
            .in2(N__22795),
            .in3(N__25197),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_LC_5_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_5_8_1 .LUT_INIT=16'b1111111010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_LC_5_8_1  (
            .in0(N__22913),
            .in1(N__23553),
            .in2(N__23438),
            .in3(N__24555),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_7 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_5_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_5_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_5_LC_5_8_2  (
            .in0(N__22788),
            .in1(N__35192),
            .in2(N__19706),
            .in3(N__29941),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_LC_5_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_5_8_3 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_LC_5_8_3  (
            .in0(N__23434),
            .in1(N__30168),
            .in2(N__31378),
            .in3(N__24557),
            .lcout(\b2v_inst11.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_5_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_5_8_4 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_0_LC_5_8_4  (
            .in0(N__24556),
            .in1(N__31365),
            .in2(_gnd_net_),
            .in3(N__30167),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_12_LC_5_8_5  (
            .in0(N__21035),
            .in1(N__23554),
            .in2(N__25088),
            .in3(N__22789),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_5_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_5_8_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_13_LC_5_8_6  (
            .in0(N__25061),
            .in1(N__19703),
            .in2(N__23095),
            .in3(N__24917),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21601),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20153),
            .in3(N__19682),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19739),
            .in3(N__19892),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__32048),
            .in2(N__19730),
            .in3(N__19883),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19880),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_9_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_9_5  (
            .in0(N__20169),
            .in1(N__20170),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_5_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_5_9_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21602),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_9_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_15_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24713),
            .in3(N__19859),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_0_LC_5_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_0_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.curr_state_0_LC_5_10_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \b2v_inst11.curr_state_0_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__19850),
            .in2(N__19817),
            .in3(N__19787),
            .lcout(\b2v_inst11.curr_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36652),
            .ce(N__32184),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21584),
            .in3(N__21558),
            .lcout(\b2v_inst11.mult1_un47_sum_s_4_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_2 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__21582),
            .in2(N__21563),
            .in3(N__21538),
            .lcout(\b2v_inst11.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_3 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_3  (
            .in0(N__21583),
            .in1(_gnd_net_),
            .in2(N__21542),
            .in3(N__21562),
            .lcout(\b2v_inst11.mult1_un40_sum_i_5 ),
            .ltout(\b2v_inst11.mult1_un40_sum_i_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_5_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_5_10_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20186),
            .in3(N__20182),
            .lcout(\b2v_inst11.mult1_un47_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_5_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_5_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21578),
            .lcout(\b2v_inst11.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_5_10_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_5_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNI4M8F1_10_LC_5_10_7  (
            .in0(N__20144),
            .in1(N__20123),
            .in2(_gnd_net_),
            .in3(N__20107),
            .lcout(\b2v_inst16.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21109),
            .lcout(\b2v_inst11.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIANKU4_14_LC_5_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIANKU4_14_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIANKU4_14_LC_5_11_2 .LUT_INIT=16'b1110111111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIANKU4_14_LC_5_11_2  (
            .in0(N__25322),
            .in1(N__24993),
            .in2(N__34286),
            .in3(N__23087),
            .lcout(\b2v_inst11.N_155_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_5_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_5_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20444),
            .lcout(\b2v_inst11.mult1_un117_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_4 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_4  (
            .in0(N__32813),
            .in1(N__27464),
            .in2(N__30688),
            .in3(N__27533),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21836),
            .lcout(\b2v_inst11.un85_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21745),
            .lcout(\b2v_inst11.mult1_un124_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22124),
            .lcout(\b2v_inst11.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20540),
            .lcout(\b2v_inst11.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21139),
            .lcout(\b2v_inst11.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21454),
            .lcout(\b2v_inst11.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21646),
            .lcout(\b2v_inst11.mult1_un131_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_12_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21962),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20240),
            .lcout(\b2v_inst11.mult1_un103_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_12_7  (
            .in0(N__21185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__21529),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__20318),
            .in2(N__20510),
            .in3(N__20312),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__21757),
            .in2(N__21704),
            .in3(N__20309),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__20471),
            .in2(N__21746),
            .in3(N__20306),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__21744),
            .in2(N__20456),
            .in3(N__20303),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_13_5  (
            .in0(N__21641),
            .in1(N__20350),
            .in2(N__20339),
            .in3(N__20300),
            .lcout(\b2v_inst11.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_13_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20378),
            .in3(N__20297),
            .lcout(\b2v_inst11.mult1_un131_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un131_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_5_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_5_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20294),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__21184),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__20492),
            .in2(N__20395),
            .in3(N__20483),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__20391),
            .in2(N__20480),
            .in3(N__20465),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__20462),
            .in2(N__20440),
            .in3(N__20447),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__20436),
            .in2(N__20414),
            .in3(N__20405),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_14_5  (
            .in0(N__21736),
            .in1(N__20402),
            .in2(N__20396),
            .in3(N__20369),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20366),
            .in3(N__20357),
            .lcout(\b2v_inst11.mult1_un124_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un124_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20354),
            .in3(N__20351),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_5_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_5_15_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_1_LC_5_15_0  (
            .in0(N__33305),
            .in1(N__31369),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.g3_0 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__30038),
            .in2(N__22090),
            .in3(N__20588),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__22086),
            .in2(N__22010),
            .in3(N__20576),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__21989),
            .in2(N__22120),
            .in3(N__20567),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__22116),
            .in2(N__21974),
            .in3(N__20558),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_15_5  (
            .in0(N__20535),
            .in1(N__21923),
            .in2(N__22091),
            .in3(N__20546),
            .lcout(\b2v_inst11.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22148),
            .in3(N__20543),
            .lcout(\b2v_inst11.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21727),
            .lcout(\b2v_inst11.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_5_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_5_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31379),
            .lcout(\b2v_inst11.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_1_c_LC_6_2_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_6_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_c_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(N__22379),
            .in2(N__22358),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(\b2v_inst20.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_6_2_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_6_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(N__24239),
            .in2(_gnd_net_),
            .in3(N__20645),
            .lcout(\b2v_inst20.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_1 ),
            .carryout(\b2v_inst20.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_6_2_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_6_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(N__24128),
            .in2(_gnd_net_),
            .in3(N__20642),
            .lcout(\b2v_inst20.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_2 ),
            .carryout(\b2v_inst20.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_6_2_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_6_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(N__22283),
            .in2(_gnd_net_),
            .in3(N__20639),
            .lcout(\b2v_inst20.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_3 ),
            .carryout(\b2v_inst20.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_6_2_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_6_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(N__22310),
            .in2(_gnd_net_),
            .in3(N__20636),
            .lcout(\b2v_inst20.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_4 ),
            .carryout(\b2v_inst20.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_6_2_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_6_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(N__22400),
            .in2(_gnd_net_),
            .in3(N__20633),
            .lcout(\b2v_inst20.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_5 ),
            .carryout(\b2v_inst20.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_7_LC_6_2_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_7_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_7_LC_6_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_7_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(N__22234),
            .in2(_gnd_net_),
            .in3(N__20630),
            .lcout(\b2v_inst20.counterZ0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_6 ),
            .carryout(\b2v_inst20.counter_1_cry_7 ),
            .clk(N__36193),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_8_LC_6_2_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_8_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_8_LC_6_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_8_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(N__20627),
            .in2(_gnd_net_),
            .in3(N__20615),
            .lcout(\b2v_inst20.counterZ0Z_8 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_7 ),
            .carryout(\b2v_inst20.counter_1_cry_8 ),
            .clk(N__36193),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_9_LC_6_3_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_9_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_9_LC_6_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_9_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__20612),
            .in2(_gnd_net_),
            .in3(N__20600),
            .lcout(\b2v_inst20.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\b2v_inst20.counter_1_cry_9 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_10_LC_6_3_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_10_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_10_LC_6_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_10_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__20788),
            .in2(_gnd_net_),
            .in3(N__20774),
            .lcout(\b2v_inst20.counterZ0Z_10 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_9 ),
            .carryout(\b2v_inst20.counter_1_cry_10 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_11_LC_6_3_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_11_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_11_LC_6_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_11_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__20771),
            .in2(_gnd_net_),
            .in3(N__20759),
            .lcout(\b2v_inst20.counterZ0Z_11 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_10 ),
            .carryout(\b2v_inst20.counter_1_cry_11 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_12_LC_6_3_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_12_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_12_LC_6_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_12_LC_6_3_3  (
            .in0(_gnd_net_),
            .in1(N__20756),
            .in2(_gnd_net_),
            .in3(N__20744),
            .lcout(\b2v_inst20.counterZ0Z_12 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_11 ),
            .carryout(\b2v_inst20.counter_1_cry_12 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_13_LC_6_3_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_13_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_13_LC_6_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_13_LC_6_3_4  (
            .in0(_gnd_net_),
            .in1(N__20741),
            .in2(_gnd_net_),
            .in3(N__20729),
            .lcout(\b2v_inst20.counterZ0Z_13 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_12 ),
            .carryout(\b2v_inst20.counter_1_cry_13 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_14_LC_6_3_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_14_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_14_LC_6_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_14_LC_6_3_5  (
            .in0(_gnd_net_),
            .in1(N__20725),
            .in2(_gnd_net_),
            .in3(N__20711),
            .lcout(\b2v_inst20.counterZ0Z_14 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_13 ),
            .carryout(\b2v_inst20.counter_1_cry_14 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_15_LC_6_3_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_15_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_15_LC_6_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_15_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(N__20708),
            .in2(_gnd_net_),
            .in3(N__20696),
            .lcout(\b2v_inst20.counterZ0Z_15 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_14 ),
            .carryout(\b2v_inst20.counter_1_cry_15 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_16_LC_6_3_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_16_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_16_LC_6_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_16_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(N__20693),
            .in2(_gnd_net_),
            .in3(N__20681),
            .lcout(\b2v_inst20.counterZ0Z_16 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_15 ),
            .carryout(\b2v_inst20.counter_1_cry_16 ),
            .clk(N__36167),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_17_LC_6_4_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_17_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_17_LC_6_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_17_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__20677),
            .in2(_gnd_net_),
            .in3(N__20663),
            .lcout(\b2v_inst20.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\b2v_inst20.counter_1_cry_17 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_18_LC_6_4_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_18_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_18_LC_6_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_18_LC_6_4_1  (
            .in0(_gnd_net_),
            .in1(N__20660),
            .in2(_gnd_net_),
            .in3(N__20648),
            .lcout(\b2v_inst20.counterZ0Z_18 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_17 ),
            .carryout(\b2v_inst20.counter_1_cry_18 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_19_LC_6_4_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_19_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_19_LC_6_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_19_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__20912),
            .in2(_gnd_net_),
            .in3(N__20900),
            .lcout(\b2v_inst20.counterZ0Z_19 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_18 ),
            .carryout(\b2v_inst20.counter_1_cry_19 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_20_LC_6_4_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_20_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_20_LC_6_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_20_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(N__20896),
            .in2(_gnd_net_),
            .in3(N__20882),
            .lcout(\b2v_inst20.counterZ0Z_20 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_19 ),
            .carryout(\b2v_inst20.counter_1_cry_20 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_21_LC_6_4_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_21_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_21_LC_6_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_21_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(N__20879),
            .in2(_gnd_net_),
            .in3(N__20867),
            .lcout(\b2v_inst20.counterZ0Z_21 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_20 ),
            .carryout(\b2v_inst20.counter_1_cry_21 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_22_LC_6_4_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_22_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_22_LC_6_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_22_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(N__20864),
            .in2(_gnd_net_),
            .in3(N__20852),
            .lcout(\b2v_inst20.counterZ0Z_22 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_21 ),
            .carryout(\b2v_inst20.counter_1_cry_22 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_23_LC_6_4_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_23_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_23_LC_6_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_23_LC_6_4_6  (
            .in0(_gnd_net_),
            .in1(N__20849),
            .in2(_gnd_net_),
            .in3(N__20837),
            .lcout(\b2v_inst20.counterZ0Z_23 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_22 ),
            .carryout(\b2v_inst20.counter_1_cry_23 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_24_LC_6_4_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_24_LC_6_4_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_24_LC_6_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_24_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(N__20834),
            .in2(_gnd_net_),
            .in3(N__20822),
            .lcout(\b2v_inst20.counterZ0Z_24 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_23 ),
            .carryout(\b2v_inst20.counter_1_cry_24 ),
            .clk(N__36322),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_25_LC_6_5_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_25_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_25_LC_6_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_25_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__20819),
            .in2(_gnd_net_),
            .in3(N__20807),
            .lcout(\b2v_inst20.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\b2v_inst20.counter_1_cry_25 ),
            .clk(N__36339),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_26_LC_6_5_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_26_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_26_LC_6_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_26_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__20804),
            .in2(_gnd_net_),
            .in3(N__20792),
            .lcout(\b2v_inst20.counterZ0Z_26 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_25 ),
            .carryout(\b2v_inst20.counter_1_cry_26 ),
            .clk(N__36339),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_27_LC_6_5_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_27_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_27_LC_6_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_27_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__21004),
            .in2(_gnd_net_),
            .in3(N__20990),
            .lcout(\b2v_inst20.counterZ0Z_27 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_26 ),
            .carryout(\b2v_inst20.counter_1_cry_27 ),
            .clk(N__36339),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_28_LC_6_5_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_28_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_28_LC_6_5_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst20.counter_28_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20975),
            .in3(N__20987),
            .lcout(\b2v_inst20.counterZ0Z_28 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_27 ),
            .carryout(\b2v_inst20.counter_1_cry_28 ),
            .clk(N__36339),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_29_LC_6_5_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_29_LC_6_5_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_29_LC_6_5_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst20.counter_29_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20963),
            .in3(N__20984),
            .lcout(\b2v_inst20.counterZ0Z_29 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_28 ),
            .carryout(\b2v_inst20.counter_1_cry_29 ),
            .clk(N__36339),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_30_LC_6_5_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_30_LC_6_5_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_30_LC_6_5_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst20.counter_30_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20951),
            .in3(N__20981),
            .lcout(\b2v_inst20.counterZ0Z_30 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_29 ),
            .carryout(\b2v_inst20.counter_1_cry_30 ),
            .clk(N__36339),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_31_LC_6_5_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_31_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_31_LC_6_5_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst20.counter_31_LC_6_5_6  (
            .in0(N__20936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20978),
            .lcout(\b2v_inst20.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36339),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_6_5_7 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_6_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_7_c_RNO_LC_6_5_7  (
            .in0(N__20971),
            .in1(N__20959),
            .in2(N__20950),
            .in3(N__20935),
            .lcout(\b2v_inst20.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_6_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_6_6_0 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_8_LC_6_6_0  (
            .in0(N__22760),
            .in1(N__25450),
            .in2(_gnd_net_),
            .in3(N__23531),
            .lcout(\b2v_inst11.un1_dutycycle_53_9_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIO6J59_8_LC_6_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIO6J59_8_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIO6J59_8_LC_6_6_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIO6J59_8_LC_6_6_1  (
            .in0(N__31221),
            .in1(N__21055),
            .in2(N__22814),
            .in3(N__23587),
            .lcout(\b2v_inst11.dutycycleZ1Z_5 ),
            .ltout(\b2v_inst11.dutycycleZ1Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_6_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_6_6_2 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_3_LC_6_6_2  (
            .in0(N__22761),
            .in1(N__24567),
            .in2(N__20915),
            .in3(N__23422),
            .lcout(\b2v_inst11.un1_dutycycle_53_3_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_8_LC_6_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_8_LC_6_6_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_8_LC_6_6_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.dutycycle_8_LC_6_6_3  (
            .in0(N__22813),
            .in1(N__21056),
            .in2(N__31244),
            .in3(N__23588),
            .lcout(\b2v_inst11.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36437),
            .ce(),
            .sr(N__31032));
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_6_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_6_6_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_3_LC_6_6_4  (
            .in0(N__23435),
            .in1(N__25451),
            .in2(N__22790),
            .in3(N__23532),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_7Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_7_LC_6_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_7_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_7_LC_6_6_5 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_7_LC_6_6_5  (
            .in0(N__21047),
            .in1(N__22914),
            .in2(N__21041),
            .in3(N__29969),
            .lcout(\b2v_inst11.dutycycle_RNI_8Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_6_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_6_6_6 .LUT_INIT=16'b0101011100010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_8_LC_6_6_6  (
            .in0(N__23543),
            .in1(N__24568),
            .in2(N__22791),
            .in3(N__25452),
            .lcout(),
            .ltout(\b2v_inst11.N_26_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_7_LC_6_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_7_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_7_LC_6_6_7 .LUT_INIT=16'b0101111100001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_7_LC_6_6_7  (
            .in0(N__25453),
            .in1(N__22915),
            .in2(N__21038),
            .in3(N__29970),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIGFG69_13_LC_6_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIGFG69_13_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIGFG69_13_LC_6_7_0 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \b2v_inst11.dutycycle_RNIGFG69_13_LC_6_7_0  (
            .in0(N__21025),
            .in1(N__33850),
            .in2(N__24731),
            .in3(N__23017),
            .lcout(\b2v_inst11.dutycycleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_13_LC_6_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_13_LC_6_7_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_13_LC_6_7_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \b2v_inst11.dutycycle_13_LC_6_7_1  (
            .in0(N__23018),
            .in1(N__21026),
            .in2(N__33887),
            .in3(N__24727),
            .lcout(\b2v_inst11.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36198),
            .ce(),
            .sr(N__31039));
    defparam \b2v_inst11.dutycycle_4_LC_6_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_4_LC_6_7_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_4_LC_6_7_2 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \b2v_inst11.dutycycle_4_LC_6_7_2  (
            .in0(N__23198),
            .in1(N__21016),
            .in2(N__22943),
            .in3(N__33854),
            .lcout(\b2v_inst11.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36198),
            .ce(),
            .sr(N__31039));
    defparam \b2v_inst11.dutycycle_RNIGQE59_4_LC_6_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIGQE59_4_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIGQE59_4_LC_6_7_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNIGQE59_4_LC_6_7_3  (
            .in0(N__33849),
            .in1(N__22939),
            .in2(N__21017),
            .in3(N__23197),
            .lcout(\b2v_inst11.dutycycleZ0Z_7 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_6_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_6_7_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_4_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21086),
            .in3(N__22781),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_6_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_6_7_5 .LUT_INIT=16'b1001100111000110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_7_LC_6_7_5  (
            .in0(N__21083),
            .in1(N__21071),
            .in2(N__21077),
            .in3(N__22918),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_6_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_6_7_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_11_LC_6_7_6  (
            .in0(N__25219),
            .in1(_gnd_net_),
            .in2(N__21074),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_6_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_6_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_11_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(N__25218),
            .in2(_gnd_net_),
            .in3(N__23546),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_6_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_6_8_0 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_2_LC_6_8_0  (
            .in0(N__23398),
            .in1(_gnd_net_),
            .in2(N__29971),
            .in3(N__33191),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_LC_6_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_6_8_1 .LUT_INIT=16'b1010010100101101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_LC_6_8_1  (
            .in0(N__31374),
            .in1(N__33707),
            .in2(N__21065),
            .in3(N__24588),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_2_LC_6_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_2_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_2_LC_6_8_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_2_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21062),
            .in3(N__33192),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_6_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_6_8_3 .LUT_INIT=16'b1101001010110100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_7_LC_6_8_3  (
            .in0(N__22917),
            .in1(N__24595),
            .in2(N__23570),
            .in3(N__23401),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_6_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_6_8_4 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_3_LC_6_8_4  (
            .in0(N__23399),
            .in1(N__31375),
            .in2(N__24621),
            .in3(N__29957),
            .lcout(),
            .ltout(\b2v_inst11.un1_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_6_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_6_8_5 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_5_LC_6_8_5  (
            .in0(N__21209),
            .in1(N__21161),
            .in2(N__21059),
            .in3(N__35184),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_6_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_6_8_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_7_LC_6_8_6  (
            .in0(N__23400),
            .in1(_gnd_net_),
            .in2(N__24622),
            .in3(N__22916),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_6_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_6_8_7 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_3_LC_6_8_7  (
            .in0(N__31373),
            .in1(N__29953),
            .in2(_gnd_net_),
            .in3(N__23397),
            .lcout(\b2v_inst11.d_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_6_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_6_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_0_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__30176),
            .in2(N__23423),
            .in3(N__31376),
            .lcout(\b2v_inst11.g0_i_a7_1_2 ),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_6_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_6_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__21203),
            .in2(N__30184),
            .in3(N__21197),
            .lcout(\b2v_inst11.mult1_un138_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_6_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_6_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__33166),
            .in2(N__24491),
            .in3(N__21194),
            .lcout(\b2v_inst11.mult1_un131_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_1 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_6_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_6_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__21191),
            .in2(N__33186),
            .in3(N__21164),
            .lcout(\b2v_inst11.mult1_un124_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_2 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_6_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_6_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__21160),
            .in2(N__21149),
            .in3(N__21119),
            .lcout(\b2v_inst11.mult1_un117_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_3 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_6_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_6_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__21116),
            .in2(N__35198),
            .in3(N__21089),
            .lcout(\b2v_inst11.mult1_un110_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_4 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_6_9_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_6_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(N__35188),
            .in2(N__21506),
            .in3(N__21473),
            .lcout(\b2v_inst11.mult1_un103_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_5 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_6_9_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_6_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(N__22661),
            .in2(N__21470),
            .in3(N__21434),
            .lcout(\b2v_inst11.mult1_un96_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_6 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_6_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_6_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__25220),
            .in2(N__21431),
            .in3(N__21398),
            .lcout(\b2v_inst11.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_6_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_6_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__25087),
            .in2(N__21395),
            .in3(N__21362),
            .lcout(\b2v_inst11.mult1_un82_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_8 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_6_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_6_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__21359),
            .in2(N__24950),
            .in3(N__21329),
            .lcout(\b2v_inst11.mult1_un75_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_9 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_6_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__21326),
            .in2(N__23076),
            .in3(N__21287),
            .lcout(\b2v_inst11.mult1_un68_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_6_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_6_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__24699),
            .in2(N__21284),
            .in3(N__21254),
            .lcout(\b2v_inst11.mult1_un61_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_6_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_6_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__24939),
            .in2(N__21251),
            .in3(N__21212),
            .lcout(\b2v_inst11.mult1_un54_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_6_10_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_6_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__23061),
            .in2(N__21614),
            .in3(N__21587),
            .lcout(\b2v_inst11.mult1_un47_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_6_10_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_6_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(N__23282),
            .in2(N__24711),
            .in3(N__21566),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_6_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_6_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__21512),
            .in2(N__24703),
            .in3(N__21548),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\b2v_inst11.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_6_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_6_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.CO2_THRU_LUT4_0_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21545),
            .lcout(\b2v_inst11.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21695),
            .lcout(\b2v_inst11.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o2_LC_6_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o2_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o2_LC_6_11_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o2_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(N__34621),
            .in2(_gnd_net_),
            .in3(N__34455),
            .lcout(\b2v_inst11.N_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21530),
            .lcout(\b2v_inst11.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_14_LC_6_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_6_11_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_14_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23309),
            .in3(N__23057),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIL6AH3_6_LC_6_12_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIL6AH3_6_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIL6AH3_6_LC_6_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIL6AH3_6_LC_6_12_0  (
            .in0(N__21797),
            .in1(N__26864),
            .in2(_gnd_net_),
            .in3(N__22459),
            .lcout(\b2v_inst5.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_6_LC_6_12_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_6_LC_6_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_6_LC_6_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_6_LC_6_12_1  (
            .in0(N__22460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36403),
            .ce(N__26865),
            .sr(N__27341));
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_6_12_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_6_12_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_6_12_2  (
            .in0(N__21791),
            .in1(N__21773),
            .in2(_gnd_net_),
            .in3(N__34932),
            .lcout(\b2v_inst6.N_192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_12_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_12_5  (
            .in0(N__34620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32873),
            .lcout(\b2v_inst11.N_161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_6_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_6_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_6_12_6  (
            .in0(N__21761),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21740),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__21694),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__21680),
            .in2(N__21904),
            .in3(N__21671),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_2_c ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(N__21900),
            .in2(N__21668),
            .in3(N__21659),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_3_c ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__21656),
            .in2(N__21647),
            .in3(N__21650),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_4_c ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(N__21645),
            .in2(N__21623),
            .in3(N__21914),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_5_c ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_13_5  (
            .in0(N__21827),
            .in1(N__21911),
            .in2(N__21905),
            .in3(N__21887),
            .lcout(\b2v_inst11.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_6_c ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_13_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21884),
            .in3(N__21875),
            .lcout(\b2v_inst11.mult1_un138_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un138_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21872),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__23342),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__21869),
            .in2(N__22045),
            .in3(N__21860),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__22041),
            .in2(N__21857),
            .in3(N__21848),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__21845),
            .in2(N__21835),
            .in3(N__21839),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__21831),
            .in2(N__21809),
            .in3(N__21800),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5  (
            .in0(N__21950),
            .in1(N__22052),
            .in2(N__22046),
            .in3(N__22028),
            .lcout(\b2v_inst11.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22025),
            .in3(N__22016),
            .lcout(\b2v_inst11.mult1_un145_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un145_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22013),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_6_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_6_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__33197),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(N__23333),
            .in2(N__22165),
            .in3(N__22001),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__22161),
            .in2(N__21998),
            .in3(N__21983),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__21980),
            .in2(N__21958),
            .in3(N__21965),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__21954),
            .in2(N__21932),
            .in3(N__21917),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_15_5  (
            .in0(N__22112),
            .in1(N__22172),
            .in2(N__22166),
            .in3(N__22139),
            .lcout(\b2v_inst11.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22136),
            .in3(N__22127),
            .lcout(\b2v_inst11.mult1_un152_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un152_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22094),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIB8QH1_0_1_LC_7_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIB8QH1_0_1_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIB8QH1_0_1_LC_7_1_0 .LUT_INIT=16'b0100000001001100;
    LogicCell40 \b2v_inst36.count_RNIB8QH1_0_1_LC_7_1_0  (
            .in0(N__23897),
            .in1(N__24054),
            .in2(N__29150),
            .in3(N__22061),
            .lcout(\b2v_inst36.un12_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIB8QH1_1_LC_7_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIB8QH1_1_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIB8QH1_1_LC_7_1_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIB8QH1_1_LC_7_1_1  (
            .in0(N__22060),
            .in1(N__29134),
            .in2(_gnd_net_),
            .in3(N__23895),
            .lcout(\b2v_inst36.un2_count_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_7_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_7_1_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_7_1_2  (
            .in0(N__26171),
            .in1(N__24055),
            .in2(N__24038),
            .in3(N__28939),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIDPQG1_11_LC_7_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIDPQG1_11_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIDPQG1_11_LC_7_1_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNIDPQG1_11_LC_7_1_3  (
            .in0(_gnd_net_),
            .in1(N__22067),
            .in2(N__22073),
            .in3(N__29135),
            .lcout(\b2v_inst36.countZ0Z_11 ),
            .ltout(\b2v_inst36.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_11_LC_7_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_11_LC_7_1_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_11_LC_7_1_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst36.count_11_LC_7_1_4  (
            .in0(N__24037),
            .in1(N__26173),
            .in2(N__22070),
            .in3(N__28941),
            .lcout(\b2v_inst36.count_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36001),
            .ce(N__29141),
            .sr(N__28938));
    defparam \b2v_inst36.count_1_LC_7_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_1_LC_7_1_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_1_LC_7_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_1_LC_7_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23896),
            .lcout(\b2v_inst36.count_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36001),
            .ce(N__29141),
            .sr(N__28938));
    defparam \b2v_inst36.count_0_LC_7_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_0_LC_7_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_0_LC_7_1_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst36.count_0_LC_7_1_6  (
            .in0(N__26172),
            .in1(N__22185),
            .in2(_gnd_net_),
            .in3(N__28940),
            .lcout(\b2v_inst36.count_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36001),
            .ce(N__29141),
            .sr(N__28938));
    defparam \b2v_inst36.count_RNI1FG91_0_LC_7_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI1FG91_0_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI1FG91_0_LC_7_1_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst36.count_RNI1FG91_0_LC_7_1_7  (
            .in0(N__22186),
            .in1(N__28937),
            .in2(_gnd_net_),
            .in3(N__26170),
            .lcout(\b2v_inst36.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI6K3V_0_0_LC_7_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI6K3V_0_0_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI6K3V_0_0_LC_7_2_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst36.count_RNI6K3V_0_0_LC_7_2_0  (
            .in0(N__24016),
            .in1(N__23950),
            .in2(N__22190),
            .in3(N__23986),
            .lcout(\b2v_inst36.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIL5VG1_15_LC_7_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIL5VG1_15_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIL5VG1_15_LC_7_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIL5VG1_15_LC_7_2_1  (
            .in0(N__22208),
            .in1(N__29147),
            .in2(_gnd_net_),
            .in3(N__24263),
            .lcout(\b2v_inst36.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_15_LC_7_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_15_LC_7_2_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_15_LC_7_2_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_15_LC_7_2_2  (
            .in0(N__24262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36192),
            .ce(N__29146),
            .sr(N__28981));
    defparam \b2v_inst36.count_RNIHVSG1_13_LC_7_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIHVSG1_13_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIHVSG1_13_LC_7_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIHVSG1_13_LC_7_2_3  (
            .in0(N__22202),
            .in1(N__29108),
            .in2(_gnd_net_),
            .in3(N__24001),
            .lcout(\b2v_inst36.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_13_LC_7_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_13_LC_7_2_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_13_LC_7_2_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_13_LC_7_2_4  (
            .in0(N__24002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36192),
            .ce(N__29146),
            .sr(N__28981));
    defparam \b2v_inst36.count_RNIJ2UG1_14_LC_7_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJ2UG1_14_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJ2UG1_14_LC_7_2_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIJ2UG1_14_LC_7_2_5  (
            .in0(N__22196),
            .in1(N__29109),
            .in2(_gnd_net_),
            .in3(N__23971),
            .lcout(\b2v_inst36.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_14_LC_7_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_14_LC_7_2_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_14_LC_7_2_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_14_LC_7_2_6  (
            .in0(N__23972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36192),
            .ce(N__29146),
            .sr(N__28981));
    defparam \b2v_inst36.count_RNI6K3V_0_LC_7_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI6K3V_0_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI6K3V_0_LC_7_2_7 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \b2v_inst36.count_RNI6K3V_0_LC_7_2_7  (
            .in0(N__23936),
            .in1(N__29110),
            .in2(_gnd_net_),
            .in3(N__23924),
            .lcout(\b2v_inst36.count_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_7_LC_7_3_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_7_LC_7_3_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_7_LC_7_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_7_LC_7_3_0  (
            .in0(N__22433),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(N__26872),
            .sr(N__27343));
    defparam \b2v_inst5.count_RNID0AN3_11_LC_7_3_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNID0AN3_11_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNID0AN3_11_LC_7_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst5.count_RNID0AN3_11_LC_7_3_1  (
            .in0(N__22521),
            .in1(N__22252),
            .in2(_gnd_net_),
            .in3(N__26856),
            .lcout(\b2v_inst5.un2_count_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_11_LC_7_3_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_11_LC_7_3_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_11_LC_7_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_11_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22522),
            .lcout(\b2v_inst5.count_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(N__26872),
            .sr(N__27343));
    defparam \b2v_inst5.count_RNIN9BH3_7_LC_7_3_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIN9BH3_7_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIN9BH3_7_LC_7_3_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIN9BH3_7_LC_7_3_3  (
            .in0(N__22259),
            .in1(N__26855),
            .in2(_gnd_net_),
            .in3(N__22432),
            .lcout(\b2v_inst5.countZ0Z_7 ),
            .ltout(\b2v_inst5.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNID0AN3_0_11_LC_7_3_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNID0AN3_0_11_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNID0AN3_0_11_LC_7_3_4 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \b2v_inst5.count_RNID0AN3_0_11_LC_7_3_4  (
            .in0(N__22253),
            .in1(N__26873),
            .in2(N__22244),
            .in3(N__22523),
            .lcout(\b2v_inst5.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIF3BN3_12_LC_7_3_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIF3BN3_12_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIF3BN3_12_LC_7_3_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \b2v_inst5.count_RNIF3BN3_12_LC_7_3_5  (
            .in0(N__22241),
            .in1(N__22504),
            .in2(N__27342),
            .in3(N__26857),
            .lcout(\b2v_inst5.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_12_LC_7_3_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_12_LC_7_3_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_12_LC_7_3_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst5.count_12_LC_7_3_6  (
            .in0(N__22505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27335),
            .lcout(\b2v_inst5.count_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(N__26872),
            .sr(N__27343));
    defparam \b2v_inst5.count_14_LC_7_3_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_14_LC_7_3_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_14_LC_7_3_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst5.count_14_LC_7_3_7  (
            .in0(_gnd_net_),
            .in1(N__24332),
            .in2(_gnd_net_),
            .in3(N__27344),
            .lcout(\b2v_inst5.count_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(N__26872),
            .sr(N__27343));
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_7_4_0 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_7_4_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_RNO_LC_7_4_0  (
            .in0(N__22235),
            .in1(N__22305),
            .in2(N__22399),
            .in3(N__22371),
            .lcout(\b2v_inst20.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_6_LC_7_4_1 .C_ON=1'b0;
    defparam \b2v_inst20.counter_6_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_6_LC_7_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst20.counter_6_LC_7_4_1  (
            .in0(N__24190),
            .in1(N__22409),
            .in2(_gnd_net_),
            .in3(N__22395),
            .lcout(\b2v_inst20.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36194),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_0_LC_7_4_2 .C_ON=1'b0;
    defparam \b2v_inst20.counter_0_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_0_LC_7_4_2 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \b2v_inst20.counter_0_LC_7_4_2  (
            .in0(N__22351),
            .in1(N__24192),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst20.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36194),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_LC_7_4_3 .C_ON=1'b0;
    defparam \b2v_inst20.counter_1_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_1_LC_7_4_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst20.counter_1_LC_7_4_3  (
            .in0(N__24191),
            .in1(_gnd_net_),
            .in2(N__22378),
            .in3(N__22350),
            .lcout(\b2v_inst20.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36194),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_7_4_4 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_7_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_RNO_LC_7_4_4  (
            .in0(N__22349),
            .in1(N__24228),
            .in2(N__22282),
            .in3(N__24120),
            .lcout(\b2v_inst20.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_5_LC_7_4_5 .C_ON=1'b0;
    defparam \b2v_inst20.counter_5_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_5_LC_7_4_5 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \b2v_inst20.counter_5_LC_7_4_5  (
            .in0(N__22306),
            .in1(_gnd_net_),
            .in2(N__24194),
            .in3(N__22322),
            .lcout(\b2v_inst20.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36194),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_4_LC_7_4_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_4_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_4_LC_7_4_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_4_LC_7_4_6  (
            .in0(N__22278),
            .in1(N__22292),
            .in2(_gnd_net_),
            .in3(N__24193),
            .lcout(\b2v_inst20.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36194),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_7_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_7_4_7 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_7_4_7  (
            .in0(N__27463),
            .in1(N__27044),
            .in2(N__27071),
            .in3(N__27532),
            .lcout(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_0_c_LC_7_5_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_0_c_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_0_c_LC_7_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_0_c_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24341),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNIKSVJ1_LC_7_5_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNIKSVJ1_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNIKSVJ1_LC_7_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_0_c_RNIKSVJ1_LC_7_5_1  (
            .in0(N__27307),
            .in1(N__26519),
            .in2(_gnd_net_),
            .in3(N__22262),
            .lcout(\b2v_inst5.count_rst_13 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_0 ),
            .carryout(\b2v_inst5.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNILU0K1_LC_7_5_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNILU0K1_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNILU0K1_LC_7_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_1_c_RNILU0K1_LC_7_5_2  (
            .in0(N__27305),
            .in1(N__26498),
            .in2(_gnd_net_),
            .in3(N__22472),
            .lcout(\b2v_inst5.count_rst_12 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_1 ),
            .carryout(\b2v_inst5.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNIM02K1_LC_7_5_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNIM02K1_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNIM02K1_LC_7_5_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_2_c_RNIM02K1_LC_7_5_3  (
            .in0(N__27309),
            .in1(_gnd_net_),
            .in2(N__26555),
            .in3(N__22469),
            .lcout(\b2v_inst5.count_rst_11 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_2 ),
            .carryout(\b2v_inst5.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_7_5_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_7_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__24437),
            .in2(_gnd_net_),
            .in3(N__22466),
            .lcout(\b2v_inst5.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_3 ),
            .carryout(\b2v_inst5.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIO44K1_LC_7_5_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIO44K1_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIO44K1_LC_7_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_4_c_RNIO44K1_LC_7_5_5  (
            .in0(N__27308),
            .in1(N__26429),
            .in2(_gnd_net_),
            .in3(N__22463),
            .lcout(\b2v_inst5.count_rst_9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_4 ),
            .carryout(\b2v_inst5.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIP65K1_LC_7_5_6 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIP65K1_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIP65K1_LC_7_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_5_c_RNIP65K1_LC_7_5_6  (
            .in0(N__27304),
            .in1(N__26398),
            .in2(_gnd_net_),
            .in3(N__22445),
            .lcout(\b2v_inst5.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_5 ),
            .carryout(\b2v_inst5.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIQ86K1_LC_7_5_7 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIQ86K1_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIQ86K1_LC_7_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_6_c_RNIQ86K1_LC_7_5_7  (
            .in0(N__27306),
            .in1(N__22442),
            .in2(_gnd_net_),
            .in3(N__22421),
            .lcout(\b2v_inst5.count_rst_7 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_6 ),
            .carryout(\b2v_inst5.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_7_6_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_7_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__24472),
            .in2(_gnd_net_),
            .in3(N__22418),
            .lcout(\b2v_inst5.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_7_6_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_7_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__27023),
            .in2(_gnd_net_),
            .in3(N__22415),
            .lcout(\b2v_inst5.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_8 ),
            .carryout(\b2v_inst5.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_7_6_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_7_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__26651),
            .in2(_gnd_net_),
            .in3(N__22412),
            .lcout(\b2v_inst5.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_9 ),
            .carryout(\b2v_inst5.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_7_6_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_7_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_7_6_3  (
            .in0(N__27313),
            .in1(N__22535),
            .in2(_gnd_net_),
            .in3(N__22508),
            .lcout(\b2v_inst5.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_10 ),
            .carryout(\b2v_inst5.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_7_6_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_7_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__24289),
            .in2(_gnd_net_),
            .in3(N__22493),
            .lcout(\b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_11 ),
            .carryout(\b2v_inst5.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_7_6_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_7_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__26535),
            .in2(_gnd_net_),
            .in3(N__22490),
            .lcout(\b2v_inst5.un2_count_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_12 ),
            .carryout(\b2v_inst5.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_7_6_6 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_7_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__24308),
            .in2(_gnd_net_),
            .in3(N__22487),
            .lcout(\b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_13 ),
            .carryout(\b2v_inst5.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_7_6_7 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_7_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_7_6_7  (
            .in0(N__27314),
            .in1(N__26615),
            .in2(_gnd_net_),
            .in3(N__22484),
            .lcout(\b2v_inst5.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_LC_7_7_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_LC_7_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_c_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30175),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_7_7_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_7_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__31350),
            .in2(N__27141),
            .in3(N__22481),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_7_7_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_7_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__27130),
            .in2(N__33196),
            .in3(N__22478),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_7_7_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_7_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__27135),
            .in2(N__23425),
            .in3(N__22475),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_2 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_7_7_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_7_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__27131),
            .in2(N__24596),
            .in3(N__22928),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_3 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_7_7_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_7_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__35183),
            .in2(N__27142),
            .in3(N__22925),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_4 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_7_7_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_7_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__29906),
            .in2(N__27143),
            .in3(N__22922),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_7_7_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_7_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__27139),
            .in2(N__22919),
            .in3(N__22817),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9J1_LC_7_8_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9J1_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9J1_LC_7_8_0 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9J1_LC_7_8_0  (
            .in0(N__33842),
            .in1(N__27118),
            .in2(N__23568),
            .in3(N__22799),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_7_c_RNIUJ9JZ0Z1 ),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJ1_LC_7_8_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJ1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJ1_LC_7_8_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJ1_LC_7_8_1  (
            .in0(N__33881),
            .in1(N__27121),
            .in2(N__22796),
            .in3(N__22670),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_8_c_RNIVLAJZ0Z1 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJ1_LC_7_8_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJ1_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJ1_LC_7_8_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJ1_LC_7_8_2  (
            .in0(N__33843),
            .in1(N__27119),
            .in2(N__22667),
            .in3(N__22541),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_9_c_RNI0OBJZ0Z1 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_9 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUF1_LC_7_8_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUF1_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUF1_LC_7_8_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUF1_LC_7_8_3  (
            .in0(N__33882),
            .in1(N__27122),
            .in2(N__25196),
            .in3(N__22538),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_10_c_RNI8IUFZ0Z1 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_10 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_11_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNI9KVF1_LC_7_8_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNI9KVF1_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNI9KVF1_LC_7_8_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_11_c_RNI9KVF1_LC_7_8_4  (
            .in0(N__33844),
            .in1(N__25037),
            .in2(N__27140),
            .in3(N__23021),
            .lcout(\b2v_inst11.dutycycle_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_11_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_12_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_7_8_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_7_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__27126),
            .in2(N__24935),
            .in3(N__23009),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_12_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_13_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_7_8_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_7_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__27120),
            .in2(N__23086),
            .in3(N__23006),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_13_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_7_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_7_8_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_7_8_7  (
            .in0(N__24704),
            .in1(N__33411),
            .in2(_gnd_net_),
            .in3(N__23003),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIANKU4_3_LC_7_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIANKU4_3_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIANKU4_3_LC_7_9_0 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \b2v_inst11.dutycycle_RNIANKU4_3_LC_7_9_0  (
            .in0(N__34289),
            .in1(N__25301),
            .in2(N__22994),
            .in3(N__23449),
            .lcout(\b2v_inst11.un1_clk_100khz_43_and_i_0_0_0 ),
            .ltout(\b2v_inst11.un1_clk_100khz_43_and_i_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI61IA9_3_LC_7_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI61IA9_3_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI61IA9_3_LC_7_9_1 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI61IA9_3_LC_7_9_1  (
            .in0(N__34799),
            .in1(N__22976),
            .in2(N__23000),
            .in3(N__22956),
            .lcout(\b2v_inst11.dutycycleZ0Z_3 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_7_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_7_9_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_3_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22997),
            .in3(N__25246),
            .lcout(\b2v_inst11.un1_clk_100khz_43_and_i_0_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI52KD2_3_LC_7_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI52KD2_3_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI52KD2_3_LC_7_9_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI52KD2_3_LC_7_9_3  (
            .in0(N__22985),
            .in1(N__33848),
            .in2(N__22961),
            .in3(N__31193),
            .lcout(\b2v_inst11.dutycycle_e_1_3 ),
            .ltout(\b2v_inst11.dutycycle_e_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_3_LC_7_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_3_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_3_LC_7_9_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \b2v_inst11.dutycycle_3_LC_7_9_4  (
            .in0(N__22957),
            .in1(N__22970),
            .in2(N__22964),
            .in3(N__34800),
            .lcout(\b2v_inst11.dutycycle_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36099),
            .ce(),
            .sr(N__31038));
    defparam \b2v_inst11.dutycycle_RNITSFK3_4_LC_7_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITSFK3_4_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITSFK3_4_LC_7_9_5 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNITSFK3_4_LC_7_9_5  (
            .in0(N__25302),
            .in1(N__34290),
            .in2(N__25250),
            .in3(N__24623),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_40_and_i_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIT35D7_4_LC_7_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIT35D7_4_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIT35D7_4_LC_7_9_6 .LUT_INIT=16'b1010101010100010;
    LogicCell40 \b2v_inst11.dutycycle_RNIT35D7_4_LC_7_9_6  (
            .in0(N__31192),
            .in1(N__34798),
            .in2(N__23201),
            .in3(N__23450),
            .lcout(\b2v_inst11.dutycycle_RNIT35D7Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIKLI69_15_LC_7_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIKLI69_15_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIKLI69_15_LC_7_10_0 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \b2v_inst11.dutycycle_RNIKLI69_15_LC_7_10_0  (
            .in0(N__23140),
            .in1(N__33846),
            .in2(N__23165),
            .in3(N__23155),
            .lcout(\b2v_inst11.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIT35D7_14_LC_7_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIT35D7_14_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIT35D7_14_LC_7_10_1 .LUT_INIT=16'b0010001010100010;
    LogicCell40 \b2v_inst11.dutycycle_RNIT35D7_14_LC_7_10_1  (
            .in0(N__31194),
            .in1(N__34804),
            .in2(N__23186),
            .in3(N__27643),
            .lcout(\b2v_inst11.dutycycle_en_11 ),
            .ltout(\b2v_inst11.dutycycle_en_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_14_LC_7_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_14_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_14_LC_7_10_2 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \b2v_inst11.dutycycle_14_LC_7_10_2  (
            .in0(N__23129),
            .in1(N__33847),
            .in2(N__23171),
            .in3(N__23111),
            .lcout(\b2v_inst11.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36394),
            .ce(),
            .sr(N__31021));
    defparam \b2v_inst11.dutycycle_RNIANKU4_15_LC_7_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIANKU4_15_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIANKU4_15_LC_7_10_3 .LUT_INIT=16'b1110111111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIANKU4_15_LC_7_10_3  (
            .in0(N__25320),
            .in1(N__24987),
            .in2(N__34285),
            .in3(N__24688),
            .lcout(),
            .ltout(\b2v_inst11.N_158_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIT35D7_15_LC_7_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIT35D7_15_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIT35D7_15_LC_7_10_4 .LUT_INIT=16'b0100000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIT35D7_15_LC_7_10_4  (
            .in0(N__27644),
            .in1(N__31195),
            .in2(N__23168),
            .in3(N__34805),
            .lcout(\b2v_inst11.dutycycle_RNIT35D7Z0Z_15 ),
            .ltout(\b2v_inst11.dutycycle_RNIT35D7Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_15_LC_7_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_15_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_15_LC_7_10_5 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \b2v_inst11.dutycycle_15_LC_7_10_5  (
            .in0(N__23156),
            .in1(N__33917),
            .in2(N__23144),
            .in3(N__23141),
            .lcout(\b2v_inst11.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36394),
            .ce(),
            .sr(N__31021));
    defparam \b2v_inst11.dutycycle_RNIIIH69_14_LC_7_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIIIH69_14_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIIIH69_14_LC_7_10_6 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \b2v_inst11.dutycycle_RNIIIH69_14_LC_7_10_6  (
            .in0(N__23128),
            .in1(N__33845),
            .in2(N__23120),
            .in3(N__23110),
            .lcout(\b2v_inst11.dutycycleZ0Z_12 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_7_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_7_10_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_14_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__24689),
            .in2(N__23312),
            .in3(N__23305),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIM50S4_LC_7_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIM50S4_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIM50S4_LC_7_11_0 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIM50S4_LC_7_11_0  (
            .in0(N__23273),
            .in1(N__34807),
            .in2(N__23261),
            .in3(N__33929),
            .lcout(\b2v_inst11.dutycycle_set_1 ),
            .ltout(\b2v_inst11.dutycycle_set_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_5_LC_7_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_5_LC_7_11_1 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_5_LC_7_11_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_5_LC_7_11_1  (
            .in0(N__23219),
            .in1(N__31191),
            .in2(N__23264),
            .in3(N__34643),
            .lcout(\b2v_inst11.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36315),
            .ce(),
            .sr(N__31020));
    defparam \b2v_inst11.func_state_RNISPKF1_0_1_LC_7_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNISPKF1_0_1_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNISPKF1_0_1_LC_7_11_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.func_state_RNISPKF1_0_1_LC_7_11_2  (
            .in0(N__29638),
            .in1(N__33415),
            .in2(N__34287),
            .in3(N__30276),
            .lcout(\b2v_inst11.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIBGDMD_6_LC_7_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIBGDMD_6_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIBGDMD_6_LC_7_11_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIBGDMD_6_LC_7_11_3  (
            .in0(N__23237),
            .in1(N__23227),
            .in2(N__23606),
            .in3(N__31190),
            .lcout(\b2v_inst11.dutycycleZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNISPKF1_1_LC_7_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNISPKF1_1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNISPKF1_1_LC_7_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.func_state_RNISPKF1_1_LC_7_11_4  (
            .in0(N__29639),
            .in1(N__33416),
            .in2(N__34288),
            .in3(N__30277),
            .lcout(),
            .ltout(\b2v_inst11.N_300_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIN71S4_LC_7_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIN71S4_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIN71S4_LC_7_11_5 .LUT_INIT=16'b1111011111110011;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIN71S4_LC_7_11_5  (
            .in0(N__33928),
            .in1(N__34806),
            .in2(N__23252),
            .in3(N__23249),
            .lcout(\b2v_inst11.dutycycle_set_0_0 ),
            .ltout(\b2v_inst11.dutycycle_set_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_6_LC_7_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_6_LC_7_11_6 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_6_LC_7_11_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_6_LC_7_11_6  (
            .in0(N__23228),
            .in1(N__31249),
            .in2(N__23231),
            .in3(N__23605),
            .lcout(\b2v_inst11.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36315),
            .ce(),
            .sr(N__31020));
    defparam \b2v_inst11.dutycycle_RNIFNB2O_5_LC_7_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIFNB2O_5_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIFNB2O_5_LC_7_11_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIFNB2O_5_LC_7_11_7  (
            .in0(N__23218),
            .in1(N__31189),
            .in2(N__23210),
            .in3(N__34642),
            .lcout(\b2v_inst11.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5DSV7_6_LC_7_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5DSV7_6_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5DSV7_6_LC_7_12_0 .LUT_INIT=16'b0000011111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI5DSV7_6_LC_7_12_0  (
            .in0(N__23321),
            .in1(N__24866),
            .in2(N__25259),
            .in3(N__34796),
            .lcout(\b2v_inst11.dutycycle_eena_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_6_LC_7_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_6_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_6_LC_7_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_6_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33049),
            .lcout(\b2v_inst11.N_200_i ),
            .ltout(\b2v_inst11.N_200_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_7_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_7_12_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_7_12_2  (
            .in0(N__33886),
            .in1(_gnd_net_),
            .in2(N__23594),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNIDQ4A1_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI9LPN6_8_LC_7_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI9LPN6_8_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI9LPN6_8_LC_7_12_3 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \b2v_inst11.dutycycle_RNI9LPN6_8_LC_7_12_3  (
            .in0(N__34797),
            .in1(N__23456),
            .in2(N__23591),
            .in3(N__25240),
            .lcout(\b2v_inst11.dutycycle_eena_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNITSFK3_8_LC_7_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITSFK3_8_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITSFK3_8_LC_7_12_4 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNITSFK3_8_LC_7_12_4  (
            .in0(N__25239),
            .in1(N__25316),
            .in2(N__34311),
            .in3(N__23569),
            .lcout(\b2v_inst11.un1_clk_100khz_32_and_i_0_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_7_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_7_12_5 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__33885),
            .in2(N__33279),
            .in3(N__25238),
            .lcout(\b2v_inst11.un1_clk_100khz_40_and_i_0_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_7_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_7_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_3_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__23424),
            .in2(_gnd_net_),
            .in3(N__30154),
            .lcout(\b2v_inst11.mult1_un145_sum ),
            .ltout(\b2v_inst11.mult1_un145_sum_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23336),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIGUKJ1_1_LC_7_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIGUKJ1_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIGUKJ1_1_LC_7_13_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \b2v_inst11.func_state_RNIGUKJ1_1_LC_7_13_4  (
            .in0(N__34457),
            .in1(N__30275),
            .in2(N__34312),
            .in3(N__33417),
            .lcout(\b2v_inst11.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_7_LC_7_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_7_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_7_LC_7_14_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst11.count_clk_RNI_7_LC_7_14_0  (
            .in0(N__28422),
            .in1(N__23615),
            .in2(_gnd_net_),
            .in3(N__23663),
            .lcout(\b2v_inst11.N_428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_8_LC_7_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_8_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_8_LC_7_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_8_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25717),
            .lcout(\b2v_inst11.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36479),
            .ce(N__28570),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI342J_8_LC_7_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI342J_8_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI342J_8_LC_7_14_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \b2v_inst11.count_clk_RNI342J_8_LC_7_14_2  (
            .in0(N__30637),
            .in1(N__28489),
            .in2(N__25721),
            .in3(N__23630),
            .lcout(\b2v_inst11.count_clkZ0Z_8 ),
            .ltout(\b2v_inst11.count_clkZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_2_LC_7_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_2_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_2_LC_7_14_3 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \b2v_inst11.count_clk_RNI_2_LC_7_14_3  (
            .in0(N__25831),
            .in1(N__25868),
            .in2(N__23624),
            .in3(N__25655),
            .lcout(),
            .ltout(\b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_6_LC_7_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_6_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_6_LC_7_14_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \b2v_inst11.count_clk_RNI_6_LC_7_14_4  (
            .in0(N__25765),
            .in1(N__28424),
            .in2(N__23621),
            .in3(N__23662),
            .lcout(\b2v_inst11.count_clk_RNIZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_3_LC_7_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_3_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_3_LC_7_14_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst11.count_clk_RNI_3_LC_7_14_5  (
            .in0(N__25863),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25732),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_7_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_7_14_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_2_LC_7_14_6  (
            .in0(N__25764),
            .in1(N__25653),
            .in2(N__23618),
            .in3(N__25830),
            .lcout(\b2v_inst11.N_379 ),
            .ltout(\b2v_inst11.N_379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_7_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_7_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_1_LC_7_14_7  (
            .in0(N__28214),
            .in1(N__28423),
            .in2(N__23609),
            .in3(N__23645),
            .lcout(\b2v_inst11.count_clk_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_9_LC_7_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_9_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_9_LC_7_15_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_9_LC_7_15_0  (
            .in0(N__25694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36481),
            .ce(N__28541),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI573J_9_LC_7_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI573J_9_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI573J_9_LC_7_15_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \b2v_inst11.count_clk_RNI573J_9_LC_7_15_1  (
            .in0(N__30635),
            .in1(N__28542),
            .in2(N__23675),
            .in3(N__25693),
            .lcout(\b2v_inst11.count_clkZ0Z_9 ),
            .ltout(\b2v_inst11.count_clkZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_1_LC_7_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_1_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_1_LC_7_15_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \b2v_inst11.count_clk_RNI_1_LC_7_15_2  (
            .in0(N__23723),
            .in1(N__25801),
            .in2(N__23666),
            .in3(N__28215),
            .lcout(\b2v_inst11.N_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_5_LC_7_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_5_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_5_LC_7_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_5_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25783),
            .lcout(\b2v_inst11.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36481),
            .ce(N__28541),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNITQUI_5_LC_7_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNITQUI_5_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNITQUI_5_LC_7_15_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst11.count_clk_RNITQUI_5_LC_7_15_4  (
            .in0(N__28539),
            .in1(N__23654),
            .in2(N__25787),
            .in3(N__30636),
            .lcout(\b2v_inst11.count_clkZ0Z_5 ),
            .ltout(\b2v_inst11.count_clkZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_5_LC_7_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_5_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_5_LC_7_15_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \b2v_inst11.count_clk_RNI_5_LC_7_15_5  (
            .in0(N__25705),
            .in1(_gnd_net_),
            .in2(N__23648),
            .in3(N__23722),
            .lcout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIQA5D_1_LC_7_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIQA5D_1_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIQA5D_1_LC_7_15_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \b2v_inst11.count_clk_RNIQA5D_1_LC_7_15_6  (
            .in0(N__28540),
            .in1(N__23636),
            .in2(N__30706),
            .in3(N__28190),
            .lcout(\b2v_inst11.count_clkZ0Z_1 ),
            .ltout(\b2v_inst11.count_clkZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_1_LC_7_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_1_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_1_LC_7_15_7 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \b2v_inst11.count_clk_1_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__28110),
            .in2(N__23639),
            .in3(N__28173),
            .lcout(\b2v_inst11.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36481),
            .ce(N__28541),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_11_LC_7_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_11_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_11_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_11_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25882),
            .lcout(\b2v_inst11.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36485),
            .ce(N__28568),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_14_LC_7_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_14_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_14_LC_7_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_14_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25918),
            .lcout(\b2v_inst11.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36485),
            .ce(N__28568),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVFGI_15_LC_7_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVFGI_15_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVFGI_15_LC_7_16_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \b2v_inst11.count_clk_RNIVFGI_15_LC_7_16_3  (
            .in0(N__28571),
            .in1(N__30634),
            .in2(N__23708),
            .in3(N__25897),
            .lcout(\b2v_inst11.count_clkZ0Z_15 ),
            .ltout(\b2v_inst11.count_clkZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_15_LC_7_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_15_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_15_LC_7_16_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNI_15_LC_7_16_4  (
            .in0(N__25930),
            .in1(N__28325),
            .in2(N__23726),
            .in3(N__28177),
            .lcout(\b2v_inst11.N_175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNITCFI_14_LC_7_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNITCFI_14_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNITCFI_14_LC_7_16_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.count_clk_RNITCFI_14_LC_7_16_5  (
            .in0(N__25919),
            .in1(N__23714),
            .in2(N__30727),
            .in3(N__28569),
            .lcout(\b2v_inst11.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_15_LC_7_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_15_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_15_LC_7_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_15_LC_7_16_6  (
            .in0(N__25898),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36485),
            .ce(N__28568),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIFESH1_3_LC_8_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIFESH1_3_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIFESH1_3_LC_8_1_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIFESH1_3_LC_8_1_0  (
            .in0(N__23686),
            .in1(N__29117),
            .in2(_gnd_net_),
            .in3(N__23696),
            .lcout(\b2v_inst36.un2_count_1_axb_3 ),
            .ltout(\b2v_inst36.un2_count_1_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_8_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_8_1_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_8_1_1  (
            .in0(N__26142),
            .in1(N__23827),
            .in2(N__23699),
            .in3(N__28916),
            .lcout(\b2v_inst36.count_rst_11 ),
            .ltout(\b2v_inst36.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIFESH1_0_3_LC_8_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIFESH1_0_3_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIFESH1_0_3_LC_8_1_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \b2v_inst36.count_RNIFESH1_0_3_LC_8_1_2  (
            .in0(N__23687),
            .in1(N__29118),
            .in2(N__23690),
            .in3(N__23877),
            .lcout(\b2v_inst36.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_3_LC_8_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_3_LC_8_1_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_3_LC_8_1_3 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.count_3_LC_8_1_3  (
            .in0(N__26143),
            .in1(N__23828),
            .in2(N__23846),
            .in3(N__28960),
            .lcout(\b2v_inst36.count_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__29145),
            .sr(N__28959));
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_8_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_8_1_4 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_8_1_4  (
            .in0(N__23860),
            .in1(N__28914),
            .in2(N__26174),
            .in3(N__23878),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIDBRH1_2_LC_8_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIDBRH1_2_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIDBRH1_2_LC_8_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNIDBRH1_2_LC_8_1_5  (
            .in0(N__29116),
            .in1(_gnd_net_),
            .in2(N__23678),
            .in3(N__23762),
            .lcout(\b2v_inst36.countZ0Z_2 ),
            .ltout(\b2v_inst36.countZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_2_LC_8_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_2_LC_8_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_2_LC_8_1_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst36.count_2_LC_8_1_6  (
            .in0(N__23861),
            .in1(N__28915),
            .in2(N__23765),
            .in3(N__26145),
            .lcout(\b2v_inst36.count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__29145),
            .sr(N__28959));
    defparam \b2v_inst36.count_5_LC_8_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_5_LC_8_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_5_LC_8_1_7 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.count_5_LC_8_1_7  (
            .in0(N__26144),
            .in1(N__23786),
            .in2(N__23809),
            .in3(N__28961),
            .lcout(\b2v_inst36.count_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__29145),
            .sr(N__28959));
    defparam \b2v_inst36.count_7_LC_8_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_7_LC_8_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_7_LC_8_2_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst36.count_7_LC_8_2_0  (
            .in0(N__24082),
            .in1(N__28920),
            .in2(N__24104),
            .in3(N__26153),
            .lcout(\b2v_inst36.count_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36263),
            .ce(N__29096),
            .sr(N__28980));
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_8_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_8_2_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_8_2_1  (
            .in0(N__28918),
            .in1(N__24103),
            .in2(N__24086),
            .in3(N__26147),
            .lcout(\b2v_inst36.count_rst_7 ),
            .ltout(\b2v_inst36.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNINQ0I1_7_LC_8_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNINQ0I1_7_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNINQ0I1_7_LC_8_2_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNINQ0I1_7_LC_8_2_2  (
            .in0(N__29095),
            .in1(_gnd_net_),
            .in2(N__23756),
            .in3(N__23743),
            .lcout(\b2v_inst36.un2_count_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_8_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_8_2_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_8_2_3  (
            .in0(N__23782),
            .in1(N__28917),
            .in2(N__23810),
            .in3(N__26146),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIJKUH1_5_LC_8_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJKUH1_5_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJKUH1_5_LC_8_2_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNIJKUH1_5_LC_8_2_4  (
            .in0(N__29094),
            .in1(_gnd_net_),
            .in2(N__23753),
            .in3(N__23750),
            .lcout(\b2v_inst36.countZ0Z_5 ),
            .ltout(\b2v_inst36.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNINQ0I1_0_7_LC_8_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNINQ0I1_0_7_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNINQ0I1_0_7_LC_8_2_5 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \b2v_inst36.count_RNINQ0I1_0_7_LC_8_2_5  (
            .in0(N__23744),
            .in1(N__23735),
            .in2(N__23729),
            .in3(N__29097),
            .lcout(\b2v_inst36.un12_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_8_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_8_2_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_8_2_6  (
            .in0(N__26148),
            .in1(N__25999),
            .in2(N__25970),
            .in3(N__28919),
            .lcout(\b2v_inst36.count_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_0_c_RNO_LC_8_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_0_c_RNO_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_0_c_RNO_LC_8_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.un2_count_1_cry_0_c_RNO_LC_8_2_7  (
            .in0(N__23935),
            .in1(N__29093),
            .in2(_gnd_net_),
            .in3(N__23923),
            .lcout(\b2v_inst36.un2_count_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_0_c_LC_8_3_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_0_c_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_0_c_LC_8_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_0_c_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__23912),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_0_c_RNI4JMI_LC_8_3_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_0_c_RNI4JMI_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_0_c_RNI4JMI_LC_8_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_0_c_RNI4JMI_LC_8_3_1  (
            .in0(N__28945),
            .in1(N__23906),
            .in2(_gnd_net_),
            .in3(N__23882),
            .lcout(\b2v_inst36.count_rst_13 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_0 ),
            .carryout(\b2v_inst36.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_8_3_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_8_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__23879),
            .in2(_gnd_net_),
            .in3(N__23849),
            .lcout(\b2v_inst36.un2_count_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_1 ),
            .carryout(\b2v_inst36.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_8_3_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_8_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__23845),
            .in2(_gnd_net_),
            .in3(N__23816),
            .lcout(\b2v_inst36.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_2 ),
            .carryout(\b2v_inst36.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_8_3_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_8_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_8_3_4  (
            .in0(N__28973),
            .in1(N__26045),
            .in2(_gnd_net_),
            .in3(N__23813),
            .lcout(\b2v_inst36.count_rst_10 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_3 ),
            .carryout(\b2v_inst36.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_8_3_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_8_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(N__23802),
            .in2(_gnd_net_),
            .in3(N__23771),
            .lcout(\b2v_inst36.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_4 ),
            .carryout(\b2v_inst36.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNILNVH1_LC_8_3_6 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNILNVH1_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNILNVH1_LC_8_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_5_c_RNILNVH1_LC_8_3_6  (
            .in0(N__28974),
            .in1(N__26066),
            .in2(_gnd_net_),
            .in3(N__23768),
            .lcout(\b2v_inst36.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_5 ),
            .carryout(\b2v_inst36.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_8_3_7 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_8_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__24099),
            .in2(_gnd_net_),
            .in3(N__24068),
            .lcout(\b2v_inst36.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_6 ),
            .carryout(\b2v_inst36.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_8_4_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_8_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25969),
            .in3(N__24065),
            .lcout(\b2v_inst36.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_8_4_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_8_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_8_4_1  (
            .in0(N__28964),
            .in1(N__29188),
            .in2(_gnd_net_),
            .in3(N__24062),
            .lcout(\b2v_inst36.count_rst_5 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_8 ),
            .carryout(\b2v_inst36.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_8_4_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_8_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__26204),
            .in2(_gnd_net_),
            .in3(N__24059),
            .lcout(\b2v_inst36.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_9 ),
            .carryout(\b2v_inst36.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_8_4_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_8_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(N__24056),
            .in2(_gnd_net_),
            .in3(N__24023),
            .lcout(\b2v_inst36.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_10 ),
            .carryout(\b2v_inst36.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIFSRG1_LC_8_4_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIFSRG1_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIFSRG1_LC_8_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_11_c_RNIFSRG1_LC_8_4_4  (
            .in0(N__28975),
            .in1(N__26336),
            .in2(_gnd_net_),
            .in3(N__24020),
            .lcout(\b2v_inst36.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_11 ),
            .carryout(\b2v_inst36.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_8_4_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_8_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_8_4_5  (
            .in0(N__28963),
            .in1(N__24017),
            .in2(_gnd_net_),
            .in3(N__23990),
            .lcout(\b2v_inst36.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_12 ),
            .carryout(\b2v_inst36.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_8_4_6 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_8_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_8_4_6  (
            .in0(N__28976),
            .in1(N__23987),
            .in2(_gnd_net_),
            .in3(N__23957),
            .lcout(\b2v_inst36.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_13 ),
            .carryout(\b2v_inst36.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_8_4_7 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_8_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_8_4_7  (
            .in0(N__28965),
            .in1(N__23954),
            .in2(_gnd_net_),
            .in3(N__23939),
            .lcout(\b2v_inst36.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_LC_8_5_0 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_LC_8_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.tmp_1_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__24173),
            .in2(_gnd_net_),
            .in3(N__30509),
            .lcout(SYNTHESIZED_WIRE_1keep_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_2_LC_8_5_1 .C_ON=1'b0;
    defparam \b2v_inst20.counter_2_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_2_LC_8_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst20.counter_2_LC_8_5_1  (
            .in0(N__24171),
            .in1(N__24251),
            .in2(_gnd_net_),
            .in3(N__24238),
            .lcout(\b2v_inst20.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_fast_LC_8_5_2 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_fast_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_fast_LC_8_5_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.tmp_1_fast_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__27045),
            .in2(_gnd_net_),
            .in3(N__24174),
            .lcout(SYNTHESIZED_WIRE_1keep_3_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_rep1_LC_8_5_3 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_rep1_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_rep1_LC_8_5_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst20.tmp_1_rep1_LC_8_5_3  (
            .in0(N__29608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24175),
            .lcout(SYNTHESIZED_WIRE_1keep_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.G_146_LC_8_5_4 .C_ON=1'b0;
    defparam \b2v_inst36.G_146_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.G_146_LC_8_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst36.G_146_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__29607),
            .in2(_gnd_net_),
            .in3(N__24170),
            .lcout(G_146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI3E27_0_LC_8_5_5 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI3E27_0_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI3E27_0_LC_8_5_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst36.curr_state_RNI3E27_0_LC_8_5_5  (
            .in0(N__29294),
            .in1(N__29242),
            .in2(_gnd_net_),
            .in3(N__29342),
            .lcout(),
            .ltout(\b2v_inst36.curr_state_RNI3E27Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_RNIPUMD_LC_8_5_6 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_RNIPUMD_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.DSW_PWROK_RNIPUMD_LC_8_5_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst36.DSW_PWROK_RNIPUMD_LC_8_5_6  (
            .in0(N__26015),
            .in1(_gnd_net_),
            .in2(N__24215),
            .in3(N__30510),
            .lcout(dsw_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_3_LC_8_5_7 .C_ON=1'b0;
    defparam \b2v_inst20.counter_3_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_3_LC_8_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst20.counter_3_LC_8_5_7  (
            .in0(N__24172),
            .in1(N__24140),
            .in2(_gnd_net_),
            .in3(N__24124),
            .lcout(\b2v_inst20.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_0_LC_8_6_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_0_LC_8_6_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_0_LC_8_6_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst5.count_0_LC_8_6_0  (
            .in0(N__24301),
            .in1(N__26940),
            .in2(_gnd_net_),
            .in3(N__27215),
            .lcout(\b2v_inst5.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36586),
            .ce(N__26800),
            .sr(N__27323));
    defparam \b2v_inst5.count_RNIH6CN3_13_LC_8_6_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIH6CN3_13_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIH6CN3_13_LC_8_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIH6CN3_13_LC_8_6_1  (
            .in0(N__24368),
            .in1(N__26798),
            .in2(_gnd_net_),
            .in3(N__24377),
            .lcout(\b2v_inst5.countZ0Z_13 ),
            .ltout(\b2v_inst5.countZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_13_LC_8_6_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_13_LC_8_6_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_13_LC_8_6_2 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst5.count_13_LC_8_6_2  (
            .in0(N__27324),
            .in1(N__26941),
            .in2(N__24371),
            .in3(N__24389),
            .lcout(\b2v_inst5.count_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36586),
            .ce(N__26800),
            .sr(N__27323));
    defparam \b2v_inst5.count_RNIMP4T1_0_LC_8_6_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIMP4T1_0_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIMP4T1_0_LC_8_6_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \b2v_inst5.count_RNIMP4T1_0_LC_8_6_3  (
            .in0(N__24359),
            .in1(N__24352),
            .in2(_gnd_net_),
            .in3(N__26796),
            .lcout(\b2v_inst5.count_i_0 ),
            .ltout(\b2v_inst5.count_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIL9B73_0_LC_8_6_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIL9B73_0_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIL9B73_0_LC_8_6_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \b2v_inst5.count_RNIL9B73_0_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__26939),
            .in2(N__24362),
            .in3(N__27214),
            .lcout(\b2v_inst5.count_rst_14 ),
            .ltout(\b2v_inst5.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_8_6_5 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_8_6_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__24353),
            .in2(N__24344),
            .in3(N__26797),
            .lcout(\b2v_inst5.un2_count_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIJ9DN3_14_LC_8_6_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIJ9DN3_14_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIJ9DN3_14_LC_8_6_6 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \b2v_inst5.count_RNIJ9DN3_14_LC_8_6_6  (
            .in0(N__26799),
            .in1(N__24328),
            .in2(N__27289),
            .in3(N__24317),
            .lcout(\b2v_inst5.countZ0Z_14 ),
            .ltout(\b2v_inst5.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIMP4T1_0_0_LC_8_6_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIMP4T1_0_0_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIMP4T1_0_0_LC_8_6_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst5.count_RNIMP4T1_0_0_LC_8_6_7  (
            .in0(N__26614),
            .in1(N__24302),
            .in2(N__24293),
            .in3(N__24290),
            .lcout(\b2v_inst5.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIU15T1_0_8_LC_8_7_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIU15T1_0_8_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIU15T1_0_8_LC_8_7_0 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \b2v_inst5.count_RNIU15T1_0_8_LC_8_7_0  (
            .in0(N__24272),
            .in1(N__24432),
            .in2(N__26848),
            .in3(N__24449),
            .lcout(\b2v_inst5.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_8_7_1 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_8_7_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_8_7_1  (
            .in0(N__27217),
            .in1(N__24460),
            .in2(N__24476),
            .in3(N__26963),
            .lcout(\b2v_inst5.count_rst_6 ),
            .ltout(\b2v_inst5.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIU15T1_8_LC_8_7_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIU15T1_8_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIU15T1_8_LC_8_7_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.count_RNIU15T1_8_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__24448),
            .in2(N__24479),
            .in3(N__26802),
            .lcout(\b2v_inst5.un2_count_1_axb_8 ),
            .ltout(\b2v_inst5.un2_count_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_8_LC_8_7_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_8_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_8_LC_8_7_3 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.count_8_LC_8_7_3  (
            .in0(N__27219),
            .in1(N__24461),
            .in2(N__24452),
            .in3(N__26964),
            .lcout(\b2v_inst5.count_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36447),
            .ce(N__26821),
            .sr(N__27303));
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_8_7_4 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_8_7_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_8_7_4  (
            .in0(N__26962),
            .in1(N__24433),
            .in2(N__24416),
            .in3(N__27216),
            .lcout(),
            .ltout(\b2v_inst5.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIH08H3_4_LC_8_7_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIH08H3_4_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIH08H3_4_LC_8_7_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst5.count_RNIH08H3_4_LC_8_7_5  (
            .in0(N__26801),
            .in1(_gnd_net_),
            .in2(N__24440),
            .in3(N__24395),
            .lcout(\b2v_inst5.countZ0Z_4 ),
            .ltout(\b2v_inst5.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_4_LC_8_7_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_4_LC_8_7_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_4_LC_8_7_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_4_LC_8_7_6  (
            .in0(N__24415),
            .in1(N__26979),
            .in2(N__24398),
            .in3(N__27220),
            .lcout(\b2v_inst5.count_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36447),
            .ce(N__26821),
            .sr(N__27303));
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_7_7 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_7_7 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_7_7  (
            .in0(N__27218),
            .in1(N__24388),
            .in2(N__26981),
            .in3(N__26536),
            .lcout(\b2v_inst5.count_rst_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_12_LC_8_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_12_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_12_LC_8_8_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \b2v_inst11.dutycycle_12_LC_8_8_0  (
            .in0(N__24812),
            .in1(N__24788),
            .in2(N__31248),
            .in3(N__24799),
            .lcout(\b2v_inst11.dutycycleZ1Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36636),
            .ce(),
            .sr(N__31037));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_12_LC_8_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_12_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_12_LC_8_8_1 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_12_LC_8_8_1  (
            .in0(N__25112),
            .in1(N__33866),
            .in2(N__25079),
            .in3(N__24827),
            .lcout(),
            .ltout(\b2v_inst11.N_396_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIANKU4_12_LC_8_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIANKU4_12_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIANKU4_12_LC_8_8_2 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNIANKU4_12_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__25321),
            .in2(N__24818),
            .in3(N__34182),
            .lcout(\b2v_inst11.N_234_N ),
            .ltout(\b2v_inst11.N_234_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICO933_12_LC_8_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICO933_12_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICO933_12_LC_8_8_3 .LUT_INIT=16'b0011101100111111;
    LogicCell40 \b2v_inst11.dutycycle_RNICO933_12_LC_8_8_3  (
            .in0(N__25056),
            .in1(N__34738),
            .in2(N__24815),
            .in3(N__33867),
            .lcout(\b2v_inst11.dutycycle_eena_9 ),
            .ltout(\b2v_inst11.dutycycle_eena_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIHFVH5_12_LC_8_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIHFVH5_12_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIHFVH5_12_LC_8_8_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIHFVH5_12_LC_8_8_4  (
            .in0(N__24803),
            .in1(N__24787),
            .in2(N__24779),
            .in3(N__31151),
            .lcout(\b2v_inst11.dutycycleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_11_LC_8_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_11_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_11_LC_8_8_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \b2v_inst11.dutycycle_11_LC_8_8_5  (
            .in0(N__31153),
            .in1(N__24767),
            .in2(N__24761),
            .in3(N__24740),
            .lcout(\b2v_inst11.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36636),
            .ce(),
            .sr(N__31037));
    defparam \b2v_inst11.dutycycle_RNICO933_11_LC_8_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICO933_11_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICO933_11_LC_8_8_6 .LUT_INIT=16'b0101011101011111;
    LogicCell40 \b2v_inst11.dutycycle_RNICO933_11_LC_8_8_6  (
            .in0(N__34739),
            .in1(N__33937),
            .in2(N__24776),
            .in3(N__25111),
            .lcout(\b2v_inst11.dutycycle_eena_7 ),
            .ltout(\b2v_inst11.dutycycle_eena_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIFCUH5_11_LC_8_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIFCUH5_11_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIFCUH5_11_LC_8_8_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIFCUH5_11_LC_8_8_7  (
            .in0(N__31152),
            .in1(N__24754),
            .in2(N__24743),
            .in3(N__24739),
            .lcout(\b2v_inst11.dutycycleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIT35D7_13_LC_8_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIT35D7_13_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIT35D7_13_LC_8_9_0 .LUT_INIT=16'b0010001010100010;
    LogicCell40 \b2v_inst11.dutycycle_RNIT35D7_13_LC_8_9_0  (
            .in0(N__31196),
            .in1(N__34743),
            .in2(N__24875),
            .in3(N__27636),
            .lcout(\b2v_inst11.dutycycle_RNIT35D7Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_11_LC_8_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_11_LC_8_9_1  (
            .in0(N__25036),
            .in1(N__25178),
            .in2(_gnd_net_),
            .in3(N__24676),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_LC_8_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_8_9_2 .LUT_INIT=16'b1100111100110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_LC_8_9_2  (
            .in0(N__33187),
            .in1(N__24632),
            .in2(N__31377),
            .in3(N__35175),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_8_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_8_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_11_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25177),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ),
            .ltout(\b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__24853),
            .in2(N__25091),
            .in3(N__25035),
            .lcout(\b2v_inst11.N_365 ),
            .ltout(\b2v_inst11.N_365_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_8_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_8_9_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_2_LC_8_9_5  (
            .in0(N__33165),
            .in1(_gnd_net_),
            .in2(N__25001),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_366 ),
            .ltout(\b2v_inst11.N_366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_1_LC_8_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_1_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_1_LC_8_9_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_1_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__33467),
            .in2(N__24998),
            .in3(N__33406),
            .lcout(\b2v_inst11.un1_func_state25_6_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIANKU4_13_LC_8_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIANKU4_13_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIANKU4_13_LC_8_9_7 .LUT_INIT=16'b1110111110101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIANKU4_13_LC_8_9_7  (
            .in0(N__24986),
            .in1(N__25312),
            .in2(N__34300),
            .in3(N__24951),
            .lcout(\b2v_inst11.N_153_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNILF063_7_LC_8_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNILF063_7_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNILF063_7_LC_8_10_0 .LUT_INIT=16'b1111101110101010;
    LogicCell40 \b2v_inst11.dutycycle_RNILF063_7_LC_8_10_0  (
            .in0(N__27622),
            .in1(N__25479),
            .in2(N__25460),
            .in3(N__25549),
            .lcout(\b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_6_LC_8_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_6_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_6_LC_8_10_1 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_6_LC_8_10_1  (
            .in0(N__33891),
            .in1(N__33281),
            .in2(_gnd_net_),
            .in3(N__29926),
            .lcout(\b2v_inst11.g2_i_a6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_LC_8_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_8_10_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_LC_8_10_2  (
            .in0(N__27662),
            .in1(N__24854),
            .in2(N__33074),
            .in3(N__33174),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDUQ02_1_LC_8_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDUQ02_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDUQ02_1_LC_8_10_3 .LUT_INIT=16'b1101110111001101;
    LogicCell40 \b2v_inst11.func_state_RNIDUQ02_1_LC_8_10_3  (
            .in0(N__34623),
            .in1(N__27389),
            .in2(N__32911),
            .in3(N__33280),
            .lcout(\b2v_inst11.func_state_RNIDUQ02Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNIDUQ02Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNILF063_0_LC_8_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNILF063_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNILF063_0_LC_8_10_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \b2v_inst11.func_state_RNILF063_0_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25325),
            .in3(N__25512),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI8H551_7_LC_8_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI8H551_7_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI8H551_7_LC_8_10_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI8H551_7_LC_8_10_5  (
            .in0(N__27575),
            .in1(N__27661),
            .in2(N__25553),
            .in3(N__25459),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_36_and_i_a2_4_0_0cf0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5ELP4_7_LC_8_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5ELP4_7_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5ELP4_7_LC_8_10_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI5ELP4_7_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__34221),
            .in2(N__25271),
            .in3(N__25268),
            .lcout(\b2v_inst11.un1_clk_100khz_36_and_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_0_LC_8_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_0_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_0_LC_8_10_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_0_LC_8_10_7  (
            .in0(N__32897),
            .in1(N__34602),
            .in2(N__34456),
            .in3(N__30895),
            .lcout(\b2v_inst11.func_state_RNI8H551Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNILBJP_1_LC_8_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNILBJP_1_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNILBJP_1_LC_8_11_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \b2v_inst11.func_state_RNILBJP_1_LC_8_11_0  (
            .in0(N__27459),
            .in1(N__27528),
            .in2(N__29637),
            .in3(N__25565),
            .lcout(),
            .ltout(\b2v_inst11.N_14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI9MT83_6_LC_8_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI9MT83_6_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI9MT83_6_LC_8_11_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst11.dutycycle_RNI9MT83_6_LC_8_11_1  (
            .in0(N__25559),
            .in1(N__27590),
            .in2(N__25262),
            .in3(N__34219),
            .lcout(\b2v_inst11.g2_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_6_0_LC_8_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_6_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_6_0_LC_8_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.func_state_RNI_6_0_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27621),
            .lcout(\b2v_inst11.func_state_RNI_6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4  (
            .in0(N__29891),
            .in1(N__30126),
            .in2(N__31364),
            .in3(N__35135),
            .lcout(\b2v_inst11.N_395 ),
            .ltout(\b2v_inst11.N_395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_5_LC_8_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_5_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_5_LC_8_11_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_5_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25223),
            .in3(N__27580),
            .lcout(\b2v_inst11.dutycycle_RNI_6Z0Z_5 ),
            .ltout(\b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI3NQD_1_LC_8_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI3NQD_1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI3NQD_1_LC_8_11_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.func_state_RNI3NQD_1_LC_8_11_6  (
            .in0(N__34016),
            .in1(N__32823),
            .in2(N__25568),
            .in3(N__35062),
            .lcout(\b2v_inst11.g0_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIA70J1_6_LC_8_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIA70J1_6_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIA70J1_6_LC_8_11_7 .LUT_INIT=16'b0000101010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNIA70J1_6_LC_8_11_7  (
            .in0(N__29886),
            .in1(N__34624),
            .in2(N__35095),
            .in3(N__25538),
            .lcout(\b2v_inst11.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_0_0_LC_8_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_0_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_0_0_LC_8_12_0 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_0_0_LC_8_12_0  (
            .in0(N__25521),
            .in1(N__33258),
            .in2(_gnd_net_),
            .in3(N__25454),
            .lcout(\b2v_inst11.un1_clk_100khz_36_and_i_o3_0_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI8H551_6_LC_8_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI8H551_6_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI8H551_6_LC_8_12_1 .LUT_INIT=16'b0000010011000100;
    LogicCell40 \b2v_inst11.count_clk_RNI8H551_6_LC_8_12_1  (
            .in0(N__33259),
            .in1(N__32874),
            .in2(N__34622),
            .in3(N__34452),
            .lcout(\b2v_inst11.g0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNILF063_0_0_LC_8_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNILF063_0_0_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNILF063_0_0_LC_8_12_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.func_state_RNILF063_0_0_LC_8_12_2  (
            .in0(N__25522),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25483),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_eena_5_d_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIANKU4_7_LC_8_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIANKU4_7_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIANKU4_7_LC_8_12_3 .LUT_INIT=16'b0011011101110111;
    LogicCell40 \b2v_inst11.dutycycle_RNIANKU4_7_LC_8_12_3  (
            .in0(N__25455),
            .in1(N__33933),
            .in2(N__25361),
            .in3(N__34277),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_eena_5_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI2IQ6C_7_LC_8_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI2IQ6C_7_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI2IQ6C_7_LC_8_12_4 .LUT_INIT=16'b0100010011000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI2IQ6C_7_LC_8_12_4  (
            .in0(N__34814),
            .in1(N__31240),
            .in2(N__25358),
            .in3(N__25355),
            .lcout(\b2v_inst11.dutycycle_RNI2IQ6CZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI4SIH2_1_LC_8_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI4SIH2_1_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI4SIH2_1_LC_8_12_5 .LUT_INIT=16'b1111010111000100;
    LogicCell40 \b2v_inst11.func_state_RNI4SIH2_1_LC_8_12_5  (
            .in0(N__27645),
            .in1(N__32875),
            .in2(N__33938),
            .in3(N__34929),
            .lcout(\b2v_inst11.count_clk_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI34G9_1_LC_8_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI34G9_1_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI34G9_1_LC_8_12_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.func_state_RNI34G9_1_LC_8_12_6  (
            .in0(N__34453),
            .in1(N__29786),
            .in2(N__35599),
            .in3(N__30820),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_1_LC_8_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_1_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_1_LC_8_12_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_1_LC_8_12_7  (
            .in0(N__33260),
            .in1(N__30286),
            .in2(N__25622),
            .in3(N__35031),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_13_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_13_0  (
            .in0(N__33501),
            .in1(N__34040),
            .in2(_gnd_net_),
            .in3(N__27803),
            .lcout(),
            .ltout(\b2v_inst11.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIICTM5_0_LC_8_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIICTM5_0_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIICTM5_0_LC_8_13_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \b2v_inst11.func_state_RNIICTM5_0_LC_8_13_1  (
            .in0(N__25619),
            .in1(N__32214),
            .in2(N__25610),
            .in3(N__28007),
            .lcout(\b2v_inst11.count_clk_en ),
            .ltout(\b2v_inst11.count_clk_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIP95D_0_LC_8_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIP95D_0_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIP95D_0_LC_8_13_2 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIP95D_0_LC_8_13_2  (
            .in0(N__25607),
            .in1(N__28025),
            .in2(N__25595),
            .in3(N__30604),
            .lcout(\b2v_inst11.count_clkZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_8_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_8_13_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_8_13_3  (
            .in0(N__25592),
            .in1(N__34066),
            .in2(N__27809),
            .in3(N__33633),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_o_N_329_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_0_LC_8_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_0_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_0_LC_8_13_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_0_LC_8_13_4  (
            .in0(N__35595),
            .in1(N__31427),
            .in2(N__25580),
            .in3(N__33419),
            .lcout(\b2v_inst11.un1_func_state25_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_1_LC_8_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_8_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_1_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__35025),
            .in2(_gnd_net_),
            .in3(N__35594),
            .lcout(\b2v_inst11.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIDQ4A1_7_LC_8_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIDQ4A1_7_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIDQ4A1_7_LC_8_13_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \b2v_inst11.count_clk_RNIDQ4A1_7_LC_8_13_6  (
            .in0(N__27844),
            .in1(_gnd_net_),
            .in2(N__33513),
            .in3(N__34041),
            .lcout(\b2v_inst11.count_clk_RNIDQ4A1Z0Z_7 ),
            .ltout(\b2v_inst11.count_clk_RNIDQ4A1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_2_LC_8_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_2_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_2_LC_8_13_7 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_2_LC_8_13_7  (
            .in0(N__30914),
            .in1(N__25577),
            .in2(N__25571),
            .in3(N__35026),
            .lcout(\b2v_inst11.un1_func_state25_6_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNINHRI_2_LC_8_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNINHRI_2_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNINHRI_2_LC_8_14_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.count_clk_RNINHRI_2_LC_8_14_0  (
            .in0(N__25679),
            .in1(N__28487),
            .in2(N__25637),
            .in3(N__30612),
            .lcout(\b2v_inst11.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_2_LC_8_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_2_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_2_LC_8_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_2_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25633),
            .lcout(\b2v_inst11.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36656),
            .ce(N__28583),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIPKSI_3_LC_8_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIPKSI_3_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIPKSI_3_LC_8_14_2 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \b2v_inst11.count_clk_RNIPKSI_3_LC_8_14_2  (
            .in0(N__25847),
            .in1(N__28485),
            .in2(N__30638),
            .in3(N__25673),
            .lcout(\b2v_inst11.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_3_LC_8_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_3_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_3_LC_8_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_3_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25846),
            .lcout(\b2v_inst11.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36656),
            .ce(N__28583),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIRNTI_4_LC_8_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIRNTI_4_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIRNTI_4_LC_8_14_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.count_clk_RNIRNTI_4_LC_8_14_4  (
            .in0(N__25667),
            .in1(N__28488),
            .in2(N__25817),
            .in3(N__30613),
            .lcout(\b2v_inst11.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_4_LC_8_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_4_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_4_LC_8_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_4_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25813),
            .lcout(\b2v_inst11.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36656),
            .ce(N__28583),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVTVI_6_LC_8_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVTVI_6_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVTVI_6_LC_8_14_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.count_clk_RNIVTVI_6_LC_8_14_6  (
            .in0(N__25661),
            .in1(N__28486),
            .in2(N__25751),
            .in3(N__30611),
            .lcout(\b2v_inst11.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_6_LC_8_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_6_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_6_LC_8_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_6_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25747),
            .lcout(\b2v_inst11.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36656),
            .ce(N__28583),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_8_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_8_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__28169),
            .in2(N__28219),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_8_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_8_15_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_8_15_1  (
            .in0(N__28127),
            .in1(N__25654),
            .in2(_gnd_net_),
            .in3(N__25625),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_8_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_8_15_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_8_15_2  (
            .in0(N__28105),
            .in1(N__25864),
            .in2(_gnd_net_),
            .in3(N__25838),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_8_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_8_15_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_8_15_3  (
            .in0(N__28128),
            .in1(_gnd_net_),
            .in2(N__25835),
            .in3(N__25805),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_8_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_8_15_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_8_15_4  (
            .in0(N__28103),
            .in1(N__25802),
            .in2(_gnd_net_),
            .in3(N__25772),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_8_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_8_15_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_8_15_5  (
            .in0(N__28129),
            .in1(_gnd_net_),
            .in2(N__25769),
            .in3(N__25739),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_8_15_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_8_15_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_8_15_6  (
            .in0(N__28104),
            .in1(N__28413),
            .in2(_gnd_net_),
            .in3(N__25736),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_8_15_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_8_15_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_8_15_7  (
            .in0(N__28126),
            .in1(N__25733),
            .in2(_gnd_net_),
            .in3(N__25709),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_8_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_8_16_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_8_16_0  (
            .in0(N__28097),
            .in1(N__25706),
            .in2(_gnd_net_),
            .in3(N__25685),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_8_16_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_8_16_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_8_16_1  (
            .in0(N__28108),
            .in1(N__28337),
            .in2(_gnd_net_),
            .in3(N__25682),
            .lcout(\b2v_inst11.count_clk_1_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_8_16_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_8_16_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_8_16_2  (
            .in0(N__28098),
            .in1(N__28351),
            .in2(_gnd_net_),
            .in3(N__25940),
            .lcout(\b2v_inst11.count_clk_1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_10 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_8_16_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_8_16_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_8_16_3  (
            .in0(N__28107),
            .in1(N__28298),
            .in2(_gnd_net_),
            .in3(N__25937),
            .lcout(\b2v_inst11.count_clk_1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_8_16_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_8_16_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_8_16_4  (
            .in0(N__28099),
            .in1(N__28358),
            .in2(_gnd_net_),
            .in3(N__25934),
            .lcout(\b2v_inst11.count_clk_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_8_16_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_8_16_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_8_16_5  (
            .in0(N__28106),
            .in1(N__25931),
            .in2(_gnd_net_),
            .in3(N__25910),
            .lcout(\b2v_inst11.count_clk_1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_8_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_8_16_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_8_16_6  (
            .in0(N__25907),
            .in1(N__28109),
            .in2(_gnd_net_),
            .in3(N__25901),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIN3CI_11_LC_8_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIN3CI_11_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIN3CI_11_LC_8_16_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \b2v_inst11.count_clk_RNIN3CI_11_LC_8_16_7  (
            .in0(N__25889),
            .in1(N__25883),
            .in2(N__28582),
            .in3(N__30574),
            .lcout(\b2v_inst11.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_9_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_9_1_0 .LUT_INIT=16'b0010110000100000;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m4_LC_9_1_0  (
            .in0(N__29247),
            .in1(N__29318),
            .in2(N__29293),
            .in3(N__26133),
            .lcout(),
            .ltout(\b2v_inst36.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNIT62Q_0_LC_9_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIT62Q_0_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIT62Q_0_LC_9_1_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.curr_state_RNIT62Q_0_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__26036),
            .in2(N__25871),
            .in3(N__30558),
            .lcout(\b2v_inst36.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_9_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_9_1_2 .LUT_INIT=16'b0000001100001010;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m6_LC_9_1_2  (
            .in0(N__29248),
            .in1(N__26132),
            .in2(N__26039),
            .in3(N__29326),
            .lcout(\b2v_inst36.curr_state_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_0_LC_9_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_0_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_0_LC_9_1_3 .LUT_INIT=16'b0101100000001000;
    LogicCell40 \b2v_inst36.curr_state_0_LC_9_1_3  (
            .in0(N__29284),
            .in1(N__29245),
            .in2(N__29334),
            .in3(N__26152),
            .lcout(\b2v_inst36.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36234),
            .ce(N__32174),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_1_LC_9_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_1_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_1_LC_9_1_4 .LUT_INIT=16'b0000000000101110;
    LogicCell40 \b2v_inst36.curr_state_1_LC_9_1_4  (
            .in0(N__29246),
            .in1(N__29325),
            .in2(N__26169),
            .in3(N__29285),
            .lcout(\b2v_inst36.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36234),
            .ce(N__32174),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNIU72Q_1_LC_9_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIU72Q_1_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIU72Q_1_LC_9_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst36.curr_state_RNIU72Q_1_LC_9_1_5  (
            .in0(N__26030),
            .in1(N__26024),
            .in2(_gnd_net_),
            .in3(N__30557),
            .lcout(\b2v_inst36.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNIRQCA_0_LC_9_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIRQCA_0_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIRQCA_0_LC_9_1_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \b2v_inst36.curr_state_RNIRQCA_0_LC_9_1_6  (
            .in0(N__30559),
            .in1(N__29249),
            .in2(N__26018),
            .in3(N__29282),
            .lcout(\b2v_inst36.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_LC_9_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.DSW_PWROK_LC_9_1_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \b2v_inst36.DSW_PWROK_LC_9_1_7  (
            .in0(N__29283),
            .in1(_gnd_net_),
            .in2(N__29333),
            .in3(N__29244),
            .lcout(\b2v_inst36.DSW_PWROK_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36234),
            .ce(N__32174),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_8_LC_9_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_8_LC_9_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_8_LC_9_2_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.count_8_LC_9_2_0  (
            .in0(N__26154),
            .in1(N__25962),
            .in2(N__26003),
            .in3(N__28935),
            .lcout(\b2v_inst36.count_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36450),
            .ce(N__29148),
            .sr(N__28982));
    defparam \b2v_inst36.count_RNIPT1I1_8_LC_9_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIPT1I1_8_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIPT1I1_8_LC_9_2_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst36.count_RNIPT1I1_8_LC_9_2_1  (
            .in0(N__29106),
            .in1(N__25982),
            .in2(_gnd_net_),
            .in3(N__25976),
            .lcout(\b2v_inst36.countZ0Z_8 ),
            .ltout(\b2v_inst36.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI4VQN1_0_10_LC_9_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI4VQN1_0_10_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI4VQN1_0_10_LC_9_2_2 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \b2v_inst36.count_RNI4VQN1_0_10_LC_9_2_2  (
            .in0(N__29149),
            .in1(N__26075),
            .in2(N__25943),
            .in3(N__26213),
            .lcout(),
            .ltout(\b2v_inst36.un12_clk_100khz_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNILGID6_1_LC_9_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNILGID6_1_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNILGID6_1_LC_9_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNILGID6_1_LC_9_2_3  (
            .in0(N__26255),
            .in1(N__26249),
            .in2(N__26243),
            .in3(N__26240),
            .lcout(),
            .ltout(\b2v_inst36.un12_clk_100khz_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI0RKG9_6_LC_9_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI0RKG9_6_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI0RKG9_6_LC_9_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNI0RKG9_6_LC_9_2_4  (
            .in0(N__26228),
            .in1(N__26342),
            .in2(N__26219),
            .in3(N__26303),
            .lcout(\b2v_inst36.N_1_i ),
            .ltout(\b2v_inst36.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_9_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_9_2_5 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_9_2_5  (
            .in0(N__28936),
            .in1(N__26200),
            .in2(N__26216),
            .in3(N__26189),
            .lcout(\b2v_inst36.count_rst_4 ),
            .ltout(\b2v_inst36.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI4VQN1_10_LC_9_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI4VQN1_10_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI4VQN1_10_LC_9_2_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNI4VQN1_10_LC_9_2_6  (
            .in0(_gnd_net_),
            .in1(N__26074),
            .in2(N__26207),
            .in3(N__29107),
            .lcout(\b2v_inst36.un2_count_1_axb_10 ),
            .ltout(\b2v_inst36.un2_count_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_10_LC_9_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_10_LC_9_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_10_LC_9_2_7 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.count_10_LC_9_2_7  (
            .in0(N__28934),
            .in1(N__26188),
            .in2(N__26177),
            .in3(N__26155),
            .lcout(\b2v_inst36.count_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36450),
            .ce(N__29148),
            .sr(N__28982));
    defparam \b2v_inst36.count_4_LC_9_3_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_4_LC_9_3_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_4_LC_9_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_4_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26060),
            .lcout(\b2v_inst36.count_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36244),
            .ce(N__29132),
            .sr(N__28962));
    defparam \b2v_inst36.count_RNICQ3V_6_LC_9_3_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNICQ3V_6_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNICQ3V_6_LC_9_3_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNICQ3V_6_LC_9_3_1  (
            .in0(N__26350),
            .in1(N__29120),
            .in2(_gnd_net_),
            .in3(N__26367),
            .lcout(\b2v_inst36.un2_count_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_6_LC_9_3_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_6_LC_9_3_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_6_LC_9_3_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_6_LC_9_3_2  (
            .in0(N__26368),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36244),
            .ce(N__29132),
            .sr(N__28962));
    defparam \b2v_inst36.count_RNIHHTH1_4_LC_9_3_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIHHTH1_4_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIHHTH1_4_LC_9_3_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \b2v_inst36.count_RNIHHTH1_4_LC_9_3_3  (
            .in0(N__26059),
            .in1(N__29119),
            .in2(_gnd_net_),
            .in3(N__26051),
            .lcout(\b2v_inst36.countZ0Z_4 ),
            .ltout(\b2v_inst36.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNICQ3V_0_6_LC_9_3_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNICQ3V_0_6_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNICQ3V_0_6_LC_9_3_4 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \b2v_inst36.count_RNICQ3V_0_6_LC_9_3_4  (
            .in0(N__29122),
            .in1(N__26369),
            .in2(N__26354),
            .in3(N__26351),
            .lcout(\b2v_inst36.un12_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIPRQ41_12_LC_9_3_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIPRQ41_12_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIPRQ41_12_LC_9_3_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIPRQ41_12_LC_9_3_5  (
            .in0(N__26330),
            .in1(N__29121),
            .in2(_gnd_net_),
            .in3(N__26316),
            .lcout(\b2v_inst36.un2_count_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_12_LC_9_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_12_LC_9_3_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_12_LC_9_3_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_12_LC_9_3_6  (
            .in0(N__26317),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36244),
            .ce(N__29132),
            .sr(N__28962));
    defparam \b2v_inst36.count_RNIPRQ41_0_12_LC_9_3_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIPRQ41_0_12_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIPRQ41_0_12_LC_9_3_7 .LUT_INIT=16'b0000001100010001;
    LogicCell40 \b2v_inst36.count_RNIPRQ41_0_12_LC_9_3_7  (
            .in0(N__26329),
            .in1(N__29189),
            .in2(N__26321),
            .in3(N__29133),
            .lcout(\b2v_inst36.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_3_LC_9_4_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_3_LC_9_4_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_3_LC_9_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_3_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26575),
            .lcout(\b2v_inst5.count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36356),
            .ce(N__26863),
            .sr(N__27302));
    defparam \b2v_inst5.count_RNIBN4H3_1_LC_9_4_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIBN4H3_1_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIBN4H3_1_LC_9_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst5.count_RNIBN4H3_1_LC_9_4_1  (
            .in0(N__26282),
            .in1(N__26297),
            .in2(_gnd_net_),
            .in3(N__26825),
            .lcout(\b2v_inst5.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_1_LC_9_4_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_1_LC_9_4_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_1_LC_9_4_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_1_LC_9_4_2  (
            .in0(N__26296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36356),
            .ce(N__26863),
            .sr(N__27302));
    defparam \b2v_inst5.count_RNIDQ5H3_2_LC_9_4_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIDQ5H3_2_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIDQ5H3_2_LC_9_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst5.count_RNIDQ5H3_2_LC_9_4_3  (
            .in0(N__26276),
            .in1(N__26261),
            .in2(_gnd_net_),
            .in3(N__26826),
            .lcout(\b2v_inst5.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_2_LC_9_4_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_2_LC_9_4_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_2_LC_9_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_2_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26275),
            .lcout(\b2v_inst5.count_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36356),
            .ce(N__26863),
            .sr(N__27302));
    defparam \b2v_inst5.count_RNIFT6H3_3_LC_9_4_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIFT6H3_3_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIFT6H3_3_LC_9_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst5.count_RNIFT6H3_3_LC_9_4_5  (
            .in0(N__26576),
            .in1(N__26561),
            .in2(_gnd_net_),
            .in3(N__26827),
            .lcout(\b2v_inst5.countZ0Z_3 ),
            .ltout(\b2v_inst5.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI_1_LC_9_4_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI_1_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI_1_LC_9_4_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \b2v_inst5.count_RNI_1_LC_9_4_6  (
            .in0(N__26540),
            .in1(N__26515),
            .in2(N__26501),
            .in3(N__26494),
            .lcout(\b2v_inst5.un12_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIJ39H3_5_LC_9_4_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIJ39H3_5_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIJ39H3_5_LC_9_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst5.count_RNIJ39H3_5_LC_9_4_7  (
            .in0(N__26903),
            .in1(N__26882),
            .in2(_gnd_net_),
            .in3(N__26828),
            .lcout(\b2v_inst5.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI7BCA2_0_10_LC_9_5_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI7BCA2_0_10_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI7BCA2_0_10_LC_9_5_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \b2v_inst5.count_RNI7BCA2_0_10_LC_9_5_0  (
            .in0(N__26633),
            .in1(N__26815),
            .in2(N__26455),
            .in3(N__27015),
            .lcout(),
            .ltout(\b2v_inst5.un12_clk_100khz_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI870S9_8_LC_9_5_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI870S9_8_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI870S9_8_LC_9_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.count_RNI870S9_8_LC_9_5_1  (
            .in0(N__26480),
            .in1(N__26471),
            .in2(N__26462),
            .in3(N__26375),
            .lcout(\b2v_inst5.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI7BCA2_10_LC_9_5_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI7BCA2_10_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI7BCA2_10_LC_9_5_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \b2v_inst5.count_RNI7BCA2_10_LC_9_5_2  (
            .in0(N__26632),
            .in1(_gnd_net_),
            .in2(N__26456),
            .in3(N__26813),
            .lcout(\b2v_inst5.un2_count_1_axb_10 ),
            .ltout(\b2v_inst5.un2_count_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_10_LC_9_5_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_10_LC_9_5_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_10_LC_9_5_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_10_LC_9_5_3  (
            .in0(N__26666),
            .in1(N__26975),
            .in2(N__26459),
            .in3(N__27330),
            .lcout(\b2v_inst5.count_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36350),
            .ce(N__26820),
            .sr(N__27329));
    defparam \b2v_inst5.count_RNI3QEK5_11_LC_9_5_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI3QEK5_11_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI3QEK5_11_LC_9_5_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst5.count_RNI3QEK5_11_LC_9_5_4  (
            .in0(N__26441),
            .in1(N__26425),
            .in2(N__26411),
            .in3(N__26402),
            .lcout(\b2v_inst5.un12_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIRFDH3_9_LC_9_5_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIRFDH3_9_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIRFDH3_9_LC_9_5_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst5.count_RNIRFDH3_9_LC_9_5_5  (
            .in0(N__26814),
            .in1(_gnd_net_),
            .in2(N__26675),
            .in3(N__26909),
            .lcout(\b2v_inst5.countZ0Z_9 ),
            .ltout(\b2v_inst5.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_9_LC_9_5_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_9_LC_9_5_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_9_LC_9_5_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst5.count_9_LC_9_5_6  (
            .in0(N__26974),
            .in1(N__27293),
            .in2(N__26678),
            .in3(N__26999),
            .lcout(\b2v_inst5.count_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36350),
            .ce(N__26820),
            .sr(N__27329));
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_9_5_7 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_9_5_7 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_9_5_7  (
            .in0(N__26665),
            .in1(N__26973),
            .in2(N__27325),
            .in3(N__26647),
            .lcout(\b2v_inst5.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIKEUB2_1_LC_9_6_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIKEUB2_1_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIKEUB2_1_LC_9_6_0 .LUT_INIT=16'b0011001111110000;
    LogicCell40 \b2v_inst5.curr_state_RNIKEUB2_1_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__32248),
            .in2(N__32237),
            .in3(N__30391),
            .lcout(\b2v_inst5.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst5.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI_1_LC_9_6_1 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI_1_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI_1_LC_9_6_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst5.curr_state_RNI_1_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26624),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.curr_state_RNIZ0Z_1 ),
            .ltout(\b2v_inst5.curr_state_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIRH7S1_0_LC_9_6_2 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIRH7S1_0_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIRH7S1_0_LC_9_6_2 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \b2v_inst5.curr_state_RNIRH7S1_0_LC_9_6_2  (
            .in0(N__32986),
            .in1(N__27357),
            .in2(N__26621),
            .in3(N__31124),
            .lcout(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ),
            .ltout(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNILCEN3_15_LC_9_6_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNILCEN3_15_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNILCEN3_15_LC_9_6_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst5.count_RNILCEN3_15_LC_9_6_3  (
            .in0(N__26600),
            .in1(_gnd_net_),
            .in2(N__26618),
            .in3(N__26588),
            .lcout(\b2v_inst5.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_15_LC_9_6_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_15_LC_9_6_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_15_LC_9_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_15_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26599),
            .lcout(\b2v_inst5.count_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36360),
            .ce(N__26819),
            .sr(N__27331));
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_9_6_5 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_9_6_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_9_6_5  (
            .in0(N__26582),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26938),
            .lcout(N_413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_9_6_6 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_9_6_6 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_9_6_6  (
            .in0(N__27019),
            .in1(N__26998),
            .in2(N__26980),
            .in3(N__27213),
            .lcout(\b2v_inst5.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_5_LC_9_6_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_5_LC_9_6_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_5_LC_9_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_5_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26902),
            .lcout(\b2v_inst5.count_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36360),
            .ce(N__26819),
            .sr(N__27331));
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_9_7_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_9_7_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst5.curr_state_RNI65HI_0_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__26696),
            .in2(N__30602),
            .in3(N__26717),
            .lcout(\b2v_inst5.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst5.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_9_7_1 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_9_7_1 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m6_i_LC_9_7_1  (
            .in0(N__32988),
            .in1(N__27382),
            .in2(N__26720),
            .in3(N__26707),
            .lcout(\b2v_inst5.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_LC_9_7_2 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.RSMRSTn_LC_9_7_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst5.RSMRSTn_LC_9_7_2  (
            .in0(N__27381),
            .in1(N__32987),
            .in2(_gnd_net_),
            .in3(N__26690),
            .lcout(RSMRSTn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36448),
            .ce(N__32176),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_7_3 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_7_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_7_3  (
            .in0(N__27358),
            .in1(N__27513),
            .in2(_gnd_net_),
            .in3(N__26706),
            .lcout(\b2v_inst5.m4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI65HI_0_0_LC_9_7_4 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI65HI_0_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI65HI_0_0_LC_9_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst5.curr_state_RNI65HI_0_0_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26689),
            .lcout(\b2v_inst5.N_2898_i ),
            .ltout(\b2v_inst5.N_2898_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_0_LC_9_7_5 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_0_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_0_LC_9_7_5 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \b2v_inst5.curr_state_0_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__27512),
            .in2(N__26711),
            .in3(N__26708),
            .lcout(\b2v_inst5.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36448),
            .ce(N__32176),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNID8DP1_0_LC_9_7_6 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNID8DP1_0_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNID8DP1_0_LC_9_7_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst5.curr_state_RNID8DP1_0_LC_9_7_6  (
            .in0(N__32990),
            .in1(N__27373),
            .in2(_gnd_net_),
            .in3(N__26688),
            .lcout(curr_state_RNID8DP1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIVF6A1_0_LC_9_7_7 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIVF6A1_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIVF6A1_0_LC_9_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.curr_state_RNIVF6A1_0_LC_9_7_7  (
            .in0(N__32989),
            .in1(N__27383),
            .in2(N__27362),
            .in3(N__30420),
            .lcout(\b2v_inst5.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_8_1_LC_9_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_8_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_8_1_LC_9_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.func_state_RNI_8_1_LC_9_8_0  (
            .in0(N__33385),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_172_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI5DLR_1_LC_9_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI5DLR_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI5DLR_1_LC_9_8_1 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \b2v_inst11.func_state_RNI5DLR_1_LC_9_8_1  (
            .in0(N__34615),
            .in1(N__32910),
            .in2(_gnd_net_),
            .in3(N__35096),
            .lcout(\b2v_inst11.un1_clk_100khz_2_i_o3_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_9_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_9_8_2 .LUT_INIT=16'b0101011111011111;
    LogicCell40 \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_9_8_2  (
            .in0(N__34619),
            .in1(N__29623),
            .in2(N__27445),
            .in3(N__27495),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_6_1_LC_9_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_6_1_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_6_1_LC_9_8_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst11.func_state_RNI_6_1_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__33384),
            .in2(_gnd_net_),
            .in3(N__33293),
            .lcout(),
            .ltout(\b2v_inst11.N_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_9_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_9_8_4 .LUT_INIT=16'b1101110011111111;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_9_8_4  (
            .in0(N__28246),
            .in1(N__33898),
            .in2(N__27056),
            .in3(N__34052),
            .lcout(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_9_8_5 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_9_8_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst5.RSMRSTn_RNI8DFE_LC_9_8_5  (
            .in0(N__27046),
            .in1(_gnd_net_),
            .in2(N__27514),
            .in3(N__27432),
            .lcout(rsmrstn),
            .ltout(rsmrstn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_9_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_9_8_6 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_9_8_6  (
            .in0(N__34405),
            .in1(N__30309),
            .in2(N__27053),
            .in3(N__29624),
            .lcout(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_8_7 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_8_7  (
            .in0(N__27499),
            .in1(N__29570),
            .in2(N__27050),
            .in3(N__27433),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_9_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_9_9_0 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_9_9_0  (
            .in0(N__32907),
            .in1(N__34614),
            .in2(_gnd_net_),
            .in3(N__34181),
            .lcout(\b2v_inst11.N_168 ),
            .ltout(\b2v_inst11.N_168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_9_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_9_9_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_9_9_1  (
            .in0(N__30515),
            .in1(N__32908),
            .in2(N__27536),
            .in3(N__34625),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_9_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_9_9_2 .LUT_INIT=16'b0101110101111111;
    LogicCell40 \b2v_inst11.VCCST_EN_i_0_o3_0_LC_9_9_2  (
            .in0(N__32906),
            .in1(N__30514),
            .in2(N__27527),
            .in3(N__27458),
            .lcout(VCCST_EN_i_0_o3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIDQ4A1_6_LC_9_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIDQ4A1_6_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIDQ4A1_6_LC_9_9_3 .LUT_INIT=16'b1010101010111111;
    LogicCell40 \b2v_inst11.count_clk_RNIDQ4A1_6_LC_9_9_3  (
            .in0(N__33477),
            .in1(N__27573),
            .in2(N__27982),
            .in3(N__33079),
            .lcout(),
            .ltout(\b2v_inst11.count_clk_RNIDQ4A1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIQK9K2_6_LC_9_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIQK9K2_6_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIQK9K2_6_LC_9_9_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \b2v_inst11.count_clk_RNIQK9K2_6_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__33407),
            .in2(N__27407),
            .in3(N__27404),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIH3DN3_6_LC_9_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIH3DN3_6_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIH3DN3_6_LC_9_9_5 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \b2v_inst11.count_clk_RNIH3DN3_6_LC_9_9_5  (
            .in0(N__34884),
            .in1(_gnd_net_),
            .in2(N__27398),
            .in3(N__34432),
            .lcout(\b2v_inst11.N_186_i ),
            .ltout(\b2v_inst11.N_186_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIN1E71_2_LC_9_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIN1E71_2_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIN1E71_2_LC_9_9_6 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \b2v_inst11.dutycycle_RNIN1E71_2_LC_9_9_6  (
            .in0(N__33098),
            .in1(N__32909),
            .in2(N__27395),
            .in3(N__34883),
            .lcout(),
            .ltout(\b2v_inst11.N_115_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAEUL3_2_LC_9_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAEUL3_2_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAEUL3_2_LC_9_9_7 .LUT_INIT=16'b0000110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIAEUL3_2_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__31211),
            .in2(N__27392),
            .in3(N__34737),
            .lcout(\b2v_inst11.dutycycle_RNIAEUL3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_0_1_LC_9_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_0_1_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_0_1_LC_9_10_0 .LUT_INIT=16'b0101110100000000;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_0_1_LC_9_10_0  (
            .in0(N__34601),
            .in1(N__32905),
            .in2(N__34454),
            .in3(N__35094),
            .lcout(\b2v_inst11.N_381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_9_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_9_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_6_LC_9_10_2  (
            .in0(N__29797),
            .in1(N__33304),
            .in2(N__27785),
            .in3(N__29942),
            .lcout(\b2v_inst11.g0_i_a7_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIUCAD1_0_0_LC_9_10_3 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIUCAD1_0_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIUCAD1_0_0_LC_9_10_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \b2v_inst16.curr_state_RNIUCAD1_0_0_LC_9_10_3  (
            .in0(N__27769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27740),
            .lcout(\b2v_inst16.N_268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_LC_9_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_LC_9_10_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_LC_9_10_4  (
            .in0(N__34014),
            .in1(N__30893),
            .in2(N__27974),
            .in3(N__27668),
            .lcout(\b2v_inst11.N_159 ),
            .ltout(\b2v_inst11.N_159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_4_0_LC_9_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_4_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_4_0_LC_9_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_4_0_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27653),
            .in3(N__27574),
            .lcout(\b2v_inst11.N_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI2MQD_0_LC_9_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI2MQD_0_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI2MQD_0_LC_9_10_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.func_state_RNI2MQD_0_LC_9_10_6  (
            .in0(N__34600),
            .in1(N__27579),
            .in2(N__27975),
            .in3(N__30894),
            .lcout(\b2v_inst11.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_ss0_i_0_a2_2_LC_9_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_ss0_i_0_a2_2_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_1_ss0_i_0_a2_2_LC_9_10_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \b2v_inst11.func_state_1_ss0_i_0_a2_2_LC_9_10_7  (
            .in0(N__32904),
            .in1(N__34599),
            .in2(_gnd_net_),
            .in3(N__34220),
            .lcout(\b2v_inst11.func_state_1_ss0_i_0_a2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_9_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_9_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_9_11_0  (
            .in0(N__30778),
            .in1(N__34015),
            .in2(N__35108),
            .in3(N__35600),
            .lcout(\b2v_inst11.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_LC_9_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_9_11_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_LC_9_11_1  (
            .in0(N__33716),
            .in1(N__31312),
            .in2(N__30144),
            .in3(N__29890),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_0 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_9_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_9_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_9_11_2  (
            .in0(N__30777),
            .in1(N__27584),
            .in2(N__27539),
            .in3(N__30896),
            .lcout(\b2v_inst11.N_406 ),
            .ltout(\b2v_inst11.N_406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVT4P1_1_LC_9_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVT4P1_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVT4P1_1_LC_9_11_3 .LUT_INIT=16'b0000001100001111;
    LogicCell40 \b2v_inst11.func_state_RNIVT4P1_1_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__34748),
            .in2(N__27872),
            .in3(N__35084),
            .lcout(\b2v_inst11.func_state_1_m2_ns_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_LC_9_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_0_LC_9_11_4 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \b2v_inst11.func_state_0_LC_9_11_4  (
            .in0(N__27869),
            .in1(N__28016),
            .in2(N__33632),
            .in3(N__28284),
            .lcout(\b2v_inst11.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36503),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_en_LC_9_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_en_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_en_LC_9_11_5 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \b2v_inst11.func_state_en_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__32824),
            .in2(N__32224),
            .in3(N__34894),
            .lcout(\b2v_inst11.func_state_enZ0 ),
            .ltout(\b2v_inst11.func_state_enZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDHTPG_0_LC_9_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDHTPG_0_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDHTPG_0_LC_9_11_6 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \b2v_inst11.func_state_RNIDHTPG_0_LC_9_11_6  (
            .in0(N__27868),
            .in1(N__33618),
            .in2(N__27860),
            .in3(N__28015),
            .lcout(\b2v_inst11.func_state ),
            .ltout(\b2v_inst11.func_state_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_0_LC_9_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_9_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.func_state_RNI_1_0_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27857),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_2946_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI5DLR_0_LC_9_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI5DLR_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI5DLR_0_LC_9_12_0 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \b2v_inst11.func_state_RNI5DLR_0_LC_9_12_0  (
            .in0(N__30290),
            .in1(N__35030),
            .in2(N__27854),
            .in3(N__30883),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINIV94_0_LC_9_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINIV94_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINIV94_0_LC_9_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.func_state_RNINIV94_0_LC_9_12_1  (
            .in0(N__27807),
            .in1(N__27823),
            .in2(N__27833),
            .in3(N__27830),
            .lcout(\b2v_inst11.func_state_RNINIV94_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF1Q43_0_LC_9_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF1Q43_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF1Q43_0_LC_9_12_2 .LUT_INIT=16'b0011011101110111;
    LogicCell40 \b2v_inst11.func_state_RNIF1Q43_0_LC_9_12_2  (
            .in0(N__27824),
            .in1(N__27808),
            .in2(N__30307),
            .in3(N__30884),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m2_ns_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINCPR4_0_LC_9_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINCPR4_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINCPR4_0_LC_9_12_3 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \b2v_inst11.func_state_RNINCPR4_0_LC_9_12_3  (
            .in0(N__27928),
            .in1(N__30841),
            .in2(N__27788),
            .in3(N__35586),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m2_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIPBBTD_0_LC_9_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIPBBTD_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIPBBTD_0_LC_9_12_4 .LUT_INIT=16'b0000001110001011;
    LogicCell40 \b2v_inst11.func_state_RNIPBBTD_0_LC_9_12_4  (
            .in0(N__30761),
            .in1(N__27884),
            .in2(N__28019),
            .in3(N__27927),
            .lcout(\b2v_inst11.func_state_1_m2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNID7Q51_0_LC_9_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNID7Q51_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNID7Q51_0_LC_9_12_5 .LUT_INIT=16'b0100110000000100;
    LogicCell40 \b2v_inst11.func_state_RNID7Q51_0_LC_9_12_5  (
            .in0(N__30882),
            .in1(N__34085),
            .in2(N__35072),
            .in3(N__35584),
            .lcout(\b2v_inst11.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_9_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_9_12_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_9_12_6  (
            .in0(N__34433),
            .in1(N__34201),
            .in2(N__30306),
            .in3(N__30623),
            .lcout(\b2v_inst11.N_382 ),
            .ltout(\b2v_inst11.N_382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI794G3_1_LC_9_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI794G3_1_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI794G3_1_LC_9_12_7 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \b2v_inst11.func_state_RNI794G3_1_LC_9_12_7  (
            .in0(N__28001),
            .in1(N__35585),
            .in2(N__27992),
            .in3(N__34048),
            .lcout(\b2v_inst11.func_state_1_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIHJNV7_0_LC_9_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIHJNV7_0_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIHJNV7_0_LC_9_13_1 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNIHJNV7_0_LC_9_13_1  (
            .in0(N__27989),
            .in1(N__31239),
            .in2(N__27983),
            .in3(N__27944),
            .lcout(\b2v_inst11.dutycycle_RNIHJNV7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI98MHC_1_LC_9_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI98MHC_1_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI98MHC_1_LC_9_13_2 .LUT_INIT=16'b1101110100001111;
    LogicCell40 \b2v_inst11.func_state_RNI98MHC_1_LC_9_13_2  (
            .in0(N__30757),
            .in1(N__27932),
            .in2(N__27914),
            .in3(N__27883),
            .lcout(\b2v_inst11.func_state_1_m2_1 ),
            .ltout(\b2v_inst11.func_state_1_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIUE8EF_1_LC_9_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIUE8EF_1_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIUE8EF_1_LC_9_13_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst11.func_state_RNIUE8EF_1_LC_9_13_3  (
            .in0(N__28258),
            .in1(N__33617),
            .in2(N__27905),
            .in3(N__28285),
            .lcout(\b2v_inst11.func_stateZ0Z_0 ),
            .ltout(\b2v_inst11.func_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI57FD1_0_1_LC_9_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI57FD1_0_1_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI57FD1_0_1_LC_9_13_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.func_state_RNI57FD1_0_1_LC_9_13_4  (
            .in0(N__30308),
            .in1(N__30603),
            .in2(N__27902),
            .in3(N__34200),
            .lcout(),
            .ltout(\b2v_inst11.N_338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIHVOG4_1_LC_9_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIHVOG4_1_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIHVOG4_1_LC_9_13_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \b2v_inst11.func_state_RNIHVOG4_1_LC_9_13_5  (
            .in0(N__28229),
            .in1(N__27899),
            .in2(N__27887),
            .in3(N__34747),
            .lcout(\b2v_inst11.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_LC_9_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_1_LC_9_13_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst11.func_state_1_LC_9_13_6  (
            .in0(N__28286),
            .in1(N__28268),
            .in2(N__28262),
            .in3(N__33622),
            .lcout(\b2v_inst11.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36661),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_1_LC_9_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_9_13_7 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \b2v_inst11.func_state_RNI_1_1_LC_9_13_7  (
            .in0(N__33418),
            .in1(N__28247),
            .in2(_gnd_net_),
            .in3(N__35083),
            .lcout(\b2v_inst11.func_state_1_m2s2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_LC_9_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_LC_9_14_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_LC_9_14_0  (
            .in0(N__28090),
            .in1(N__28223),
            .in2(_gnd_net_),
            .in3(N__28155),
            .lcout(\b2v_inst11.count_clk_RNIZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_0_LC_9_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_0_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_0_LC_9_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.count_clk_0_LC_9_14_1  (
            .in0(N__28156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28089),
            .lcout(\b2v_inst11.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36657),
            .ce(N__28572),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI8F1AB_2_LC_9_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI8F1AB_2_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI8F1AB_2_LC_9_14_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_off_RNI8F1AB_2_LC_9_14_2  (
            .in0(N__35681),
            .in1(N__35886),
            .in2(_gnd_net_),
            .in3(N__35699),
            .lcout(\b2v_inst11.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIAI2AB_3_LC_9_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIAI2AB_3_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIAI2AB_3_LC_9_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_off_RNIAI2AB_3_LC_9_14_3  (
            .in0(N__35887),
            .in1(N__36728),
            .in2(_gnd_net_),
            .in3(N__36746),
            .lcout(\b2v_inst11.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNICA5EB_13_LC_9_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNICA5EB_13_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNICA5EB_13_LC_9_14_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_off_RNICA5EB_13_LC_9_14_4  (
            .in0(N__35711),
            .in1(N__35890),
            .in2(_gnd_net_),
            .in3(N__35726),
            .lcout(\b2v_inst11.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNICL3AB_4_LC_9_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNICL3AB_4_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNICL3AB_4_LC_9_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_off_RNICL3AB_4_LC_9_14_5  (
            .in0(N__35888),
            .in1(N__36701),
            .in2(_gnd_net_),
            .in3(N__36719),
            .lcout(\b2v_inst11.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIED6EB_14_LC_9_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIED6EB_14_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIED6EB_14_LC_9_14_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_off_RNIED6EB_14_LC_9_14_6  (
            .in0(N__31439),
            .in1(N__35891),
            .in2(_gnd_net_),
            .in3(N__31454),
            .lcout(\b2v_inst11.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIEO4AB_5_LC_9_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIEO4AB_5_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIEO4AB_5_LC_9_14_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_off_RNIEO4AB_5_LC_9_14_7  (
            .in0(N__35889),
            .in1(N__36674),
            .in2(_gnd_net_),
            .in3(N__36692),
            .lcout(\b2v_inst11.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_10_LC_9_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_10_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_10_LC_9_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_10_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28369),
            .lcout(\b2v_inst11.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36552),
            .ce(N__28538),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_12_LC_9_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_12_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_12_LC_9_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_12_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28315),
            .lcout(\b2v_inst11.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36552),
            .ce(N__28538),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI111J_7_LC_9_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI111J_7_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI111J_7_LC_9_16_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.count_clk_RNI111J_7_LC_9_16_0  (
            .in0(N__28385),
            .in1(N__28554),
            .in2(N__28397),
            .in3(N__30680),
            .lcout(\b2v_inst11.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_7_LC_9_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_7_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_7_LC_9_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_7_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28393),
            .lcout(\b2v_inst11.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36541),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIEN0E_10_LC_9_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIEN0E_10_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIEN0E_10_LC_9_16_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIEN0E_10_LC_9_16_2  (
            .in0(N__28556),
            .in1(N__28379),
            .in2(N__28373),
            .in3(N__30681),
            .lcout(\b2v_inst11.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIR9EI_13_LC_9_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIR9EI_13_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIR9EI_13_LC_9_16_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIR9EI_13_LC_9_16_3  (
            .in0(N__28598),
            .in1(N__28589),
            .in2(N__30725),
            .in3(N__28558),
            .lcout(\b2v_inst11.count_clkZ0Z_13 ),
            .ltout(\b2v_inst11.count_clkZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_10_LC_9_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_10_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_10_LC_9_16_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNI_10_LC_9_16_4  (
            .in0(N__28297),
            .in1(N__28352),
            .in2(N__28340),
            .in3(N__28336),
            .lcout(\b2v_inst11.un2_count_clk_17_0_o2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIP6DI_12_LC_9_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIP6DI_12_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIP6DI_12_LC_9_16_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIP6DI_12_LC_9_16_5  (
            .in0(N__28316),
            .in1(N__28304),
            .in2(N__30724),
            .in3(N__28557),
            .lcout(\b2v_inst11.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_13_LC_9_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_13_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_13_LC_9_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_13_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28597),
            .lcout(\b2v_inst11.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36541),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_1_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_LC_11_1_0  (
            .in0(_gnd_net_),
            .in1(N__32102),
            .in2(N__32687),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_1_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNID98I1_LC_11_1_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNID98I1_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNID98I1_LC_11_1_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_RNID98I1_LC_11_1_1  (
            .in0(N__32616),
            .in1(N__31574),
            .in2(_gnd_net_),
            .in3(N__28445),
            .lcout(\b2v_inst6.count_rst_12 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_1 ),
            .carryout(\b2v_inst6.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_1_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31615),
            .in3(N__28442),
            .lcout(\b2v_inst6.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_2 ),
            .carryout(\b2v_inst6.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_1_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31495),
            .in3(N__28439),
            .lcout(\b2v_inst6.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_3 ),
            .carryout(\b2v_inst6.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_1_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_1_4  (
            .in0(_gnd_net_),
            .in1(N__32015),
            .in2(_gnd_net_),
            .in3(N__28436),
            .lcout(\b2v_inst6.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_4 ),
            .carryout(\b2v_inst6.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_1_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_1_5  (
            .in0(_gnd_net_),
            .in1(N__28628),
            .in2(_gnd_net_),
            .in3(N__28433),
            .lcout(\b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_5 ),
            .carryout(\b2v_inst6.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_1_6 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_1_6  (
            .in0(_gnd_net_),
            .in1(N__28682),
            .in2(_gnd_net_),
            .in3(N__28430),
            .lcout(\b2v_inst6.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_6 ),
            .carryout(\b2v_inst6.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_1_7 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_1_7  (
            .in0(_gnd_net_),
            .in1(N__32455),
            .in2(_gnd_net_),
            .in3(N__28427),
            .lcout(\b2v_inst6.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_7 ),
            .carryout(\b2v_inst6.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_2_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__29425),
            .in2(_gnd_net_),
            .in3(N__28619),
            .lcout(\b2v_inst6.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNILPGI1_LC_11_2_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNILPGI1_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNILPGI1_LC_11_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_9_c_RNILPGI1_LC_11_2_1  (
            .in0(N__32617),
            .in1(N__28775),
            .in2(_gnd_net_),
            .in3(N__28616),
            .lcout(\b2v_inst6.count_rst_4 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_9 ),
            .carryout(\b2v_inst6.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_2_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_2_2  (
            .in0(_gnd_net_),
            .in1(N__31847),
            .in2(_gnd_net_),
            .in3(N__28613),
            .lcout(\b2v_inst6.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_10 ),
            .carryout(\b2v_inst6.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIU1QP1_LC_11_2_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIU1QP1_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIU1QP1_LC_11_2_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_11_c_RNIU1QP1_LC_11_2_3  (
            .in0(N__32618),
            .in1(N__31754),
            .in2(_gnd_net_),
            .in3(N__28610),
            .lcout(\b2v_inst6.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_11 ),
            .carryout(\b2v_inst6.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNIV3RP1_LC_11_2_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNIV3RP1_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNIV3RP1_LC_11_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_12_c_RNIV3RP1_LC_11_2_4  (
            .in0(N__32620),
            .in1(N__31682),
            .in2(_gnd_net_),
            .in3(N__28607),
            .lcout(\b2v_inst6.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_12 ),
            .carryout(\b2v_inst6.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI06SP1_LC_11_2_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI06SP1_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI06SP1_LC_11_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_13_c_RNI06SP1_LC_11_2_5  (
            .in0(N__32619),
            .in1(N__31787),
            .in2(_gnd_net_),
            .in3(N__28604),
            .lcout(\b2v_inst6.un2_count_1_cry_13_c_RNI06SPZ0Z1 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_13 ),
            .carryout(\b2v_inst6.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNI18TP1_LC_11_2_6 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNI18TP1_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNI18TP1_LC_11_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_14_c_RNI18TP1_LC_11_2_6  (
            .in0(N__32621),
            .in1(N__28691),
            .in2(_gnd_net_),
            .in3(N__28601),
            .lcout(\b2v_inst6.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_10_LC_11_2_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_10_LC_11_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_10_LC_11_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_10_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28794),
            .lcout(\b2v_inst6.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36510),
            .ce(N__32422),
            .sr(N__32651));
    defparam \b2v_inst6.count_15_LC_11_3_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_15_LC_11_3_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_15_LC_11_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_15_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28700),
            .lcout(\b2v_inst6.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36556),
            .ce(N__32429),
            .sr(N__32607));
    defparam \b2v_inst6.count_13_LC_11_3_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_13_LC_11_3_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_13_LC_11_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_13_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31712),
            .lcout(\b2v_inst6.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36556),
            .ce(N__32429),
            .sr(N__32607));
    defparam \b2v_inst6.count_RNIT5A54_15_LC_11_3_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIT5A54_15_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIT5A54_15_LC_11_3_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst6.count_RNIT5A54_15_LC_11_3_2  (
            .in0(N__32361),
            .in1(N__28706),
            .in2(_gnd_net_),
            .in3(N__28699),
            .lcout(\b2v_inst6.countZ0Z_15 ),
            .ltout(\b2v_inst6.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIPV754_0_13_LC_11_3_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIPV754_0_13_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIPV754_0_13_LC_11_3_3 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \b2v_inst6.count_RNIPV754_0_13_LC_11_3_3  (
            .in0(N__31696),
            .in1(N__32362),
            .in2(N__28685),
            .in3(N__31711),
            .lcout(\b2v_inst6.count_1_i_a3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_7_LC_11_3_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_7_LC_11_3_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_7_LC_11_3_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.count_7_LC_11_3_4  (
            .in0(N__28681),
            .in1(N__31942),
            .in2(N__28667),
            .in3(N__32615),
            .lcout(\b2v_inst6.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36556),
            .ce(N__32429),
            .sr(N__32607));
    defparam \b2v_inst6.count_RNIV0AS3_7_LC_11_3_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIV0AS3_7_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIV0AS3_7_LC_11_3_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst6.count_RNIV0AS3_7_LC_11_3_5  (
            .in0(N__28642),
            .in1(N__32360),
            .in2(_gnd_net_),
            .in3(N__28649),
            .lcout(\b2v_inst6.un2_count_1_axb_7 ),
            .ltout(\b2v_inst6.un2_count_1_axb_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIIJDI1_LC_11_3_6 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIIJDI1_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIIJDI1_LC_11_3_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_c_RNIIJDI1_LC_11_3_6  (
            .in0(N__28663),
            .in1(N__31941),
            .in2(N__28652),
            .in3(N__32614),
            .lcout(\b2v_inst6.count_rst_7 ),
            .ltout(\b2v_inst6.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIV0AS3_0_7_LC_11_3_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIV0AS3_0_7_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIV0AS3_0_7_LC_11_3_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \b2v_inst6.count_RNIV0AS3_0_7_LC_11_3_7  (
            .in0(N__28643),
            .in1(N__32363),
            .in2(N__28634),
            .in3(N__32014),
            .lcout(\b2v_inst6.count_1_i_a3_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIALQ32_1_LC_11_4_0 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIALQ32_1_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIALQ32_1_LC_11_4_0 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \b2v_inst6.curr_state_RNIALQ32_1_LC_11_4_0  (
            .in0(N__29729),
            .in1(N__32547),
            .in2(_gnd_net_),
            .in3(N__31209),
            .lcout(\b2v_inst6.count_en ),
            .ltout(\b2v_inst6.count_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNITT8S3_6_LC_11_4_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITT8S3_6_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITT8S3_6_LC_11_4_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \b2v_inst6.count_RNITT8S3_6_LC_11_4_1  (
            .in0(N__32548),
            .in1(N__31655),
            .in2(N__28631),
            .in3(N__31672),
            .lcout(\b2v_inst6.countZ0Z_6 ),
            .ltout(\b2v_inst6.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNICITT3_0_10_LC_11_4_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNICITT3_0_10_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNICITT3_0_10_LC_11_4_2 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \b2v_inst6.count_RNICITT3_0_10_LC_11_4_2  (
            .in0(N__32367),
            .in1(N__28796),
            .in2(N__29348),
            .in3(N__28808),
            .lcout(),
            .ltout(\b2v_inst6.count_1_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI3F438_12_LC_11_4_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI3F438_12_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI3F438_12_LC_11_4_3 .LUT_INIT=16'b0101000000110000;
    LogicCell40 \b2v_inst6.count_RNI3F438_12_LC_11_4_3  (
            .in0(N__31748),
            .in1(N__31730),
            .in2(N__29345),
            .in3(N__32368),
            .lcout(\b2v_inst6.count_1_i_a3_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNINSDS_0_LC_11_4_4 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNINSDS_0_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNINSDS_0_LC_11_4_4 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \b2v_inst36.curr_state_RNINSDS_0_LC_11_4_4  (
            .in0(N__29341),
            .in1(N__29292),
            .in2(N__29243),
            .in3(N__31210),
            .lcout(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ),
            .ltout(\b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIR03I1_9_LC_11_4_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIR03I1_9_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIR03I1_9_LC_11_4_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \b2v_inst36.count_RNIR03I1_9_LC_11_4_5  (
            .in0(_gnd_net_),
            .in1(N__29168),
            .in2(N__29192),
            .in3(N__29156),
            .lcout(\b2v_inst36.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_9_LC_11_4_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_9_LC_11_4_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_9_LC_11_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_9_LC_11_4_6  (
            .in0(N__29167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36402),
            .ce(N__29126),
            .sr(N__28972));
    defparam \b2v_inst6.count_RNICITT3_10_LC_11_4_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNICITT3_10_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNICITT3_10_LC_11_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNICITT3_10_LC_11_4_7  (
            .in0(N__28807),
            .in1(N__28795),
            .in2(_gnd_net_),
            .in3(N__32366),
            .lcout(\b2v_inst6.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_11_5_0 .C_ON=1'b0;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_11_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.un8_rsmrst_pwrgd_4_LC_11_5_0  (
            .in0(N__28766),
            .in1(N__28751),
            .in2(N__28739),
            .in3(N__28718),
            .lcout(SYNTHESIZED_WIRE_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIKNFI1_LC_11_5_2 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIKNFI1_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIKNFI1_LC_11_5_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_c_RNIKNFI1_LC_11_5_2  (
            .in0(N__32542),
            .in1(N__29407),
            .in2(N__29426),
            .in3(N__31954),
            .lcout(\b2v_inst6.count_rst_5 ),
            .ltout(\b2v_inst6.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI37CS3_9_LC_11_5_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI37CS3_9_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI37CS3_9_LC_11_5_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNI37CS3_9_LC_11_5_3  (
            .in0(N__32365),
            .in1(_gnd_net_),
            .in2(N__28709),
            .in3(N__32467),
            .lcout(\b2v_inst6.un2_count_1_axb_9 ),
            .ltout(\b2v_inst6.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_9_LC_11_5_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_9_LC_11_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_9_LC_11_5_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.count_9_LC_11_5_4  (
            .in0(N__32649),
            .in1(N__29408),
            .in2(N__29396),
            .in3(N__31955),
            .lcout(\b2v_inst6.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36568),
            .ce(N__32428),
            .sr(N__32648));
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNIJLEI1_LC_11_5_5 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNIJLEI1_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNIJLEI1_LC_11_5_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_c_RNIJLEI1_LC_11_5_5  (
            .in0(N__32451),
            .in1(N__31952),
            .in2(N__29390),
            .in3(N__32541),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI14BS3_8_LC_11_5_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI14BS3_8_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI14BS3_8_LC_11_5_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst6.count_RNI14BS3_8_LC_11_5_6  (
            .in0(N__29372),
            .in1(_gnd_net_),
            .in2(N__29393),
            .in3(N__32364),
            .lcout(\b2v_inst6.countZ0Z_8 ),
            .ltout(\b2v_inst6.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_8_LC_11_5_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_8_LC_11_5_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_8_LC_11_5_7 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.count_8_LC_11_5_7  (
            .in0(N__29389),
            .in1(N__31953),
            .in2(N__29375),
            .in3(N__32543),
            .lcout(\b2v_inst6.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36568),
            .ce(N__32428),
            .sr(N__32648));
    defparam \b2v_inst6.curr_state_1_LC_11_6_0 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_1_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_1_LC_11_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.curr_state_1_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29354),
            .lcout(\b2v_inst6.curr_state_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36635),
            .ce(N__32183),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_0_LC_11_6_1 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_0_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_0_LC_11_6_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \b2v_inst6.curr_state_0_LC_11_6_1  (
            .in0(N__31951),
            .in1(N__29514),
            .in2(N__29704),
            .in3(N__29537),
            .lcout(\b2v_inst6.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36635),
            .ce(N__32183),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_11_6_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_11_6_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m4_0_LC_11_6_2  (
            .in0(N__29515),
            .in1(N__29535),
            .in2(N__29705),
            .in3(N__31949),
            .lcout(),
            .ltout(\b2v_inst6.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI5DHS1_0_LC_11_6_3 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI5DHS1_0_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI5DHS1_0_LC_11_6_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.curr_state_RNI5DHS1_0_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__29363),
            .in2(N__29357),
            .in3(N__30597),
            .lcout(\b2v_inst6.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_LC_11_6_4 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_LC_11_6_4 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m6_i_LC_11_6_4  (
            .in0(N__29536),
            .in1(N__31950),
            .in2(_gnd_net_),
            .in3(N__29725),
            .lcout(\b2v_inst6.N_42 ),
            .ltout(\b2v_inst6.N_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI8KCH_1_LC_11_6_5 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI8KCH_1_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI8KCH_1_LC_11_6_5 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \b2v_inst6.curr_state_RNI8KCH_1_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__29546),
            .in2(N__29540),
            .in3(N__30595),
            .lcout(\b2v_inst6.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst6.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI_1_LC_11_6_6 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI_1_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI_1_LC_11_6_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst6.curr_state_RNI_1_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29522),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.N_3053_i ),
            .ltout(\b2v_inst6.N_3053_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIM6FE1_1_LC_11_6_7 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIM6FE1_1_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIM6FE1_1_LC_11_6_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIM6FE1_1_LC_11_6_7  (
            .in0(N__29516),
            .in1(N__29756),
            .in2(N__29519),
            .in3(N__30596),
            .lcout(\b2v_inst6.curr_state_RNIM6FE1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI_0_LC_11_7_1 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI_0_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI_0_LC_11_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.curr_state_RNI_0_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29451),
            .lcout(\b2v_inst6.N_3034_i ),
            .ltout(\b2v_inst6.N_3034_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIUP4B1_1_LC_11_7_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIUP4B1_1_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIUP4B1_1_LC_11_7_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIUP4B1_1_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__29436),
            .in2(N__29501),
            .in3(N__29754),
            .lcout(\b2v_inst6.N_276_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIUP4B1_0_LC_11_7_3 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIUP4B1_0_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIUP4B1_0_LC_11_7_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIUP4B1_0_LC_11_7_3  (
            .in0(N__29755),
            .in1(_gnd_net_),
            .in2(N__29441),
            .in3(N__29452),
            .lcout(\b2v_inst6.curr_state_RNIUP4B1Z0Z_0 ),
            .ltout(\b2v_inst6.curr_state_RNIUP4B1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU8MF3_LC_11_7_4 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU8MF3_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU8MF3_LC_11_7_4 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU8MF3_LC_11_7_4  (
            .in0(N__29680),
            .in1(N__29713),
            .in2(N__29498),
            .in3(N__32215),
            .lcout(),
            .ltout(\b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_LC_11_7_5 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_LC_11_7_5 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIIJ994_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29495),
            .in3(N__34927),
            .lcout(N_222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_7_6 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_7_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_7_6  (
            .in0(N__29453),
            .in1(N__29440),
            .in2(_gnd_net_),
            .in3(N__29753),
            .lcout(N_241),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_7_7 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_7_7 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_7_7  (
            .in0(N__29714),
            .in1(N__29697),
            .in2(N__32225),
            .in3(N__29681),
            .lcout(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36449),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_LC_11_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_LC_11_8_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst11.func_state_RNI_1_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__34061),
            .in2(_gnd_net_),
            .in3(N__35109),
            .lcout(\b2v_inst11.N_172 ),
            .ltout(\b2v_inst11.N_172_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_3_LC_11_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_3_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_3_LC_11_8_1 .LUT_INIT=16'b1010100000001010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_3_LC_11_8_1  (
            .in0(N__33078),
            .in1(N__29672),
            .in2(N__29657),
            .in3(N__33311),
            .lcout(),
            .ltout(\b2v_inst11.g0_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIKAJP_6_LC_11_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIKAJP_6_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIKAJP_6_LC_11_8_2 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIKAJP_6_LC_11_8_2  (
            .in0(N__29654),
            .in1(N__33377),
            .in2(N__29642),
            .in3(N__34919),
            .lcout(\b2v_inst11.g0_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINGLA1_1_LC_11_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINGLA1_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINGLA1_1_LC_11_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.func_state_RNINGLA1_1_LC_11_8_3  (
            .in0(N__35110),
            .in1(N__30047),
            .in2(N__30326),
            .in3(N__29636),
            .lcout(),
            .ltout(\b2v_inst11.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI4KE12_LC_11_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI4KE12_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI4KE12_LC_11_8_4 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI4KE12_LC_11_8_4  (
            .in0(N__29585),
            .in1(N__34495),
            .in2(N__29573),
            .in3(N__35111),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_11_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_11_8_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__32896),
            .in2(_gnd_net_),
            .in3(N__34494),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_0_o3_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_11_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_11_8_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_0_LC_11_8_6  (
            .in0(N__29561),
            .in1(N__31332),
            .in2(N__33314),
            .in3(N__30143),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.N_224_i_LC_11_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.N_224_i_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.N_224_i_LC_11_8_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.N_224_i_LC_11_8_7  (
            .in0(N__34421),
            .in1(N__34241),
            .in2(N__30325),
            .in3(N__30598),
            .lcout(\b2v_inst11.N_224_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI34G9_0_LC_11_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI34G9_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI34G9_0_LC_11_9_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.func_state_RNI34G9_0_LC_11_9_2  (
            .in0(N__34422),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34064),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNII5M67_2_LC_11_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNII5M67_2_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNII5M67_2_LC_11_9_3 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \b2v_inst11.dutycycle_RNII5M67_2_LC_11_9_3  (
            .in0(N__29980),
            .in1(N__30007),
            .in2(N__30020),
            .in3(N__29995),
            .lcout(\b2v_inst11.dutycycleZ0Z_2 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_11_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_11_9_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30041),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_2_LC_11_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_2_LC_11_9_5 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_2_LC_11_9_5 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \b2v_inst11.dutycycle_2_LC_11_9_5  (
            .in0(N__30019),
            .in1(N__30008),
            .in2(N__29984),
            .in3(N__29996),
            .lcout(\b2v_inst11.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36207),
            .ce(),
            .sr(N__30984));
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_11_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_11_10_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_0_LC_11_10_1  (
            .in0(N__29962),
            .in1(N__29809),
            .in2(N__30166),
            .in3(N__31310),
            .lcout(\b2v_inst11.N_293_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_11_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_11_10_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_0_LC_11_10_2  (
            .in0(N__31311),
            .in1(N__29963),
            .in2(N__29813),
            .in3(N__30142),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_2_1_LC_11_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_11_10_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst11.func_state_RNI_2_1_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__34059),
            .in2(_gnd_net_),
            .in3(N__35091),
            .lcout(\b2v_inst11.func_state_RNI_2Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNI_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIN1E71_1_LC_11_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIN1E71_1_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIN1E71_1_LC_11_10_4 .LUT_INIT=16'b1111111100110001;
    LogicCell40 \b2v_inst11.func_state_RNIN1E71_1_LC_11_10_4  (
            .in0(N__32895),
            .in1(N__34931),
            .in2(N__29771),
            .in3(N__29768),
            .lcout(\b2v_inst11.N_119_f0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_LC_11_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_LC_11_10_5 .LUT_INIT=16'b1000000010010001;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_1_LC_11_10_5  (
            .in0(N__35583),
            .in1(N__34060),
            .in2(N__30785),
            .in3(N__35093),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_ss0_i_0_o3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIHVOG4_0_1_LC_11_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIHVOG4_0_1_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIHVOG4_0_1_LC_11_10_6 .LUT_INIT=16'b1111110111111101;
    LogicCell40 \b2v_inst11.func_state_RNIHVOG4_0_1_LC_11_10_6  (
            .in0(N__34810),
            .in1(N__30230),
            .in2(N__30764),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI57FD1_1_LC_11_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI57FD1_1_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI57FD1_1_LC_11_10_7 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \b2v_inst11.func_state_RNI57FD1_1_LC_11_10_7  (
            .in0(N__34250),
            .in1(N__35092),
            .in2(N__30705),
            .in3(N__30324),
            .lcout(\b2v_inst11.N_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIN52J1_LC_11_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIN52J1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIN52J1_LC_11_11_0 .LUT_INIT=16'b1111101111110001;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIN52J1_LC_11_11_0  (
            .in0(N__35105),
            .in1(N__30224),
            .in2(N__33515),
            .in3(N__30898),
            .lcout(\b2v_inst11.dutycycle_1_0_1 ),
            .ltout(\b2v_inst11.dutycycle_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIB6O76_1_LC_11_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIB6O76_1_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIB6O76_1_LC_11_11_1 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIB6O76_1_LC_11_11_1  (
            .in0(N__31236),
            .in1(N__31051),
            .in2(N__30209),
            .in3(N__31256),
            .lcout(\b2v_inst11.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_0_LC_11_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_0_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_0_LC_11_11_2 .LUT_INIT=16'b0111000011111000;
    LogicCell40 \b2v_inst11.dutycycle_0_LC_11_11_2  (
            .in0(N__30206),
            .in1(N__31238),
            .in2(N__30200),
            .in3(N__30056),
            .lcout(\b2v_inst11.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36416),
            .ce(),
            .sr(N__31036));
    defparam \b2v_inst11.dutycycle_RNIAA6Q3_0_LC_11_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAA6Q3_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAA6Q3_0_LC_11_11_3 .LUT_INIT=16'b0101010111111101;
    LogicCell40 \b2v_inst11.dutycycle_RNIAA6Q3_0_LC_11_11_3  (
            .in0(N__34808),
            .in1(N__30115),
            .in2(N__34938),
            .in3(N__31387),
            .lcout(\b2v_inst11.dutycycle_eena ),
            .ltout(\b2v_inst11.dutycycle_eena_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI0QQU5_0_LC_11_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI0QQU5_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI0QQU5_0_LC_11_11_4 .LUT_INIT=16'b0010101011101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI0QQU5_0_LC_11_11_4  (
            .in0(N__30196),
            .in1(N__31235),
            .in2(N__30188),
            .in3(N__30055),
            .lcout(\b2v_inst11.dutycycleZ0Z_0 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_LC_11_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_LC_11_11_5 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_0_LC_11_11_5  (
            .in0(N__30897),
            .in1(N__33509),
            .in2(N__30059),
            .in3(N__35104),
            .lcout(\b2v_inst11.dutycycle_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAA6Q3_1_LC_11_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAA6Q3_1_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAA6Q3_1_LC_11_11_6 .LUT_INIT=16'b0011111100111011;
    LogicCell40 \b2v_inst11.dutycycle_RNIAA6Q3_1_LC_11_11_6  (
            .in0(N__34926),
            .in1(N__34809),
            .in2(N__31391),
            .in3(N__31309),
            .lcout(\b2v_inst11.dutycycle_eena_0 ),
            .ltout(\b2v_inst11.dutycycle_eena_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_LC_11_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_1_LC_11_11_7 .LUT_INIT=16'b0111111100100000;
    LogicCell40 \b2v_inst11.dutycycle_1_LC_11_11_7  (
            .in0(N__31237),
            .in1(N__31061),
            .in2(N__31055),
            .in3(N__31052),
            .lcout(\b2v_inst11.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36416),
            .ce(),
            .sr(N__31036));
    defparam \b2v_inst11.count_off_RNIL5413_0_LC_11_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIL5413_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIL5413_0_LC_11_12_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.count_off_RNIL5413_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__35326),
            .in2(_gnd_net_),
            .in3(N__35271),
            .lcout(),
            .ltout(\b2v_inst11.count_off_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI8BS7B_0_LC_11_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI8BS7B_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI8BS7B_0_LC_11_12_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_off_RNI8BS7B_0_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__35231),
            .in2(N__30917),
            .in3(N__35929),
            .lcout(\b2v_inst11.count_offZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_11_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_11_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_11_12_2  (
            .in0(N__30848),
            .in1(N__31420),
            .in2(_gnd_net_),
            .in3(N__30827),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_330_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_0_LC_11_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_11_12_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.func_state_RNI_0_0_LC_11_12_3  (
            .in0(N__35106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30902),
            .lcout(\b2v_inst11.func_state_RNI_0Z0Z_0 ),
            .ltout(\b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8BVM1_0_LC_11_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8BVM1_0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8BVM1_0_LC_11_12_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.func_state_RNI8BVM1_0_LC_11_12_4  (
            .in0(N__30842),
            .in1(N__30826),
            .in2(N__30803),
            .in3(N__35577),
            .lcout(),
            .ltout(\b2v_inst11.N_315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIL5413_1_LC_11_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIL5413_1_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIL5413_1_LC_11_12_5 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \b2v_inst11.func_state_RNIL5413_1_LC_11_12_5  (
            .in0(N__35107),
            .in1(N__35587),
            .in2(N__30800),
            .in3(N__30797),
            .lcout(\b2v_inst11.N_125 ),
            .ltout(\b2v_inst11.N_125_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIL5413_1_LC_11_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIL5413_1_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIL5413_1_LC_11_12_6 .LUT_INIT=16'b0011000011000000;
    LogicCell40 \b2v_inst11.count_off_RNIL5413_1_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__35362),
            .in2(N__31430),
            .in3(N__35325),
            .lcout(\b2v_inst11.count_off_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_11_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_11_12_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_11_12_7  (
            .in0(N__34493),
            .in1(N__32894),
            .in2(N__34445),
            .in3(N__34301),
            .lcout(\b2v_inst11.N_382_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_11_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__35327),
            .in2(N__35363),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIJ7933_LC_11_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIJ7933_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIJ7933_LC_11_13_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_RNIJ7933_LC_11_13_1  (
            .in0(N__35272),
            .in1(N__35626),
            .in2(_gnd_net_),
            .in3(N__31409),
            .lcout(\b2v_inst11.count_off_1_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_1 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIK9A33_LC_11_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIK9A33_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIK9A33_LC_11_13_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_2_c_RNIK9A33_LC_11_13_2  (
            .in0(N__35276),
            .in1(N__35416),
            .in2(_gnd_net_),
            .in3(N__31406),
            .lcout(\b2v_inst11.count_off_1_3 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_2 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNILBB33_LC_11_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNILBB33_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNILBB33_LC_11_13_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_3_c_RNILBB33_LC_11_13_3  (
            .in0(N__35273),
            .in1(N__35392),
            .in2(_gnd_net_),
            .in3(N__31403),
            .lcout(\b2v_inst11.count_off_1_4 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_3 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNIMDC33_LC_11_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNIMDC33_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNIMDC33_LC_11_13_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_4_c_RNIMDC33_LC_11_13_4  (
            .in0(N__35277),
            .in1(N__35653),
            .in2(_gnd_net_),
            .in3(N__31400),
            .lcout(\b2v_inst11.count_off_1_5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_4 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNINFD33_LC_11_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNINFD33_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNINFD33_LC_11_13_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_5_c_RNINFD33_LC_11_13_5  (
            .in0(N__35274),
            .in1(N__35671),
            .in2(_gnd_net_),
            .in3(N__31397),
            .lcout(\b2v_inst11.count_off_1_6 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_5 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIOHE33_LC_11_13_6 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIOHE33_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIOHE33_LC_11_13_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_6_c_RNIOHE33_LC_11_13_6  (
            .in0(N__35278),
            .in1(N__35458),
            .in2(_gnd_net_),
            .in3(N__31394),
            .lcout(\b2v_inst11.count_off_1_7 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_6 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNIPJF33_LC_11_13_7 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNIPJF33_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNIPJF33_LC_11_13_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_7_c_RNIPJF33_LC_11_13_7  (
            .in0(N__35275),
            .in1(N__35437),
            .in2(_gnd_net_),
            .in3(N__31478),
            .lcout(\b2v_inst11.count_off_1_8 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_7 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIQLG33_LC_11_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIQLG33_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIQLG33_LC_11_14_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_8_c_RNIQLG33_LC_11_14_0  (
            .in0(N__35297),
            .in1(N__35210),
            .in2(_gnd_net_),
            .in3(N__31475),
            .lcout(\b2v_inst11.count_off_1_9 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNIRNH33_LC_11_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNIRNH33_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNIRNH33_LC_11_14_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_9_c_RNIRNH33_LC_11_14_1  (
            .in0(N__35301),
            .in1(_gnd_net_),
            .in2(N__35813),
            .in3(N__31472),
            .lcout(\b2v_inst11.count_off_1_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_9 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI35P63_LC_11_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI35P63_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI35P63_LC_11_14_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_10_c_RNI35P63_LC_11_14_2  (
            .in0(N__35298),
            .in1(N__35782),
            .in2(_gnd_net_),
            .in3(N__31469),
            .lcout(\b2v_inst11.count_off_1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_10 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNI47Q63_LC_11_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNI47Q63_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNI47Q63_LC_11_14_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_11_c_RNI47Q63_LC_11_14_3  (
            .in0(N__35303),
            .in1(N__35756),
            .in2(_gnd_net_),
            .in3(N__31466),
            .lcout(\b2v_inst11.count_off_1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_11 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNI59R63_LC_11_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNI59R63_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNI59R63_LC_11_14_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_12_c_RNI59R63_LC_11_14_4  (
            .in0(N__35299),
            .in1(N__35506),
            .in2(_gnd_net_),
            .in3(N__31463),
            .lcout(\b2v_inst11.count_off_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_12 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNI6BS63_LC_11_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNI6BS63_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNI6BS63_LC_11_14_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_13_c_RNI6BS63_LC_11_14_5  (
            .in0(N__35302),
            .in1(N__35482),
            .in2(_gnd_net_),
            .in3(N__31460),
            .lcout(\b2v_inst11.count_off_1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_13 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DT63_LC_11_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DT63_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DT63_LC_11_14_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_14_c_RNI7DT63_LC_11_14_6  (
            .in0(N__35300),
            .in1(N__35524),
            .in2(_gnd_net_),
            .in3(N__31457),
            .lcout(\b2v_inst11.un3_count_off_1_cry_14_c_RNI7DTZ0Z63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_14_LC_11_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_14_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_14_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_off_14_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31453),
            .lcout(\b2v_inst11.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36618),
            .ce(N__35941),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIGG7EB_15_LC_11_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIGG7EB_15_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIGG7EB_15_LC_11_15_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_off_RNIGG7EB_15_LC_11_15_0  (
            .in0(N__31568),
            .in1(N__31559),
            .in2(_gnd_net_),
            .in3(N__35937),
            .lcout(\b2v_inst11.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_15_LC_11_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_15_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_15_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_off_15_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31567),
            .lcout(\b2v_inst11.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36489),
            .ce(N__35942),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIGR5AB_6_LC_11_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIGR5AB_6_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIGR5AB_6_LC_11_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_off_RNIGR5AB_6_LC_11_15_2  (
            .in0(N__31541),
            .in1(N__31552),
            .in2(_gnd_net_),
            .in3(N__35934),
            .lcout(\b2v_inst11.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_6_LC_11_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_6_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_6_LC_11_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_off_6_LC_11_15_3  (
            .in0(N__31553),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36489),
            .ce(N__35942),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIIU6AB_7_LC_11_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIIU6AB_7_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIIU6AB_7_LC_11_15_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_off_RNIIU6AB_7_LC_11_15_4  (
            .in0(N__31523),
            .in1(N__31534),
            .in2(_gnd_net_),
            .in3(N__35935),
            .lcout(\b2v_inst11.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_7_LC_11_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_7_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_7_LC_11_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_off_7_LC_11_15_5  (
            .in0(N__31535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36489),
            .ce(N__35942),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIK18AB_8_LC_11_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIK18AB_8_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIK18AB_8_LC_11_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_off_RNIK18AB_8_LC_11_15_6  (
            .in0(N__31505),
            .in1(N__31516),
            .in2(_gnd_net_),
            .in3(N__35936),
            .lcout(\b2v_inst11.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_8_LC_11_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_8_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_8_LC_11_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_off_8_LC_11_15_7  (
            .in0(N__31517),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36489),
            .ce(N__35942),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIFDAI1_LC_12_1_0 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIFDAI1_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIFDAI1_LC_12_1_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_c_RNIFDAI1_LC_12_1_0  (
            .in0(N__31945),
            .in1(N__31645),
            .in2(N__31496),
            .in3(N__32623),
            .lcout(\b2v_inst6.count_rst_10 ),
            .ltout(\b2v_inst6.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIPN6S3_4_LC_12_1_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIPN6S3_4_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIPN6S3_4_LC_12_1_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNIPN6S3_4_LC_12_1_1  (
            .in0(_gnd_net_),
            .in1(N__31627),
            .in2(N__31499),
            .in3(N__32397),
            .lcout(\b2v_inst6.un2_count_1_axb_4 ),
            .ltout(\b2v_inst6.un2_count_1_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_4_LC_12_1_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_4_LC_12_1_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_4_LC_12_1_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.count_4_LC_12_1_2  (
            .in0(N__31947),
            .in1(N__31646),
            .in2(N__31637),
            .in3(N__32626),
            .lcout(\b2v_inst6.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36349),
            .ce(N__32432),
            .sr(N__32635));
    defparam \b2v_inst6.count_RNIPN6S3_0_4_LC_12_1_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIPN6S3_0_4_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIPN6S3_0_4_LC_12_1_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \b2v_inst6.count_RNIPN6S3_0_4_LC_12_1_3  (
            .in0(N__31611),
            .in1(N__31634),
            .in2(N__32431),
            .in3(N__31628),
            .lcout(\b2v_inst6.count_1_i_a3_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIEB9I1_LC_12_1_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIEB9I1_LC_12_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIEB9I1_LC_12_1_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_c_RNIEB9I1_LC_12_1_4  (
            .in0(N__31944),
            .in1(N__31591),
            .in2(N__31616),
            .in3(N__32622),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNINK5S3_3_LC_12_1_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNINK5S3_3_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNINK5S3_3_LC_12_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNINK5S3_3_LC_12_1_5  (
            .in0(_gnd_net_),
            .in1(N__31580),
            .in2(N__31619),
            .in3(N__32396),
            .lcout(\b2v_inst6.countZ0Z_3 ),
            .ltout(\b2v_inst6.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_3_LC_12_1_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_3_LC_12_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_3_LC_12_1_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.count_3_LC_12_1_6  (
            .in0(N__31946),
            .in1(N__31592),
            .in2(N__31583),
            .in3(N__32625),
            .lcout(\b2v_inst6.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36349),
            .ce(N__32432),
            .sr(N__32635));
    defparam \b2v_inst6.count_11_LC_12_1_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_11_LC_12_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_11_LC_12_1_7 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.count_11_LC_12_1_7  (
            .in0(N__32624),
            .in1(N__31855),
            .in2(N__31973),
            .in3(N__31948),
            .lcout(\b2v_inst6.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36349),
            .ce(N__32432),
            .sr(N__32635));
    defparam \b2v_inst6.count_14_LC_12_2_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_14_LC_12_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_14_LC_12_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_14_LC_12_2_0  (
            .in0(N__31796),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36530),
            .ce(N__32430),
            .sr(N__32650));
    defparam \b2v_inst6.count_RNILH4S3_2_LC_12_2_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNILH4S3_2_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNILH4S3_2_LC_12_2_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst6.count_RNILH4S3_2_LC_12_2_1  (
            .in0(N__31764),
            .in1(N__31780),
            .in2(_gnd_net_),
            .in3(N__32373),
            .lcout(\b2v_inst6.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_2_LC_12_2_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_2_LC_12_2_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_2_LC_12_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_2_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31766),
            .lcout(\b2v_inst6.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36530),
            .ce(N__32430),
            .sr(N__32650));
    defparam \b2v_inst6.count_RNIR2954_14_LC_12_2_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIR2954_14_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIR2954_14_LC_12_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIR2954_14_LC_12_2_3  (
            .in0(N__31802),
            .in1(N__31795),
            .in2(_gnd_net_),
            .in3(N__32376),
            .lcout(\b2v_inst6.countZ0Z_14 ),
            .ltout(\b2v_inst6.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNILH4S3_0_2_LC_12_2_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNILH4S3_0_2_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNILH4S3_0_2_LC_12_2_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \b2v_inst6.count_RNILH4S3_0_2_LC_12_2_4  (
            .in0(N__32377),
            .in1(N__31781),
            .in2(N__31769),
            .in3(N__31765),
            .lcout(\b2v_inst6.count_1_i_a3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNINS654_12_LC_12_2_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNINS654_12_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNINS654_12_LC_12_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNINS654_12_LC_12_2_5  (
            .in0(N__31723),
            .in1(N__31743),
            .in2(_gnd_net_),
            .in3(N__32374),
            .lcout(\b2v_inst6.un2_count_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_12_LC_12_2_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_12_LC_12_2_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_12_LC_12_2_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_12_LC_12_2_6  (
            .in0(N__31744),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36530),
            .ce(N__32430),
            .sr(N__32650));
    defparam \b2v_inst6.count_RNIPV754_13_LC_12_2_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIPV754_13_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIPV754_13_LC_12_2_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst6.count_RNIPV754_13_LC_12_2_7  (
            .in0(N__31710),
            .in1(N__31697),
            .in2(_gnd_net_),
            .in3(N__32375),
            .lcout(\b2v_inst6.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_6_LC_12_3_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_6_LC_12_3_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_6_LC_12_3_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst6.count_6_LC_12_3_0  (
            .in0(N__32611),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31676),
            .lcout(\b2v_inst6.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36367),
            .ce(N__32427),
            .sr(N__32613));
    defparam \b2v_inst6.count_RNI_0_0_LC_12_3_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_0_0_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_0_0_LC_12_3_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst6.count_RNI_0_0_LC_12_3_1  (
            .in0(N__32711),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32076),
            .lcout(\b2v_inst6.N_394 ),
            .ltout(\b2v_inst6.N_394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIGFBI1_LC_12_3_2 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIGFBI1_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIGFBI1_LC_12_3_2 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_c_RNIGFBI1_LC_12_3_2  (
            .in0(N__32609),
            .in1(N__31993),
            .in2(N__31649),
            .in3(N__32013),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIRQ7S3_5_LC_12_3_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRQ7S3_5_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRQ7S3_5_LC_12_3_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNIRQ7S3_5_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__31979),
            .in2(N__32018),
            .in3(N__32358),
            .lcout(\b2v_inst6.countZ0Z_5 ),
            .ltout(\b2v_inst6.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_5_LC_12_3_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_5_LC_12_3_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_5_LC_12_3_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.count_5_LC_12_3_4  (
            .in0(N__32612),
            .in1(N__31994),
            .in2(N__31982),
            .in3(N__31923),
            .lcout(\b2v_inst6.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36367),
            .ce(N__32427),
            .sr(N__32613));
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNITVOP1_LC_12_3_5 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNITVOP1_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNITVOP1_LC_12_3_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_c_RNITVOP1_LC_12_3_5  (
            .in0(N__31966),
            .in1(N__31943),
            .in2(N__31856),
            .in3(N__32610),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNILP554_11_LC_12_3_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNILP554_11_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNILP554_11_LC_12_3_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNILP554_11_LC_12_3_6  (
            .in0(N__32359),
            .in1(_gnd_net_),
            .in2(N__31877),
            .in3(N__31874),
            .lcout(\b2v_inst6.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIM6FE1_0_LC_12_3_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIM6FE1_0_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIM6FE1_0_LC_12_3_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst6.count_RNIM6FE1_0_LC_12_3_7  (
            .in0(N__32710),
            .in1(N__32077),
            .in2(_gnd_net_),
            .in3(N__32608),
            .lcout(\b2v_inst6.count_RNIM6FE1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNISCBO3_0_LC_12_4_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNISCBO3_0_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNISCBO3_0_LC_12_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNISCBO3_0_LC_12_4_0  (
            .in0(N__32699),
            .in1(N__31865),
            .in2(_gnd_net_),
            .in3(N__32331),
            .lcout(\b2v_inst6.countZ0Z_0 ),
            .ltout(\b2v_inst6.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIM6FE1_1_LC_12_4_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIM6FE1_1_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIM6FE1_1_LC_12_4_1 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \b2v_inst6.count_RNIM6FE1_1_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(N__32680),
            .in2(N__31859),
            .in3(N__32582),
            .lcout(\b2v_inst6.count_rst_13 ),
            .ltout(\b2v_inst6.count_rst_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNITDBO3_0_1_LC_12_4_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITDBO3_0_1_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITDBO3_0_1_LC_12_4_2 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \b2v_inst6.count_RNITDBO3_0_1_LC_12_4_2  (
            .in0(N__31854),
            .in1(N__32662),
            .in2(N__31826),
            .in3(N__32330),
            .lcout(),
            .ltout(\b2v_inst6.count_1_i_a3_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIOD8DF_1_LC_12_4_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIOD8DF_1_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIOD8DF_1_LC_12_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNIOD8DF_1_LC_12_4_3  (
            .in0(N__31823),
            .in1(N__31814),
            .in2(N__31805),
            .in3(N__32264),
            .lcout(),
            .ltout(\b2v_inst6.count_1_i_a3_12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI9EPHV_2_LC_12_4_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI9EPHV_2_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI9EPHV_2_LC_12_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNI9EPHV_2_LC_12_4_4  (
            .in0(N__32735),
            .in1(N__32729),
            .in2(N__32720),
            .in3(N__32717),
            .lcout(\b2v_inst6.N_389 ),
            .ltout(\b2v_inst6.N_389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_0_LC_12_4_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_0_LC_12_4_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_0_LC_12_4_5 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \b2v_inst6.count_0_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(N__32078),
            .in2(N__32702),
            .in3(N__32583),
            .lcout(\b2v_inst6.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36480),
            .ce(N__32423),
            .sr(N__32641));
    defparam \b2v_inst6.count_RNITDBO3_1_LC_12_4_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITDBO3_1_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITDBO3_1_LC_12_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNITDBO3_1_LC_12_4_6  (
            .in0(N__32663),
            .in1(N__32693),
            .in2(_gnd_net_),
            .in3(N__32332),
            .lcout(\b2v_inst6.un2_count_1_axb_1 ),
            .ltout(\b2v_inst6.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_1_LC_12_4_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_1_LC_12_4_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_1_LC_12_4_7 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \b2v_inst6.count_1_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(N__32100),
            .in2(N__32666),
            .in3(N__32584),
            .lcout(\b2v_inst6.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36480),
            .ce(N__32423),
            .sr(N__32641));
    defparam \b2v_inst6.count_RNI37CS3_0_9_LC_12_5_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI37CS3_0_9_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI37CS3_0_9_LC_12_5_0 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \b2v_inst6.count_RNI37CS3_0_9_LC_12_5_0  (
            .in0(N__32474),
            .in1(N__32468),
            .in2(N__32456),
            .in3(N__32372),
            .lcout(\b2v_inst6.count_1_i_a3_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_1_LC_12_6_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_1_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_1_LC_12_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst5.curr_state_1_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32255),
            .lcout(\b2v_inst5.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36598),
            .ce(N__32178),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_0_LC_12_6_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_0_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_0_LC_12_6_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \b2v_inst6.count_RNI_0_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__32101),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.N_3036_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_7_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_7_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_7_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst31.un6_output_LC_12_7_7 .C_ON=1'b0;
    defparam \b2v_inst31.un6_output_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst31.un6_output_LC_12_7_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst31.un6_output_LC_12_7_7  (
            .in0(N__34928),
            .in1(N__33011),
            .in2(N__33005),
            .in3(N__32972),
            .lcout(vccinaux_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_0_LC_12_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_0_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_0_LC_12_8_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_0_LC_12_8_1  (
            .in0(N__33730),
            .in1(N__33312),
            .in2(_gnd_net_),
            .in3(N__32927),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI7FEU3_0_LC_12_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI7FEU3_0_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI7FEU3_0_LC_12_8_2 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI7FEU3_0_LC_12_8_2  (
            .in0(N__33920),
            .in1(N__32750),
            .in2(N__32918),
            .in3(N__34062),
            .lcout(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_rn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GPIO_FPGA_SoC_4_RNI8H551_LC_12_8_3.C_ON=1'b0;
    defparam GPIO_FPGA_SoC_4_RNI8H551_LC_12_8_3.SEQ_MODE=4'b0000;
    defparam GPIO_FPGA_SoC_4_RNI8H551_LC_12_8_3.LUT_INIT=16'b0100010000000000;
    LogicCell40 GPIO_FPGA_SoC_4_RNI8H551_LC_12_8_3 (
            .in0(N__34388),
            .in1(N__32915),
            .in2(_gnd_net_),
            .in3(N__34604),
            .lcout(G_6_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_12_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_12_8_4 .LUT_INIT=16'b0100011111001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_2_LC_12_8_4  (
            .in0(N__33150),
            .in1(N__32762),
            .in2(N__33731),
            .in3(N__34063),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_172_m1_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQK9K2_2_LC_12_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_2_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_2_LC_12_8_5 .LUT_INIT=16'b1110101011100000;
    LogicCell40 \b2v_inst11.dutycycle_RNIQK9K2_2_LC_12_8_5  (
            .in0(N__32761),
            .in1(N__33500),
            .in2(N__32753),
            .in3(N__33921),
            .lcout(\b2v_inst11.un1_dutycycle_172_m1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_5_1_LC_12_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_5_1_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_5_1_LC_12_8_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \b2v_inst11.func_state_RNI_5_1_LC_12_8_7  (
            .in0(N__33378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33313),
            .lcout(\b2v_inst11.N_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.g0_0_0_0_LC_12_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.g0_0_0_0_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.g0_0_0_0_LC_12_9_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.g0_0_0_0_LC_12_9_0  (
            .in0(N__34395),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34603),
            .lcout(),
            .ltout(\b2v_inst11.g0_0_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI0GIO3_6_LC_12_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI0GIO3_6_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI0GIO3_6_LC_12_9_1 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI0GIO3_6_LC_12_9_1  (
            .in0(N__34813),
            .in1(N__32744),
            .in2(N__32738),
            .in3(N__34284),
            .lcout(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_0_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQK9K2_3_LC_12_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_3_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_3_LC_12_9_2 .LUT_INIT=16'b0000110000101110;
    LogicCell40 \b2v_inst11.dutycycle_RNIQK9K2_3_LC_12_9_2  (
            .in0(N__34065),
            .in1(N__33206),
            .in2(N__33514),
            .in3(N__33918),
            .lcout(),
            .ltout(\b2v_inst11.g0_13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQK9K2_0_5_LC_12_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_0_5_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_0_5_LC_12_9_3 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \b2v_inst11.dutycycle_RNIQK9K2_0_5_LC_12_9_3  (
            .in0(N__33205),
            .in1(N__33146),
            .in2(N__33533),
            .in3(N__35200),
            .lcout(),
            .ltout(\b2v_inst11.N_4690_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIK9J85_5_LC_12_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIK9J85_5_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIK9J85_5_LC_12_9_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \b2v_inst11.dutycycle_RNIK9J85_5_LC_12_9_4  (
            .in0(N__33527),
            .in1(N__33437),
            .in2(N__33530),
            .in3(N__33019),
            .lcout(\b2v_inst11.N_6063_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_7_1_LC_12_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_7_1_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_7_1_LC_12_9_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst11.func_state_RNI_7_1_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__33380),
            .in2(_gnd_net_),
            .in3(N__33307),
            .lcout(\b2v_inst11.N_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQK9K2_5_LC_12_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_5_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_5_LC_12_9_6 .LUT_INIT=16'b1110010011101110;
    LogicCell40 \b2v_inst11.dutycycle_RNIQK9K2_5_LC_12_9_6  (
            .in0(N__33521),
            .in1(N__33674),
            .in2(N__35204),
            .in3(N__33508),
            .lcout(\b2v_inst11.un1_dutycycle_172_m0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_12_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_12_9_7 .LUT_INIT=16'b1111001011111110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_3_LC_12_9_7  (
            .in0(N__33431),
            .in1(N__33379),
            .in2(N__33023),
            .in3(N__33306),
            .lcout(\b2v_inst11.N_3099_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_12_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_12_10_1 .LUT_INIT=16'b1000100010011001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_2_LC_12_10_1  (
            .in0(N__35089),
            .in1(N__33170),
            .in2(_gnd_net_),
            .in3(N__34056),
            .lcout(\b2v_inst11.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_3_1_LC_12_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_3_1_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_3_1_LC_12_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.func_state_RNI_3_1_LC_12_10_3  (
            .in0(N__35090),
            .in1(N__33086),
            .in2(N__33080),
            .in3(N__34058),
            .lcout(\b2v_inst11.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_5_LC_12_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_5_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_5_LC_12_10_4 .LUT_INIT=16'b1100110000010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_5_LC_12_10_4  (
            .in0(N__34057),
            .in1(N__35199),
            .in2(_gnd_net_),
            .in3(N__35088),
            .lcout(),
            .ltout(N_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GPIO_FPGA_SoC_4_RNI498D2_LC_12_10_5.C_ON=1'b0;
    defparam GPIO_FPGA_SoC_4_RNI498D2_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam GPIO_FPGA_SoC_4_RNI498D2_LC_12_10_5.LUT_INIT=16'b0000000001111111;
    LogicCell40 GPIO_FPGA_SoC_4_RNI498D2_LC_12_10_5 (
            .in0(N__34961),
            .in1(N__34249),
            .in2(N__34949),
            .in3(N__34930),
            .lcout(),
            .ltout(b2v_inst11_un1_clk_100khz_52_and_i_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINTLA9_0_LC_12_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINTLA9_0_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINTLA9_0_LC_12_10_6 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNINTLA9_0_LC_12_10_6  (
            .in0(N__34826),
            .in1(N__34078),
            .in2(N__34817),
            .in3(N__34795),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIBNRBI_5_LC_12_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIBNRBI_5_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIBNRBI_5_LC_12_10_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNIBNRBI_5_LC_12_10_7  (
            .in0(N__34661),
            .in1(_gnd_net_),
            .in2(N__34652),
            .in3(N__34649),
            .lcout(\b2v_inst11.dutycycle_eena_14_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_4_i_a2_LC_12_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_4_i_a2_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_4_i_a2_LC_12_11_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_4_i_a2_LC_12_11_1  (
            .in0(N__34555),
            .in1(N__34396),
            .in2(_gnd_net_),
            .in3(N__34248),
            .lcout(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_rn_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_12_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_12_11_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_12_11_2  (
            .in0(N__34067),
            .in1(N__33919),
            .in2(_gnd_net_),
            .in3(N__33726),
            .lcout(\b2v_inst11.g0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_12_11_5 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_12_11_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__33665),
            .in2(_gnd_net_),
            .in3(N__33639),
            .lcout(\b2v_inst16.N_208_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI9CS7B_1_LC_12_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI9CS7B_1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI9CS7B_1_LC_12_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_off_RNI9CS7B_1_LC_12_12_0  (
            .in0(N__35339),
            .in1(N__33539),
            .in2(_gnd_net_),
            .in3(N__35930),
            .lcout(\b2v_inst11.count_offZ0Z_1 ),
            .ltout(\b2v_inst11.count_offZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_1_LC_12_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_1_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_1_LC_12_12_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.count_off_RNI_1_LC_12_12_1  (
            .in0(N__35672),
            .in1(N__35654),
            .in2(N__35630),
            .in3(N__35627),
            .lcout(),
            .ltout(\b2v_inst11.un34_clk_100khz_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_0_1_LC_12_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_0_1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_0_1_LC_12_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.count_off_RNI_0_1_LC_12_12_2  (
            .in0(N__35468),
            .in1(N__35369),
            .in2(N__35603),
            .in3(N__35819),
            .lcout(\b2v_inst11.count_off_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_15_LC_12_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_15_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_15_LC_12_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_15_LC_12_12_3  (
            .in0(N__35528),
            .in1(N__35513),
            .in2(N__35489),
            .in3(N__35332),
            .lcout(\b2v_inst11.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_3_LC_12_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_3_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_3_LC_12_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_3_LC_12_12_5  (
            .in0(N__35462),
            .in1(N__35441),
            .in2(N__35420),
            .in3(N__35393),
            .lcout(\b2v_inst11.un34_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_1_LC_12_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_1_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_1_LC_12_12_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.count_off_1_LC_12_12_6  (
            .in0(N__35295),
            .in1(_gnd_net_),
            .in2(N__35333),
            .in3(N__35358),
            .lcout(\b2v_inst11.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36579),
            .ce(N__35939),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_0_LC_12_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_0_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_0_LC_12_12_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.count_off_0_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__35328),
            .in2(_gnd_net_),
            .in3(N__35296),
            .lcout(\b2v_inst11.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36579),
            .ce(N__35939),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_9_LC_12_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_9_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_9_LC_12_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_off_9_LC_12_13_0  (
            .in0(N__35219),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36603),
            .ce(N__35940),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIM49AB_9_LC_12_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIM49AB_9_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIM49AB_9_LC_12_13_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_off_RNIM49AB_9_LC_12_13_1  (
            .in0(N__35225),
            .in1(N__35218),
            .in2(_gnd_net_),
            .in3(N__35896),
            .lcout(\b2v_inst11.count_offZ0Z_9 ),
            .ltout(\b2v_inst11.count_offZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_9_LC_12_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_9_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_9_LC_12_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_9_LC_12_13_2  (
            .in0(N__35783),
            .in1(N__35812),
            .in2(N__35822),
            .in3(N__35755),
            .lcout(\b2v_inst11.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIVLRAB_10_LC_12_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIVLRAB_10_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIVLRAB_10_LC_12_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_off_RNIVLRAB_10_LC_12_13_3  (
            .in0(N__35789),
            .in1(N__35797),
            .in2(_gnd_net_),
            .in3(N__35897),
            .lcout(\b2v_inst11.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_10_LC_12_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_10_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_10_LC_12_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_off_10_LC_12_13_4  (
            .in0(N__35798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36603),
            .ce(N__35940),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI843EB_11_LC_12_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI843EB_11_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI843EB_11_LC_12_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_off_RNI843EB_11_LC_12_13_5  (
            .in0(N__35762),
            .in1(N__35770),
            .in2(_gnd_net_),
            .in3(N__35898),
            .lcout(\b2v_inst11.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_11_LC_12_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_11_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_11_LC_12_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_off_11_LC_12_13_6  (
            .in0(N__35771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36603),
            .ce(N__35940),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIA74EB_12_LC_12_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIA74EB_12_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIA74EB_12_LC_12_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_off_RNIA74EB_12_LC_12_13_7  (
            .in0(N__35744),
            .in1(N__35732),
            .in2(_gnd_net_),
            .in3(N__35895),
            .lcout(\b2v_inst11.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_12_LC_12_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_12_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_12_LC_12_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_off_12_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35743),
            .lcout(\b2v_inst11.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36665),
            .ce(N__35938),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_13_LC_12_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_13_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_13_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_off_13_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35725),
            .lcout(\b2v_inst11.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36665),
            .ce(N__35938),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_2_LC_12_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_2_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_2_LC_12_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_off_2_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35695),
            .lcout(\b2v_inst11.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36665),
            .ce(N__35938),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_3_LC_12_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_3_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_3_LC_12_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_off_3_LC_12_14_3  (
            .in0(N__36742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36665),
            .ce(N__35938),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_4_LC_12_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_4_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_4_LC_12_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_off_4_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36715),
            .lcout(\b2v_inst11.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36665),
            .ce(N__35938),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_5_LC_12_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_5_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_5_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_off_5_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36688),
            .lcout(\b2v_inst11.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36665),
            .ce(N__35938),
            .sr(_gnd_net_));
endmodule // TOP
